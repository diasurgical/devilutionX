MPQ    c�    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h��G����|I��+N���
V��I�S���a�г} �7	M�9'�,x��0l���,���:z��e�u���{�b;'�ߝ����E�D�FɽWD�[a�ɛ>;��(k�����uKW�YF�Y#b�{�R�N���
��9�J�vn,����q�!�Z����<oLx��s-�E�5�甓�:]v]�%�ɝCѯ�{�1�'#��
��Ս[
�-9�i1{��S�&����k�R꼯-��g�?�IO�[�o�X8v1G
FE��w&j���Z/��N�����T~���S�=_������������3Ltl�	�̲+�
��Zi�׷�镻���ٽ?"q�!$A���n�0�c���n}m����ͣ��1���qR&�ӗ�ZRw�NI�+�̎����u��[V�*���(^Რ]�b����̒�\����_����m� 蟌�q5����rU��X�e��oٰ��������*[��l��He��x�t�u��u��}������ŮN�PjAbZ�5��7�ŋ�m�>��h�d������=�s��-�7����G p���x�� ���)����%J�=�:P�?LQ�)�A�A�~��
�Ƴ���rYB��~q�	BY��,��[�<�#�䖧QoX �}�+/r��z�e��]���{�Ux�[h���(�=$�{ד���q���iBI��^b�����I�f��7�ʟ�qc��XK�z�����7.���DU��e�J䥆��Y5ʧoS�L;��Z� 
���fXaknqIT�(A��~c�;�6��(�w6!ac�{�w�8
Y����6��h1C�W%�b�i�B-EI�Ϥt"&��^c_��0+��c�[�Ņ��%������Cm!Ɇ�B�;�G\�I��t���Ԗ3�0Oen1�Ъ����@�p/����?ͧ����Gs�6d�B���6;-aQ��2��I����Y���K�� H�q�@J�;Kg���G�P�'oo�'7�l	�{{�~��o�i~e�7��䋶:��qD������0ۂY���6u����u��C�8�z3�r-�q�
�d�ܾ�QIz>�j���G	���+��t.����*��g=����ǄW�k����Y�5ލ���.�����z�M��S`��\�Z����7�>���NÿT�����R����`k�
�-��=���L汣���,T]�����w/�������Pm�n͋���F��%�S8���4��������T�y9.��"�qn]�z*(��Y�j(�u���q�,Yp$��P���X�B�Q�-me�lW�]Z��'��Eᒠc��<��H
��)tCh�{0��Y٣qQ�x�s�9iF#te�1��S�/wP�ζ�iY<J�m�fxJ8g`3�KM=�1��a�2i�n�3���;���s*�1�2@��tO��.a�Sҏp1�5)!F�K ���~��1�"	4�W�N!�_ȤqA���=$�P�-?��̝����޷<I6
�y�F9�Z�(d��pK����k����ϼ�]�+|&W	����.�#{���Ɔ������{u�7�����1�F(� ���u�H�탼�������^�XAP��#.s_���ǘ$#��Ԫ(.#��(�����Τ#��[��/PW������	��L� �����M���ŏ
�gB��v,�jk����X�>���� ]�êp�K�l������ٹ|g�����ӈs���b���O
�/�����T��\�u\�Q�إ���'Κ%�>~��o�?�������}�ܯ�y"5�Q�5F�H��D�����0ɑy�x�Pzѫpz~x|�:�.Di�:��֛��b�4��q����m�����ru��h�qjR�{��j�U˘s��;��j��t� h|�a��s��i~��a𾔃�H�VnhDV��A����`d�!� y��4̈��Iw�	m���M����gEB�P�~q��-hD�K}��w{��d��޻��.cE��A�Kp9��[Y��.lI�����䐷�&7oKVVQs˚��B�`~��O���$"%�ǭ�=N��V.�����#Z��[C�˽h]��gW�~�0;*�K�H3��r��������	~G}�y)��#�̃l8� �'o9]����Bʊ�\�]�ג�.�4�8����3�7C���#��Fu��Hb��M���^���"�JU�����ry�geSk�U���܏��*�Ԉe]O��~��w���iQ���V����ߕ��mR>����|�e?�� �������q# ����ri$�^&�?̝y������{Wl��� ��B�57qe���MO�Յ��ޔܿ��w���"9�|̗E�X#AT��Y���p����j�40&��?�JBY�yR��;�k�B��V�KDi����{����h2���'�E�z�9�qYPeo�@��IܻJ�\�0�˥,�gV��iyCP�qW�Ó���f���"#0�QN=zﱒK��B���@z<f���P{�6u��Ǣ]b6�gmrRO#��V�0=��+[p�-� �%��D^s���|ps�#eQ�J�I/�6k�%�>�H�-])R���0ml�l4ax�;�k��pp_�he��+�5�\�>�U*��fCy�w��3�$k���ͅ���&��j*K�\)�>}!q_C�>�=�����^�����hWP��9�0̣yH:с7J��*�J"�߯EX��5>8L���9~�C�q�&Z���V�N#���-��� ����z٪����q �wF�"/�|���A��N u��־m{^#升ɇ%t�|��5�~Ş�;��C��}�1t���,�����fu���{��z����<����ױ���Oݜ�,���f��|+�d��A��}�HE�\�Qh_��F�D�9pԝ>�G��3���"U��hr 2d�1i�/vt��猩�9d�m!e�X�Z�|���%�'|��ߥ�n���T{�����#�5i��}�S7��J�kx�F�|u�" �N+����-9s�@F�H<+o\�Y]ω(�D�ޒ�h�Avd�I2 a�*H�"2׷'���؀k,Ӥ��Ub��ѵ-��nm�k�bb�Z��[�PM�pQk�.	��gi�"���|���)a�r�Y��{k��NE
)y�9����4��(�q��3GՀ�Puo�o�E�����N:�+�vx�p%NoC���{�.��lh�K���[�69
�w1�u�Sv�Q&(�b�I �M2¯�'�gCrIjf�ܚ<�X�GE^=���r!}���p�u_N�PE�m�g��S�`���*�����Gg�3Y7�%�	0k+��J���{�r���d��G�?�D%!?�G�
0~���}���A��%t���&�	��KE�)rx+��l�\��͜�t{Q��J;�-���65���������_=k8��-��������:�U�A��`��o4%K©Ԅ�����5�����3��eM �x�2�t-�0� ,���5�U-(�ƃ���mj���0�7ݏ��(�>� 6�d��k(ϮX-"B���G[e0���;rL�}¿�ǽA�`г=6��P�mL������-!�������\��aB�xq��r�2W���w����<�0���d}���(z}����}�r�7K��Q�]]��{��S���'�9(�{D$3˓^�q�i��1�$Z�^���f�RI�璽��ɽ����ڐys'r���[�U|
]��xJ��M����5E%�S�y�����*� wG��z-k���Io �A�g�c_H63��!\��y��wV1^Y���4hƬW`�*�H-@�	����"�^^"^b5+�+p=�cE� �� !��XhiC:|{!�tE�D;� \�=��T�υ��h��O ��1�>�Q��@���/V�?�����f�Fƿ���6�7�,4ce$;hk�)�ҰD���}��E�ЧX����!�v`�p�<�K�o_��'��L	�c��ԙJ��T�#en_�ߦ$�.3�,
n�r&�,���]����u:�e�p�섞S��5�oэ����-��?�ݾ$�ezٯ�ϳ�G^�H��^����t�m5��E��Y=/d���C:W�f��^M^�P�4��`Ag�ǉMSV<`�)�\M�˿��R�M�LCÚ0 ��L�RJ\�[}�eԛ׭�P�"��LaI�ȧ���g�f�.Ǎ�g�/KN�����OZmDQ��k%=Á,%th8�]4��Q�}�>�y�[���}�n�F�*�<Y��p�sG����G.�$! @�b'7�}��W�e������Zڦ̖B�XE\VRc~�&���:��`$}��D�{��Y�N�Q$�osh�F^�D�*1�mkϊ�b��u�it�>��)�x%��g���šv�=�n� �2$�-nǴ�|V;��rse^���l�o���
kS�d�1ѡg)�5�K۔�,9~�́<	/ı���s_�-A�@GԸ^P�X�?�W��#�{�/��H�
vdeFT	����ɷK�Z�c���̱�X��+7�	�ε��#V�c�b��]����y��`�7��J���6�(�+���uk�]�~W�y��Ϥ�a$�ӧ���M�#id��G��Oǔ/V��$��m&٣{.�؛w��@��>;��&�W���}%�*�N�pI� ����$��M\�@Ŋ̋g�	�1F5��/ե)`�����]��p���loۢ�5��r�3C��cUQ��
Qb��i�Jb/6W�砗��w7�\X/c؀=��b��%Un՝���?,�钛���*}Kl�TZvӌ�{5�{uH� �D�A1�d�>��a�������Rw~��6:@4iŐu3���ϡ̽@4H�-�k�ԟ�BO�UC�u�$êjɦװ�U���s�!�*�}:P� c`n�1�.�Hi���ak���,�V�ǒ���A��#߻m*��~�y)|@�ш^w�sX�^��M��>�a�B�`�~���-�.�K������26�ގ��ڍ�c R1A�=�9L�[4z*.��N�!�_�
~o|xQ���?�`YN{OL"ʭo�%
_����	v-VIZ�;�##5�"[~���V�b$���^;�W��r�/3��,�X��j���ՏadG8J_)�<¼G��8\��'��텈F4�=q���D_��.��ݚ���#O34�m�t����*���x�>}�����zV���e޺��3Ǎ�m�+g�/,r��p[��WҖg@h�VU]�É�y��wn��$D���εp���I��m�����|륞���:X_�LĶ�}r[a�Y�q?'�3������lo"��y���}�5�&���Z�O-^���,�ޯ�ƍr戫]`/��UEn(�X?bTF�×��)��ͪ�~��CJ���yM�w�^����x�q�D�mK��B���ۅ	bv'�N�z`6��%ye�߂�Јh�����8�0�`),%�L��)�y^�q�L��ڒf�9"��oQI�T��q�O�����KG���'�q�	�;��]]@����R
��q==j��[K-��[0C���"n�TL2�s���Q���I�o�k�H>B/��:�)M�hǋM�X�a����T&p��_��Ͻ|�P5���י�
*�>f^���3���k9��� ���!Yt�z��K���)�w0!��yC�*-x��җ6�Y[�	GW�b90�,�!�Hh7�s�ŏ���x�Cv	�>S[���;YJ?C�b��~:��__��~B#�]w-���q��kx������l�w��/u��դz�^H� Pw$j�mY/��T�_2i�7�dP����c���e�^}j�����5��d����ف0�a���U����参�ȃ����O8 ��`��)�|�b������5fEo������_N���H�TC��4���w��aU�hmz^d7�$��Z���c�Y9��HĞI"Z��v��j-'�kd�`@,�6�-T����)��^n$��;�x��7E�ˊ�e�aCua�L�)pm� �U-�Z�@A��<����㲉C�Ys�C��v�۟2�r�a����}�	���v���,N�6�0�����8�m�Y�DEfb���v�yM�k�tãil�5s��7��F<�a�p�Ya��{F��N��g
�T9���,��l�q�ӌ�S����}o ͩ
�E��V�J��:�hov��S%�X�C��{(�]�}� ��;.�[���9%z1qSQҔ&c%���H�c��`g�ĬI���*vX�2G��i�"&�"�Y_�ySN��t����BUS*�/�.՝��-Ģ$�3��^���	��+d����N��"�-`����?�8!Z�����O0YDFs�}��q���ܗp8��jO�&�_��Pe?���+Hu�����ޜ��s�&�`�I�*��F�i�>�����_i�!:͐�6 $��/}�R��IU,
�[o����d�B���� 0����an3�e�LXx��6t�q�]�������rۡx��ĕ�jwqg�+�:78z����#`d}�9�F�b���-���bG�z�fڡ�VJԅ��B�� ۛv[=��CPทL����*�H�� Ǫ��R}�J��B���q����AǕ���� <������yVl<}�P�rp�߮���]�F�{}������\�(���$�ޞ��_q��i8�+��P!^�y �&I�����L�OA������Tm������Uw"C�!J����J5��rS`�T��'��  ZW��9k�iVI�E�AxP�c:6n{j�Q�!W����55wJY�7Y�,@Uh�h�W��f���-;>�Z.{"��^=ym��+K��cUNŻ��e�Գ+�C���!7����;}Rdʪ���ʔ����=O�k31�����A@��x/��p�P��\���p���a6���姓>�(;��y���%�?���R��o���n���Y�汕ߢo��FY�o�-�'�>Q	��t�%<���e	����N�Ȥ����h��O�8ٻ�Yqu�D�k賄�(��@Ѩ
��g���N�_��ztͨ�ʄ�G��!��Z�� W�t$D����ߔn<=��S���WG����kzؕ��̳;���V3=M�I]`���\��D�z�©m ��Ǉ��u,n��R�i�V�
�E��hWm�=�L� �Ȃ?<��8���Y��d�/����S!þ�nm�SыFw�ü�n%��8�G�4_f��;z�:HKy/���z=n���*^��Y�pu��9��R͎�b#�$����=�e����cb&e�-�GZ�o�]��E�9�cY ��*���7�I�Y��{�9Y-Q��
sC�F��߼b1�a���=�DT�i��[�c��x 3�g֛X�<��=zc��{~n2�Vn�Uu�;t%2s�-��h�P�jC7���SHY�1�-+)E�K���g5�g��	*���_>��Aķ��3��P��?�d���Lv��g8
1oFox_��3�/KKM��Zp���P���^+�1	�n��k#1�c�<]���'���/w+��7@��I��rR(�֗*�wu���y�*�q��P����N.����V#�ue��Ս����!��[��{f�Mp�����<<��⺹�=�WZ�J?��E�܄�eL yF��_�M��Ņ��g�*H��"��l������L��1E�]+��p~�]liX�]n����̱����>W�� H�b2k|�E��/��S�[�ɒ�\�,t�[��ǝ>�%�䝙ն?�4�V�F�E�}�M��/���Q85|6�H�DP����F���U�~�D:�Y�i	�n�
̿u����8�4�^��FZ��㫈���'u��\�kjȚ���U��srk��e3��K� ^Ϝ?�-���i�7.a�/�l0�V�F��FUA� ���З�#(yDB���C�9.�w1�7��o�M��)／�BB�C~���-^9)K�ڃ�V�5o���^��5]�c��A�O9���[�.�i9�D�]����e�o���Q��0�c`4�]O���
*�%���c�F�VdB����#:�[����8��]U��4$;������>f3�����z<�ð���RG�0�)����f}87b!'�2�#��88��� �MV.)Cu���j�3o�l�@��J<�;˼w;;��U,��m�mؘ�����hAg,�-	�����4�B��JCY]DX�t��wɴA��VM�U�}���x,-��m�-�}ץ|J�W�`<:�t��P��'����r��v�T�4?�xN�n�W���l�e^�TF"׸P5m�ܭ��O��y����֍�t}�8����ާE	iX��Ta��RN��D�D�}���!��)hJx�yH�Z�\9ϸT����D
�K�o���.�8�܅L�'Ox]z�ᶧ
eeO1�����6����0�),��B�L	�yy��qM'����fO<�"Y��QD��gq��
� ���2Q�������|��V�]X����UR��ގ��=�D[&�h�����"��i����sN�Q�Z�I%6k�q>}�i�Ah�)Hy���Mdd"a����a;�p���_2+ν=5�9���`*w�8fy5Dm�3�F7ktuZͻ�"��Q����KX��)��+!J�Cc6c���2�wTTQ�m�W�1�9K�̙�H��7�&�`ip﷯�}/1A�>n�s����4��CZ���\�*��7X�VV#j H�S��[	F����6T�+8��gF�w��P/0���{���� +/{V�m�s�C���_���__k�BŔ�w��U�Hh=}d��Ƽ�K�L��o�ٜ������0���6���,�G���#O��*�O����|!���m�@��	8E
�½��[_�YO����o���4	�a�?�=�uU�t�hh�d���ӥ_������X��#��LZ5�ĉ��A'2p����Q!Tqr&и�뿙cMk���s).7�m�����|�)u�mE��|�;�Q-ob@<��<�U�ψډ^N���s���Av��I2F�}aӖ�����Z��,����×G��Ӷ�m�����bh����"�M�}�k���A�0~�M�8��[aˎUY��A{!��N8�=
_��9��ׇ!�'�Oq�ܾ)�o�f�Vo���D)�E��1���:J��v���%D�UCb��{Oj��_��gL얊�[;��9@Y-1��S,��&�r����C"��>Og�7lI��lܐ7�X�L{G��ɥ�q�����4QNӚl���jSe�ɟP��9��e3}J��E�	W�+?�$�T����W�<���H?SL�!u��� ڝ04=P��<}>(d���#��k�%�& ���˞e��#�+��A�����ے*�lt�G��A���#��Z>�ց��م���I�_�/�����Ql��x���<�NO�U���V׭o�m��4�4ۢ��J�˪I����e���x��6t�P�v����o�Kئ�|����EBj)��&T�7����p�60�d�?.�!b��$�~-X?ޥ��G�j�!���qBD�s���}sn��<w=l��P���LbXt�rm�c���{���h
���,BSz�q��(j)��P���#f{<�3����Z�����6}�'K@�)r+8���2]S#l{X9z���]+�(�g$�R��ŏq ,i����gL^l��sI�M��H���
�~���r�/����ݑ.�UrZ��vT�J=�	��>5;��S;3P�J���U)) �\#�w�k>/I���A�XKc#06��	��2!Rmh�/��ŵ2Y��짓bh�+�W֬�:�u-6�nϵ�"W�p^X��+H|+&��c�w��V1��(�9C��?!R��;�;X2lG���Er���Â��dO�E<1�>�G0�@]\�/��u�뵽ͮ���xA6��Y�"q#;����_��:|���&�*��V�p��-���깢�k��A�o�G'h�y	'�*���Q ��)
e����<5K�VҢ���q�"y��I)4Ōup��fW�T�/���ò8��d����/��T�z<��u�G�z�Av�;�t�:������=e�,����W�����zS����*޳*둿�M�]�`�W\.1�5�;���D�B�PH��P[�R��,�Q���#n�XD�LW���]�����.�d���;/`%�i����jm:v��!����f�%���8�/O4�M,����Ur�y������n�3*���Y�#6�)L��+H�}8�$Q�����\���ve���hMZPXx�ER=zc4�K�eS���k|��y��{a�Y*�Q�s3lFԟ�z��1�u��@�g��R�i�^���<�x���g����-�=uB���<�2��n�Pr�7;O��s�/�d��e���?��Sn�1�V)�tlK��t�����	%�ڧ_��_�#�A�N.Ԯ3�P��j?7j���\`qM��M��
��F��]��Tr��KY[�<r���«�=+��g	�� �#���wx�������?�k�7�5����ͺ(y�e�du����t?���ٻ�EȆ���D�i#ߦƅ}.�����_�n�ة�ٙ>�����Ux�,�r��t�W���!��`�f�� T��e�M��.ŀ�AgSl�����k����ß�l��]�0�pyRZl�ě�f���ԯ�)���y��;��b�o'�@r�/�e��}Yɭ�\NJ1�6�Q�ئm%�-���8l?��l����`��}A�H�
*���H5�H�<D��P�ښU�ʡ���4!��x�~)��:v�oi�H+#�0�áԹ4>]ɰ!(�5V����u�o�yYj�IP��PU�GIsM����ǲpg� Y^�Lꋤ�iϨ�aa�GTLV�'�A�z��q�W�R�y_�86s!��Fwl�Քa
M���T(B��~��-�c@K��փF7���ˢ��N���L�cv� A܁�9	�[꣮.*X�ߐT��˷��o|'�Q��'�5$�`ΐO���\% K�ǾV�7VJ�1�#봿[���9��X�Ȍ�;;P/��Ă��3��F#�� �r�ߧ�{-G�7)1�w�=H83@' �+��)�3��m�����.D�ݐ���E�E3��?�����������2X��
�p��H���0��i:&�c��gvH�谱�ya�M�e���Pq]�%�ow$��ʚ��෵��Ө�?hym#=�x�O|�\D����2���0i��;��F�Xr:Pd�O`�?���)+&�"<ele���/��G:5�����O���4����]�h#~�<��-�E���X�T����_��������J>�d��J\iyC�yL{@�s>����KD�֗�Jʉ�i�9U5��U'���z�����e��K��fQ����-\D0��,�d9�	Ky��5q��*��� f���"���Q?�����ł;�4�%�v��mo��e$�q�:]S���xl'R�ꎧ�!=`�=[~��z���4d-���s	��Q��I�ƗkcF
>�(�ܵ")Cz^�An���a�?K��A�p���_m�`���5�{�OgU*2Z�f�ù�>�3��Hk���V��gk�0m�K�)Jo!��C>bi�j��3�O����+�W��c9fz]���H��7��V��b�ޯ.J�Y>�ك�w�.�C�I0��'���/�gM�#%�cc�g��!�t�+�ߪ���b	�wW��/�e��D�T�� "��GmL���~����sڭX������w����F�}����@��5;�>�ٷ��W7
����q�����#�~�O�&M]^,��1|��A�Hlk�.��E�o��/_(��w1������<_7�x�]UQ[�hc��d�<�`����s�O�%��MR��qZ����T�'�������l&�T��Г���x�?c�ny7�R.�I��ƗG|uWC��Y��v�-
�9@7�?<<~1��NF�y˙�O����9vH2�wAa�|U�3�Xb��)YG,D������n�/m�`���b#�{��u�M4Xk�`�|�.��ɓ����ja��QYW��{���Ns"�
���9��G��Kq�9��.�A��o8���gE~�h� �:BvɥQ%�gkC=b{���ݓ	��D���[��9[X�1g��SK&�߂���>�z���]gt�OI����e�X�)�G�f^�X�v����nGN�o,�~v���S��P�d�����!�X�T38����	+:�F�Q�CN���X�!?��!�-}�{��0���T}��n��]��&����&l%�F���@+����=��1��Ǐ���\m��r+5rּ�V�t&�ͳ�_�.�VD�l�H���8��M��	�Ub��QSoEB.�ړ��O25���˅�Z��e]x���t>P$��`���&���]��W�m�:�j� U�!�7�Y���Q]Nds���A��_��-���;Gl�ܻ�֌Z����X�,�#=1eP�Z�L���-�"�~���s����'��w�B��q}��������>T�<�䝸�Q�=�k�Si}����r�T��|�]�8{3�ųGŸ�K(�a�$D�擏�q�i.Md���g^N~07k7I��	��ΟŐ�3U��
�(#�$�,�JUm���ѫ�J�.�1�5�]&S�{��.��Xk ���ҡk��KI�/RAn��c�Z�6����!�!M[���p*w�۲Y0���"\h��W�:���!-1m����"��^s��+��c�����j�M��i�Ckh�!m!/��M;3k|�����M�����yLOQ?	15ժ��@8@"/PO������\�Wrs�3ƶ6Я�坲A��;Jr��85�5a�����O�!]��[a~g�'`��A���<�opl�'#T�	B�
�j0��)�Ke?�J�з��]H�])5�C��������oP�u
 �aTք���f�}��z��]0���瀾��rz�hǩ���Go
T����V�tQH���I�
�a= ^��wW�쪏AD桖Õ�s����k�M$�G`��\^����Hy��,�����+�z���R���Ls�v�'���R�s�*L��V�8�'��
��獐�/\<���Ѝ�?m����zF�24P%Ef�8�7�4U� ��p�iy%�ۛ���nIo�*�{�Y�����~��ȨE��mt$�)נ�~��.f�מe|$��_�ZaӖ��6E�`�c&���A��m!�X`�}b{A�YE	Q�res�p�F��1|�[ϛ�Z��q�i�T�Y��x��"gL�d�r�~=pA��12U�*n�r��;*-!s,�՞Z �`� ��S���1"��)�yKl�+�'ڝF[	 #���2W_��wA���)΃P���?r�p�S)l�˷��
���F���:}M(�K����ש����¼i�+h��	7�0T#��S�����.Mt����� �7���7W�I(T����u<��o Ə'��� �:+D�D���w�#��������@�)����^�Px�i��ΐ�P�ǉb�˘W�;�"��{&ф��� /�!���FM-��{�&g��z�b����;ҥ|��êZ`��	�]a��pt?�lQ2��}a����������b�v"�bh�j�;*�/Gq������,\ɇ�����/%&�+����?=���	��{f�}�>i����=X�5��H���D
�S���qk�<���~d5�:i���[~��%����4�{���ПY޷�&U=u�S"�t�j>��(C�U�1s(}��{[�D T���f�_B'i�9�a����"��VZ�v�sBA��u��9��Ϳyz3�rk����w�r��/s�M�2t�r8tB�O�~�i�-T��Ks$チ��kH=��^���[c1��A��49��	[��.X
��zx��W�P�o7�wQ�����`�O��p�@�
%����r:H�V�r��R#�O6[/�:�ԓ�S���$�;��43,3pE,^���;���z��r6�Gi^�)L׎���>8�#'[�؅Y�w�.&��ȗ��ÙL._������ �y3���E;���s�����c�(�_����#F��k���&�^-�gфo�x��8c��Y������}�]z���jj�wc�U�u,�(�s�Ӄ���<0m�|��s�| �p���s�M~x�����݂����ur��)�J^N?8ӣ��X�=��l�LQ�
r�.��5�5��UO>���� � ������r�hqE?J�X�nT 9��+B�zP�s�u������NJ�Gy>F����.H9����D ;0�%�.����ԫ���'+@z����Ide[�҃a��6��D0�ߜ,6�/��(y��"qCܺ�k�f�&g"�"CQ:}��Х��-��O�Y(�_�HdN�"���f�]N����V9R;:9�¤W=�E1[ܬ����X��_��]�s�fwQ���I��k>�>��Z�w#�)>��ǜ���� a���WhKps��_�m��M��5��ת��*�0f�qWc�*3_h
k�͑��6E��܋�K�}A)1��!���C�?)z
�h�PJ8R�#�"W<�9���̏צH��x76�{��|vi���6��>�H��e���`C�&����Ӹ�G��d�#��~m��v���j�f矪a���]��w�#/��&֤ϡm ����m�d�y�p��hq����Ŋ�c�|{m�DW};�������Ω������!e�ҵC��4Ƭ���b��yO�OI��G��۲|_��#eF�i�E@����?__��2���t?�*���U�a�h^�dHט�ɘ�/�;�����ٜ���@�Zk�ɉ���'��GߑO}���Tg���n������ەi�x7V���Ʋ�vu�8;���+˱/�-��%@2�<�N�E4���hF���M���vP]�2|*�aɂg�����L�D�`,�R������N��	ҵm�l�U�qbމ}���%M�
�keS��,�fo-e��)��wpa+vY��u{�*�N��
���9����=�ߏ��q	O�9:��xos�m�zƨEy���[��:��9v��l%:�C�{�N��.ӎ��A>�L��[��9vw1⿬S�g�&m`�2e9���g/}WI���܆��X&�G1�&��	ݿj�����N	e���&әqS�-ߵ��>��=�ĳ�3�-��n	���+�h�������ê�|H至{?��!��I��^0��> }tɑ��Q��2)ꛋ$&6"���q6�U�+�a���Ly���w�".m=���w��7������������=t_z��kKt��dw�n�8]�O���2U��Lato�6z��j�O���)�`}��e���x��
t�o`�kS��J�A��2�u�jH�ߙ
�7I���|��l�qd� |��A�Ϛ�@-��ڥ��qG�z%��ܩ֧�܅i�S�3�[�L)=���P���Lyѻ�噙�#�q�۳]�Ԇ��HB��PqxEO �����/�Yb�<v���Z���x��'��}�5����r�~5��u�]I<P{q᳂�I�((�C�$��Z�J?�q6ԭi������r^�����sI܇���.��hP�N$����庞^ [���HUh*��,#�J��V�9�51[S�l׋�d�틨e ����-D�k�ҬI���A��%c˲X6D�"ܽ!Hi^��=�wBT�YK��읚AhxlWLIӵp�-,F��k��"ͭr^���!�+�4�c*�Ō�����5�C&��!���1Ҩ;�<�N��{I����9��d�OY�1P&_�=�@D//B���!c � g������j76���r~�`�;T�ܝ�
�0f�cO��D�<���e�Y��b����� �7i�o�;U'�7	]����j����@J�e�=t��R6Xz�a�P�ݽ�w�Ɉ����u�9�\�1�
)`�!SJ��b��%�BB��_zE�J����G�Z�����qpnt���`�9�ERR=�F&��s)WX�ѪJ(��T�� ����D��8�M��`��\�ZJ˫�z���[�8���8���)R�E^�G�Yי���LLM�Q��S)d㍋�/�8���Xy�1��m0��,��m!�%��<8�_�4p|ԣ=I��&�y�Qԛi1�n�g�*/{Y�������F�����$"��Άҏii�4B�ew���wZƉH���PEH�Rc��0��O������/&�{���Y`;�Q%s��>FJ����1w����W�u��i�j�����x��Ug����e�=k`�ߌ2T\n3��h(�;�PsQ[��9q�[�o���ZSy��1=��)�3�KGP�b�8�U	����_o�CA�5Ԥ��P\��?��K��Pg-����
bOF�^S��?�(ݵK�۫�r���8���qT+#��	"�G�z#�MD��������c<�N7qhR��|�O(/�Cۅ�u���jፏ����U�	Ϳ�$�Re>#UiE��?l�?ɔ�C�տ��fُ�>�D_���Pi�b���zB�Wk=s{D�7�\{� 

��T�Mȁ}�vhg	O�9C�������Å��m]�ÚpoL�lz��ێ�͹��
��ަ��vb�E�6�/��/��h����\D��찣�N��%�lc��^?���W�Ζk}7�U��y��xf5M&�H���Da7�P,�� b,����b�~��$:���i���᳗���ȡ8jS44����#D������E�u�W�/�j�h�C	`U:Fs6��P���; OܐP�����i�aW�R��� V��]:�AƎI�'����y���,�!���Jw�\��ʤMʗ���<�Bsߜ~��/-�KN����6��o�ʎA�F�jc���AFJ9�a�[�M�.�
2��j����v�o�R�Q�\n�+`���O8����!�%��?�tA��x�V��3'�#�
[j���oq��N���E�;Ɔ'���N3K�������&�uw���G$�_)g�ͼ3�a8�4�'��9��T��)M�#���~k�.z�s݆����R}3 b��;�����L������C��ft
���ަU���-��Y�ig,�0^`���Ce�������]� �e�uw���O@GTA���P�^O�ޔmY��np�|[����v�h3��&�{��t��J�rp�ǡE|�?�������X\Ll[���B�ik5>=U��>7O��������T4�^࣫ɗ���E��mX
O TrSÃ���Ƴ���f�{���ڔsJIS�y9�l���q���Z�D{�� ң��o"����.'`��zLI����-e�]Ń<���q��c��0��,��&�}h�y�#�q��֓Fz/f ��"*odQ5]��x�L�;��j�5�!��#y��]���]I,��.a�R��̎ݱU=V��[�l��G]��Z�Q�G�sGvQ��I��k��>.���))9�D��j�G�a��(�ҮpN�g_�>B���5����^ *�'f�?�A�3:)|k%�;͌�*��R�湨K���)L��!v�C��da~��AE�\�~΁W���9��.�
��H��7q|��1��	֞��B�b�0>��<�mؼő�C$N�-Q�����R#�(���y�]4��k���	�X�w�v/a��Ay/�J�� �`�Gm����tM�˧��#�����R<�W>P�b�}�mX��1;�\����Z���\��MT����-��ʳ��J$�t��O��r����\|�H���}��F�E��8����_�$��������Ν�F���Ɩ����U��chY��d����-\�J�k�Ew˴��5��Z����g'C=��L?K���,T�q��I�!�JA<�dy�7�Q������uMN8������~-@9�@-j�<�Ҫ� :ꉯ%��E5Z���v��@2�PaĨU��l���c\�_�b,:���������q��4m�]���ub����{oM� Dk@�M��A�	!�Ie�2va��YM&R{��N��
0�9�	lט�v�X�q$��ő����o�#��E�EtA���:{�Ev�-�%���C�x�{ �l�ɼ���^��_[l]�9���1]�KS��A&OR�P��4z�Ol�g�O�I��f� XZCvGl�#��P$����ye
�N$z�t�x�aS�����y�ػ��ZU3����#	u�+�۴��^%�yY��w���lT?�G!���qe�0�6�2@}����e����&�V��&Q�\�<��p�+4FJ�s����x�}����������9��2��������u_Ջ�&`�����-�8B���hU�I�G�o�J��P�d��@�Z�;G�Z�WeT?�x�2�t����I�7�����o��⮰	j�#�j7�c6��1=ч]di��an�ՠ-)g���G"��R������K��t�ۇO�==�fP�|Ls9@��p,��0D���8j�6�4B$$�qs�{�,ǁT��t�|<��5�O���-ºv}�l�Q�r\`ڮ�]�x�{�<ͳ�3�.W(�E�$�#���xqQ�i$<M�kln^�m~(I�T�Y�Q�;`��i%������$�}��b��Uc�����Jn��T�5�x�S�9c����& �%����ko�QI��Ad2Ec�*e6Z����!C���@+�w���Yf8W�NhS4tW��ߵdb-'?���ϊ"�ѹ^�%���4+�[cA���'�%����y!C�5!�t�0;�<���)�e]���/�ZOǒ�1k�[ĸ��@�g/}n~�����zͧ����/�6H�Q'�/�;�~;�0�$�+�����[���W˥����4;E杪��w!��2Y�o&+'���	x�`���{
keuV��Q\r����Ok�?��ZۤXR���uAOJ�W@i�en���C{�km�S'U놽s�Kw�z��Ʃ�|G%ˆ�r���cet���;ù߀3�=6OG���kW�/W�/��2O�������B$MZX`�l2\!w�fL@�لӡ�y~��[ǖ�RQ${�B��,K��T
ɹ� dL����Է��<�^V���\/Ui�? i�L+�m��j���Gè.�%{�A8ǧL4��أ�Eց��(yy�D�n��*ʚ�Y����:C��>��7'$�:㠩�A���\���wer��yz�Z��!��ESE��cūK�~������W��?{��"Y{�Q���s�L�F��^K31rq��QK �0di��_�O�(xl9g��@Ũ0�=f�(��7�2�=RnN��l�;�Ps����ԧP�V�:�P9�S4lS1X�J)��K"�jS����i�	���p��_*�A0��c�P7�8?�9;��",b��^%�
�WF�@J�
ew��K
Lޭy!���%�<�+���	=� ��l#�̈́�(��d�[��G���17,��miZ���|(
��ur:�e�Q����v?�pQ��:���-;#��b�N�;�������v�)���
�0�����5����u�%WƳj6������z �5��K�Mc��qvgd�-�����إrn��`��N)]���pjy9l��_�I>�b�����Ӫ�i��|rb�=��1��/���G�&��y\�bq��ݔǉ�%\<S��!�?���B�Gα�7}����Qnӳ�r5�`HHֆ)D��Q�%g�rՉ2��=��~��:G0Ti�A�<,1�a��Se,4����QH�ϐ7�\V�u�{X���j��^�#U��s��QD�Azk J˯�W���U�i �$aҙ���CVЃ�� �A�Hy߂,����y�r`��C��)�wg?�e��M���(aB.�m~�-J��K)�,���塡:���c����c�7�A-�9z7=[{�].�*�갧������$�o�!Qڽ�%N`��	Os�.�v��%�����M���V�"����#|�s[��*�
o�IY%̠��;�b�B^W*�}3&1��^b�q\��p�5�(~G�z)�35����8�e�'�"O��(��$���~Ĩ�9]�.�'Y�#c��.Q3[c��{zW�����P�cn�^�3����3���a�:׏�T�og�]�hx����������682]���`��w5�g���.b>�i/�9,�;m�[�i�|�s��L�Ƀ��r�r���ͬr�=�@��?�y�Z���s�lֳ���Q�פ��5ْm��GZO���e��6�c���ȫ�up�ރ�Eu�cX#�Tͦi�>����\~�iL��V���9MJ�~�y4d@]��Ϥ�����D�cE�����
�Q��3�'�]�z�_eQM$��7��_f� �0�),��8Ȳy�z�q91�!�f;��"��Q0]��Ӯ���É���̘��X��vS�B�K]D����R�����=��|[�L���8�����U����s:H�Q"��I�Ek�v>in��^�)4=��R��P�/a��M�p)�_0����@5�)��`	�*c>�f�-Y�U3
�k`���'H�� �A�5KD��)gu�!�{sCϥ\�h�Ҟ��@�ß���W�$9�f3̅FuH\:7�����]c9�?o�`�>چ���j{�srCFA���ݸ��T�x��#Vk���������������66�S�wh�/o�\�P���E �N�B*�m�o;�&U���4ׁ�ŀ� �2!�4�A}qs게�^�o>���i������"o���H�o7EO��u�Jj�H-|R��ٶ�ߚ�Ev�%��J_S�����۶�� �A�ͪ��)^U"�ShT��d�i�ӑ��e����ˏ���p��Z�Ʈ���l'����O���@T]\1�$T��x��4��_)473�z+h��duȃ�p���'K-��&@(��<M�G��_"������2��v�S;2��a���Dr���ЙzQL,����w��3[u�?m�m�n2��bT���.�Mx�k�أ-O)����=�����qa7G7YȇZ{�,%N$ǟ
�Ώ9�n��zΏ3�q?AXr5����o��Ͱ��Eo�6�͆:6x5v��%0�4C�_\{;�"�d���� �<+['�w9��1�$wS�k�&��W���K/����sJg�B�IC��|�2X5�G��T�)0p��� < ��N?���ISQ���5
���Y�i�e3i�)�	�$+�n��L=���r���i��??ۦ!������N0�t m}�����W�7y���(&l�4շķ�K:+oJ��Dؠ�ε���f�.%魰T� %��B�m�q�E������_0��ᔀ����d}}M$�:��U3�{�Bk+oV�s7��������1I���e�YxÒOtO9��?�:�Ź7���� ��F^j~G�@�7�����Ѣ�d�A����9��R-�	8��sG}�`�~N��b�_Ǧ��^	�o=���P�=0L�/�^\��ϓl�gg9� ��q�B��Mqn=�֖7�<�d���w<l�H�
W��T]�Q}�ÿ��1rbC�"Ȧ]?�d{�(�����ɥu(�g�$U���89ql��i��c�FZ^�to8UI�A��'���w2��"��{4������� U^z���qPJ)�3�o��5'��S�&�6U>���� 稬���8k*;I&Aߺ0c���6���X��!>�Ŀ�8�w���Y���!�h.w�W�e`����-"X
�!�"C�^���+��ic|\�����o�z�YC�tz!��R'��;���3�]ʱ�������a�O��1�(��3Bz@ɫ�/�-ԍW����h>�d�6!�~�Q<�P;�H���Ѱ&�Ǭ����r2��v��|����s�-i�o�:�'T�	����u�lT9��He�����'���ҎLI�j�;��H  �Cuܡ3�R�|����T�/����Rq�aX��m�z{A:��ygG�[��-%&�vdt�T��	�߻4�=�w�����W�|��U���0ѕXܳ���}0LM��K`�s�\od�!�ɩ�m��.�;ü�%�<��R�"��=���\��GZ���LCv���a�ɣC��A��5�/m�Ղ��\�g��m&@o������[9%��8��4&+�������Zy�ʛK�n��*e�qY�/����a���֑��,$s���� ����jw(em�q�7#Z<;_���=E>��c��֛Q���>�S���n{M�.Y��Q~�s��QF�Dd���1mIϬ^�덙i�D���xG_�g�P=�Cq=a���Bv(2�Gni[�^��;�� s�p�o���Q�a䫢�S� �1s�)~r*K�m��6�n+�	���ˏ;_���AK�]Ԛ]�P4�?#�>�$O�]�䷹��
؄�F�B�����ަUKE�D��Z��.q�z&�+��7	X}���+#xm�c%�����Ἕ�� u7�xO�A��r{�(�<Q��u���`�8��1�$��͵�4�1T#˫���#��r�Q��KM��D� مDO�����A�����p��W!J"���̑܄R�C �����JM��,�l��g��W���"�'hx��uj�;�B�X �]2�vpe�&l0������9ь�RaӅ@�'Z�b9�đ,B/X���t�\: �آ*��ć`%�+����?N@u��R����3}-���vI�����5���H�4�D���=5�6�f��Bu�D�~�T:���i���J��ݡn�4*�����ܟ
�U����u���^OjoD�y�Uu��s��X��� E�
F]���i;��aM�想#6V���'�A�"��%3�>;�y�N�"1҈�xwX��� h�M��XB�^B~._�-�MK�i�2L��<~���N"��Iccb��AH�m9�,Y[Vw�.	k��K�`��c�,�ioh��Q0w��!fY`{M}O��g%��*�Kk:�V�T�#W�:[�Dѽ��s�D*�����;<^�]��V�3�<����;�k����(�G��8)��ļ)�+8~��'��*���q��
+��na.�p��|�9��*�3��ԕ������1O�y��\�7�ک�:��ՠ��O��g���ԏm6��9��K,�qŚ]K}�[b[w�YAʆ�A}Hk��`��)oT��m��܀dvQ|fw�1Iɞ���S�n.�2q�r����;�?I�t��Hَ��lQ�(蛤2��@l5t~��pyOO0!� C�Qʛ�T��s��=�E�qX xT(r��g���q���ͻ1. �P��J�1y/#P�4��_%߱}=Dq(���Y��U���o�뽳''�z��.��e�\��d��93�"0�~m,Gv��G�y �q�������fvvI"`hoQ+}A�.����펉�O��L���&��f�����]?�9����Rl���,�=L��[mL���3��)WyPEyn�s�h�Q=37I��Wk�1�>�t��H,)/�ǭ/�a5'�ț�p8�_YAt��5�u�׻�k*u�f <!��-3�
pk�«�����+ܜ��K�b�)�nN!l�VC�Q�ڏ��9�+;~��4��Wmq9�J�� �~H7�K7����g���P�����7>�U�c�{uC�~��c�Ÿ�OZ��j�#���;1�S���n�`�2��NUqwê%/�\w�:�@d r��}}�m��1�jI���"
ڙ{#����X��$fo�d}�~���&�W��*B��#3��C�8�w���]}��3L��j�OZ�I�q�#�&|�{������E�J�޹�_p�i�c�r��ŝ�K���6�d�FU�5�hO��dY���LW�����;ֻ�jI����Z<�U����'�e,��~����T�fR��d���HrqӕZ�{7g�t�5����WuC�6�K���b�K-vh;@#�}<��$�v�������;Vףe�;v��2M�a�T�����D姙�9,0u��R> �n����mޟpfG�b=��M�M`k���h�7������;����aR�YC	�{h��N_��
f"D9�w��N!�Τ�qZ���>%��3�o$�/�K��EjE��l� :�t	v56/%��C�f�{v�����������]8B[�Ln9ǔ�1S�.Ssy&��q←�*�����g`UGI'����Z�XݸG⇹��/t��4�{m>�%�NZ��j��dQ_S�׃��tx��\��4�3$ցDFF	khI+�!��2[ɺ����m�M�Ĝ�?���!��gb�0{���*|}E+����*��L��� &�5�2���&�+�nԍ��۠��.�3�n�a�ȱ*�D����֨�"��q����_�����\���s�������u2�U�,a�= �o��^��R���ϭ����:��e���x�\t����Kl�Uo��������&��j�љ��7Z���E��ѽQ�d_���hU�K7�-_̪��>Gؚ����6�����b���i�����=s'IP�CL)��hF�����Mz��=��|�BZ5�qi��1����au��L�<��ٸ�j�)����d}�:3:r҃p�=!x]�Qa{�4�3"�d4(Ω�$���{��q�@$i��!�5^:���I�N!��ԟ�����QYw�X�v�a�vݘE�UYRv�=I�J�y؆���5��S�3�q���\W� �K%�>��k�[hI,��AZc�c\zn6�����c!9S¿�e�ws~�Y����{h	��W�#U�AO�-�'�|`�"�x�^߻Z�@�+m�c�%c�]�A���G��_2CWcc!�yY��;���nkE�L�������jO=f�1��,Į�@�7/����VI鎮����6<`L�p�`-�;3՝f?��!5r�t��ѓ�������D���u+��:��(��o�i�'�a	���V+bG����Ze��Aݼ���I��^\��;��ZX�[�uw��M�l�Y��R�	�J���I�y�<'����z���
OG�����5�©kt���nj��U�=l�ѵ�'DWi�B�{�p�O{��9ʳ]��\8M���`��F\�����w����D×�T�w/�R�A��8{J�#�ʣϹ��=L���Ȥ�@��>5R��|�/��A���T����m� �h���%�x8��W4��A�n]��$�yǛ�$n5z* :�Ŷ����y������$~��_^�3�B�eh�/	Z�� ��eE�.c{�ћ�:B��7<?@�{оY�|"Q�l�se��F������1h�%��f��,si1mR�Eux"�g8����'2=\}�ߝ�Z2Aq�n����U�;���s��
u��L��,�S��j1�K)�A�K�,j�Є�		���&D�_�"�Af">�x�P흽?^dV����Xmz��A
�OOFe0� "���K��߭C�J���x��0�+TT�	s�*y2�#S-���������M67�YY�9���v�(�w��x�u�5��[DΏ�{��������0����F7#}Z���#��r����D��_p1� ֙��AN�|��3XS�kg�W| ��i��J�ͰY �����IM���g�Tg�a�N�h�B��h�f�����}]��p`3�l�ۿ+�T`���^�`��bW�b�fh�'JZ/�:-���4�e\����}�����%�;[�{�?���� ���:�}���Qa�)�56H��Dr2��vg�Q�߉(����~P�:}�oi�SP�|��t�����4�5��h�E���׉u�#�@B]j*�ڦ�$U�s� ��ǌw�r @	�aTڋK�	iV��a��"����VF��.N>A���8_����y�J.��̈[�Yw��{՛��M�����	�B�N~IF|-@�K�˶�m����z����|�W�c�Ac\{9pB![1<�.D����V��<෇yqo#�QK4���0`V�@O�p=��9u%��Vǅ��&˰VS����#2�q[��@���?K�V��;�y?xd� M�3ܜbJA�§���fK!��c�GU9�)�|���8Y','G���/�����4qm��.�����\��Fi3�q̕�WԨ�V4�]S���e�n��ך���}�W��p���J��g=�u��f-u���#�d����r]�s��VJ�w�@;�Agx�r|�_����Es�]m*�[�_)�|lx��ɹ����p�I��m44rA屡6��?����v٩��l̚H�vS��5������O����۶-�l�ۍ�k7�Z���T�E���X�*^T��ôfU��苙__C��(���J6�y*������.>�D�����㯐�B@F��g 'q�z}'>�I:�eG�&�����"4�4d�0��U,�����ay�(q/t��wnf�{"�YQ&�`��l~��Ѻ꘴w#�ww�x�]:�*�?@R'Q�.� =���[Hl���NC���&K�ɧ�s���QX��IPVk���>ߚ���y)*_���6�JOaPO��CB�p߭�_�r뽹p�5�����*�ˎfj_O�13�+�k��q�]�+��9q����K�Dh)���!�ԅC�������$6����2�W(��9�Nu�{5�Hr7"��#$����'��/�>E����V��C�ۑ���F�����.p#�PU����,�hr%�RȨ�����I��wm�/�j��h줻�N M��mS�&�ew7����Tw�P�vN��F��}�}���~���moe��e��>ΎѾ��R�zƘ����ٱe��O�7\��>4H|�#�����U��E�����H�_�|���y,������>�|SUX�<hJP�d�|�����Hl���/�E���)xZ׉t����'T*��}����ITS���������Ϋ�U�_7¿֊�����u�N8�&��˝p�-0@;�<�A�1_� ʁ�H�@��v<�,2�4�a��H������㙰A�,����-�\�����u�m�����bʸ��3�|Mn� k�ݞ�������<Z׵�c�Uam�Y���{C�^N�	
�09�^(ש罏�6�qu��+a���}o_��怷Ee���Ǐ�:���vP��%&=-C��^{��jݚ97��u��TY[��h9�31�	rSN�,& ��!E�%��`�g��IB7J�r(fX�Y"G�R�_O0��t��߀��qNuy���9?y�S��b�k�;�����Ҧ3�f_��	��b+a�5�m�ɺJ���h,�e�?�bH!eδ�p0VPi�cx}����a��?��F�&�:]խ���9�+岧�D���,䜎�`)�b���H���|U�����{�����_��W^���B�Z|r�*�����Uiξ�8��oH�R����
�}�H��d�X�e%Ox��t-��zּ�pQ�-�E۞�z�a�j�=���7�b�� ����d���C��φ��-�������G3��������U����w�8��=u�P�RL�:��ԓ��Ց]Tǳɋ+��rB��qd���.ǲ*����<b<����u�dm�ů}���b��r��a�X��]5�{z`q�n����J(�t$��6�fq���i��Ջ��^u�>I�{��j��l%���?���QJU��3�1UTJ���@DJ�\����5�+S]`'���M��&� �Z���k���IG��A�+lc7Rk6����!4᛿Q��w.wY���(h�\-W8����-�@����"���^����Z+H,8c�x�������;�0�Cr�!�_���;zg�_���w��}x�@�O���1���)@��/.���=�H)����=#6W����;\�;@=�������� ��Cp��`�lψ�h�N�~�H�F�#�
o7��'�9c	�D�� �">4,�eFLݷ�	m�������\��5�L��u���H�8�v�A��f�eC���	n����z�
���2G6��������zt��������1��=);����W����6��(�M�;�8H����M+sg`|�*\%4~˗�)�*��$���r�S����R"��3�=ߒׅ )����L9�w�O_�?H.����w��/#j��p�P���^m��C4C�Y�%L��8�?�4�Y��)�V���y�Gp����np�$*���Y��(�KZѯo�6�W�$�Cp�:�o�U�Q�,ec��OZ�l�&�E4�cV�<����t��D��M{��Y�'�Q�z�s@��F6W+a�1c��b�y�a��iL���u]x�PgsyR�yS+=W���RM2���n�=[T��;q�0s=X�ե.�G���a�LSe��1���)t1K����ڤ�	����_[��A�y�Ԑ�JP�'�?�)��ZQSm��oó
N:F,��{����K�\��ޟ����<�0[�+ʸ	��[�#.'�ٻݲ5Z�Ჩ���7]Z��Q,�h��(���^zuC�O�V������⧂I��pͫ[u�|�#An4��;��.��1*�ZU�z^��{���"�η�Ԋ��[�f^�W���gG�$��H�� vy(���M4|<�b\gu�K�	,��]�������,5��$]hj3p[�ul��$�zԧ�o,�W��;�l��t�bo+��"�/�l�x-9�O��\0���X$��:��%-ks�v*?%��s����}#��,���d�5��NH���D�,��<���lbA��	����"~�,U:��i�MU���X���4 ���C����N�-H�u����Ej�I��a`Uk�QsoY��4�J ;Xu�����iq�aC7��iˋV�A�ɔA�61ߓ�ᗴ$Syg1P3�6v�w�E�6��M�k*�9��B_^�~dM�-�JK�����r�+���s����cاRA~N19�w�[!�.KW��7����S�o�)Qf]�G�`1MTO$�­G,�%�l���g�{/V!��#6[VQz��'>�:,�̱��;��T�u�cR3������BV��a'��9�oG �)ӭ[�q�84�k'��ǅ`cJ�)џ��o�j�C.�b��r���g��3)��L����ʤ���`����R�j�Aޒ�G��2�Ejg��7J?dH�e�/f�?O���?�]��9�QR�wFHU��Y���5��[��ʂ��5�mŚ��Z��|Ǫ�},��G7��Z�$�'���r�/��14�?�e���2���lG�T�Q���U�=5�S���"�O!���J�އ�#�Jڀ�5�%�EF��X�^`T�`c�o����Ι�������J��fy%$n�-��X"�I�Dg��la��˗��<���1�'�Iz8\A�dde��Ƀ����]N���L0���,���i�?y6@�q�����aNf��"���Q!��l)�'c���s7�����Q�I�W�<�]5����TR�&ÎI&=B��[#���3��_|�F$]*sk
[QsFI��@k���>�%�~'�)% ��c���6%ak�E���p�C�_����T�X5�m��q�7*�Bf6����a3�l$k[���h������R�\KuF�)���!b1C`	�P>��o+v1� �꓾W�j�9s�����H히7]�����;���P��NG>+T�Y��1مC�X{��#`���9���d#�����Ij�C_�Pm�h��D;�wyO�/M���Mf�6 (���9m���`ţ�7���.(�������É<�}BD��y��ȧT�����Y�-�9�-���ӯ�i�F�`�O�?�Vm�Yڑ|~.��j!��W�EG�<���_&�N��k��,
ܝ�XB�^��;4U�b5hEʶd6��� S���<�1�� ��!�UZr���d'�p�8>����T��8еxK�6���J�P��7�X���G�9T6u9��,��P�-��@<^����c�Z_�1�����vw�#2���a����UB!��惙�iz,&���T)���8�F�m�a�H�b�TE�N�M��k�#ڣ��Xm���P������=a��Y9l|{��NՋ�
�)U9�e���U�D�Iq�� �7�cKo���́E`�A�"��:g�]vk�%���C_��{���5������p[X�g9���1I�AS)��&;�� Zc��IXg�ڛI]����X���GX�������p�1rQ�FN��`���S>��������z��3���z&		aOh+<�����=�����c�҇zM�?pV_!2�ô]�01�e�}{����%�HS^�B��&����(�D�܁d+ /�ߦ����՜�%~��'������WI��}�D(���_AqY���z��+���k���U���3�`og���<r����ͭ��n˧��F�e�1�x�rIt`�n�5�1��S빨��y�����jO�`��[7MU�H9���dU�2�!|��M�-����=iG��
�>`4�.�������z���s(�=��P�@]L�z����p� }��z �����"��B��}q_��x�m��Z<ݭ�������)$.	3}����FrH'�s3�]��>{U�������Q�(č�$fi����q�(�i�0�ׇ�^��C�$�I���ŌX�'����mE�,���2���.(UObh��W�JZ_���mQ5�.dS8�s��#� ��J��O�k[W�Ib�AP�cJ�6F���)a`!/�Q�� w��Y�8��\�h���Ws ��w��-cV�2q�"t��^���*+#z�c-!œɽ��Lԋ��C͠!!f���;U`P�s1ʂW������yO���1כĤ�@Z7�/i+΍(D�" �y*~���6r���;{g?����_;�*e�GP��'���y��b�承��Ӕ�Yo�()'���	���L�����gKe�cݲ9�6ҿ���x��������3�u�Y �C��������F(р˺�?�N��蚾7�zL:f���G����^����o�t�w��[�l��=�����?�Wݮ��_�C�G��\*����.-M�fI`wHK\�z��R���E郡�k;�M�"���HR��_�.�@�P��@�f��L�<��Z�m�z�k�ԍŗ/~�+�P���cm��ŋ�Ô��%��E8��47!+��Pt��y�ś���n� *6Y^Y��Li�*;͑:L�$t܌����Y��;7Ke^x��/�Zm5p�5nE��c17�wY��m�O�{~WkY��_Qw��s�'Fq��A�1^�3ϽX-��ig���;�qx���g�=k��\=R�*�S��2�$�n��.Ͼ�;LDqsx'��@���B 伞�S 1��)�@�K�
*?e@�?0D	A���!_}A���JP�т?����N�z���E
	E�FG	���:}oE�K�L��y�T�������E+�_�	�Uo�/#	���~�мL�_�7{�ىB���h(v�ye�uް��Q&;�I��b."�_�&�'�ҭ#|���l��zĔb�J|���l��X���#���q�i��auW2��"�=�q���i Q%��7��Mϊ��]>gе��x��x�ǥ^L��̃��	W�]�EpVm�lA;��5�(���Ǳ�	���8�ر*b
x�_/i	��3���jB�\��0�3�:�u z%ȺC�qm�?_��.���e�}����ӟk�5T�VH���D(����G�����#���~Ɗ:�li����M��M\ܡ���4���I���u(����u�K�hYj��[����U��BsJ�%�=U��Z 6Ǆ�����i�@�a���D��V���d�LA�p���1��o��y����%�w	Ј��|,M�p��2>B��~t-66K�_�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸���r(K!�1�#l����_�)��ToڬrN�'|W�lc4�MS�i��(�gwGJ%
qAڲtva�V`o�,����D��	8ZZ��x7���l~$�aF��'*��[�'KJ#<A��v��c˔7-f�YA��ɓ.�:虖^�T���=$Lt����9?1�Ά�{�b7��\}RND����Q#�kubDIM�o����sM^�6
��	��yRn�.��g�ɓM��]�2���t.ܙBf�-S*�C䉁X�,LÐ�|en=Ph� X�dC䉗O�}� &��A���%ۥ4�xC�	
/��˴���#����.22B�ɹec��`vʌ13<�mh�̘�B�I}j�����Þs���d��%1�0C�	:>���Q��k.���E�}G�B�I8$yhM@�D
�!d��t��r2�B��<'��Տ��6>4�%�?N��B�.wͪ\���.a�X	r���l��B�	(�L�����{.TQ�[�&����d�>�q�(]fpX�	�)(�0�˟|Ex�W-��	D?�Ƽ���!M�n�Z%�Th�5�䐺�M$�I�{������>���[�\u�܈��)F��@!�[}��S�'�<!Gxr�R5h�Ҍ�.G_9
E��Kp�<yg� 2  ��$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Z    �q�5�oN�b�ǐ�o��h�"LO�L)����u8��'���J��T�g�.u��\�z��Ш4�.$�(�!    ���v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   �  �  
    	&   �m�%O8���b���8f��p��'l���4"S
�����?�)O����O��S�0��t	�>=��l(լ��h��m9
OX�����s�f�(w/����e��Px"���}���J)X0i!����&���9���?�J>1+O1�r.I�b�~!R��D������y�#�Z <cEfذ:!�]C&�)�'P6��O��`������2wꕈ|@��_�l2�����$�h�)�gy�ν(-��2��6���dA�y�GA��@)b�E�V�\rWgܴ�y���)b��w	�5!��P��]$�y��M�(ez��k�-��]��J3�Px2�PQ8,�벡Ԁ3�jUQG��>�tuF}r,M�h��uJ0c�8Q�pІ_}��x+����	CX��r&ET�'̐�$�	f��/?D���WBL�P�*�i�k��F�	r5�:D�lp4*T3��Jd�@�S� M�2�-D����D�.�+�Ğ�kt܌�!.&O�PDy�Y �Z��7jчi����'��/�~"%��O�I�Op���>��F�]+�8������@]�<��a̋b���EH�H\��M�W�<�@�e� ra��9Vi��nV�<)F�B�}2���peA�'���J�ƃQ�<aPm�i�(͢���J�Ɩ�7)��'�`"=�B�ǐ09�����9d���!�,�/Du̡�pj��$�O����<�'�?i�O���A��=S����r�E�!ٚp�)��2]�H���A/I�i�R`Q��8�D�w�'�}���S�3�r��0
C�;���bR$��?�s�iD7��O�ʓ�?��}�សrx-Ye�T�zU�$��y�
z��D�1o�x�)���<��':vmB��'��	�g��]w{�S�� a��
���r�)эn�:Ը�����?��E%�`QS�:�$�,-n�e!^�^=�$`ӆT�}ayn�$Ѱ�$��y��٨L���рGOG���",OX�+��'�B\��GO1z����fG$1�LQ׃����I���?���,��T�Q,ސ;������x(<�ዙ�f:~8�A��� Q��	b����$_*O]F�o��b�b�IS��+�hA2_09fKk�aS$`��"���'�P��e�'1O�<9"�s��|�g���_�AKuJ�L≙U��"<�~Rd������2��z}���!��G�I	�����O����b��A��!E���h篁�����A��kX�����Q�p�ݎ~�T탤�"O�5Dy҃��A�x�C'l�t���0fL�$RF���O�ʓ!���S�T�	�L�'�h���$&�z�v&Q(c�(��}b.�%��<����:t����A���qÔ��k�Y��5���.cj��С�IJ)�fG��q0�,�"�|Ǉ��?�}&��
#+��^���SRDRr@Vtqw�*T��'�Q��dq�&��!6D�B�>1�i>�'�`��L,�N�}�6��gm=id��s�i.��'��V��S������5`j����bCL��`�f.���l��=�O֠�&��0r590�1�B��.uh<�s�ڏ1#������t��	x��=�v���S�| �H��ݖs�N`��������!�M����$�OLc��@��B0^��'�M+q��'�"D��Eb�}q
��2����vV8��l��F�'��IPڶ j�4-�xpߴ_JI��e�����&[K�@��U�'N�I؟��	��|��L�:ܚ]��A~�lz���*وT+$�4�?d4Zr
�8����E��I��4@�bܵc)�T�łڠ��z7I���� ��@,iBb�Ê�$K+���'hJ6mv�X�!ďJ
s�4	�G(P�ę� ��_y��'��O���C��ƹ%��L�Q�(�L�k
O
��P,
�xi�g��7 jdHt�ûB�����<i�9�^�c�'���?᯻3�$�ho��N�"D��b!E9��'�"�\7�y�T>�*��p�怦W��В�&4t�h'���&�)�!e��{�̜�36�X���S�iT~OdԱ��'�2��D��$��4r��	�TA@.$�V1�U��5��'���'{��ƨҹ*���y aʹU�D��5Q���� �1/2 !Ǯ\3� ��c����g�u������?�O� ��ـ+Z��Ɋ�L�,'�3�"O,,�g/��#����L���U"O�����'V�J��JX6$	8�w"Op���P,xtk�� ��*"Oܔ*�\;sj���Ò'C�����>���)��'pE����$	�'���ǩOǬ�'��}x�'j�|J~��n�%V��Y҃��l����blB�ɵ4����ۘ#xY���:_nB�	*B�1k�!�D����γj�*B�*H0ၡ�'p}�Q&ϩp�>C��-B�T:pj�Uݶ��W�Xvp�O�E~2���?A��6=�@�v��5J
�S�QTxҒ|����ɤa���ܡ [�}�4��Ou�B�I�q���	��.m����-����B䉙h"b��.O�bY�<N�&B�I<G�~��B��u�E�B�R�\D"B�I#?�	ç.I)�6pK��Q9 ���T�I�l�}"$�T8_�i3u�_�W��%:�g�7B���'a}�,y�� ��k٦	��]Ytk��y�KB�N���>'���F ��y�l�$�T����C:h����� �y@4[+l��S�Ϟ �d�h���p<I��I��:<YD����]3ee0��	�}�0#<ͧ�?1���G�<
������<*�*IQ��S�!�d�*g-t��5/L�Y�:�A#�\�!�!�$�#|Xx�*A��+l�L2�@�9A!�ġ=���c�_�5nbp��o��o'!�$�;���e+�cN��nA��N9���?���̤u��W�W�$?�e�4 4}2@C'H�'�ɧ�.���s�ß�ȁB�1Q��u��;���{�K�*l����2Wø��ȓ]&���V�������/f0i����{�E�8?�̤J�	R|0u��{1VmQ�d�.x-���`U�qX���=�G�ɩB���ձmgN���T�X��ʗ+ZP!X���^�	̟"|�'��a2�׋s�\��2��<~F�@�'�B)��j�>Hf��1�ÿr�F)�'�4	��9ج�k
�w�\1��'���Ù1Hu�6��p�	�'�t��@_�iB�:\}\m �o�R�'��)��)U������^���8�A�_]����؟(��	"
]^�e���Q�Pi��P�VC�ɍ? \��Iȫ,�!�Z�=ӀB�ɼ<���g��	@*֡�5%T2-5B��]��Tk
�.��`�Q�Q���R�'ݢ-q���giz���˛>;z���'�zŰ��4�x���OZ�&��I��NtX[nR{^�}����`��8NH��ڥ��a������T�$�*�$h�#�*t���gĢ�Y6�S�!V(�6g	1� �ȓvM���C|:U��NA�dR��O܉Ez����O���Ĝ�w$<�Id��2��I��}��ퟴ%���|l�]%pi�Q��/y p��"O��#�N�a4��/̳��أc"OĘԈ_�S2���V@�W�Ri��"Ob���E'D�S�G@�d��"O|��ɻ/)�碉�V��d��$�T�'�x���a����:N�a$��	�6���'<�'���Y��F,��\���ѷ&̉Mv��7)D�c�ݩ3=ʬ�e"W;'����F1D�#$�3a�҉!���._p����/D�h9��24k2�a!���j��S��2�`
vmZ��D)��8��ǌԟ�Q�(�g�6�'oȈ�����7���U)�:P8Q��'i�֧� �� �!�\$؍ ��ؾ�4"O�u��Ϗ	?��B"�FN����g"Or�!���l J�*
��}@q"On �f� @6	���V��Y�'}��<�� T(&q~ȣ��\tX%��ɌU?q��J����'�X�H�6�G15�������wG��D�(D����<EB�TN�>�����#D�h��!��V�k�^7���	5�%D�L��]�nܩ�Ѡ��
��*�&&D��B���8*dy*�* �f�BP3�I8}��*�S��`�D���#W���c�I�	Y���OP�Hf��Or��5�����OU�=�歎�E>��(�!��yҢ�?���Iޖ;��@�wgK;�y��ݍs��+Q���n} 7*��y���%5
�r�H�u)z��Aɘ��y�JO6rx�x	��ڷ6~�1tFGĸ'$#?)��՟D3U,ɪ����D�6.< �C4�?iI>	�S����ʔe��8�S���^=�@���Łs�!�DӒkg�,z�X5	 ����F,0�!��_�J��S`��1g�&-ِѨ	�!�E+j%<l��A6A����-�Sԡ�Dʊ��)a�ڹ%���ω��p؂��D�.m)�>U�IM�1v4 k��Gu	��z5�N��?��ΰ>1vÍ������A�x6$�$�	d�<qՆ� V�9s�TZ�
%��e�<����,������Oᮄ���G�<y1,A,6���׉�;g���y�KC8�\ً�ĉ�{�=k�@P�qw�����)o���y}����m}��	e�BQ�`�Q�KS�|�D��y���rˌA�%�պ5����C-� �y2GT����!5�Ԁ$�̪�yRnSIp&��b�"v�\A��
.�y��ÂF
�;�M�6t�ryA7d���I�HO�c�1\�F�
6B��:�h1�Ւ>��[��?a���S�S�j��1B�ҏ8�=�/۱`��B䉕9�Ġ��`ӥa�t��Y�hr�B䉴^D����A2b!˔g�O>�B�ɶo� 1��� #Ԛ!2J��TTB�0":��H��L$���R�үP4➨ҍ��ޫr�bhN<̡��TZHfR�~����!�D�O>�EX��c�Z���h��Dt'���ȓ��LTj	$-�H"`�n40Ʉȓ+�h�9�%u�
�����OVl�ȓl��#�A\�)��ۓ$V�n{Bȇ��-"4Z�U�R��	�+RvHedN.�=�^xD��f#~�n�s'"�v�"h���W?[od���OB���\"t�Jmyb�T���'	J�(S!�D��A9�m�;���ŊI�1q!�dEj�搀�_��+p\�5Q!�d	5�H�`,�,'g�H!B�+K>�xҊ<ʓ�F	�' �*O�,�@�A�8�΍��~o@�Fx�ONB�'���6l�`�Q�sv�1�S'H��B�I&r�� ��F�<?�!�Q*ѧ/�`B��z�� ��L��e��O�� �>B�I�4� �ױ�n�˔�X�Om�C�	:) �$��@�`6 b�3V� �'>�#=��s��0*�9A�lSԘJ��K^�$�}Y�D�O�O�O���P�-��^c����!\�I��:�'��A1�؟P�D�5���Lf�\z	�'(�2Ц�"n�����C��@��'ඐA�o����T�t扣.}�dh�' lBC���r�ؤbO�nG�pr�{BH2�Mc"��	/l�8J5�m��U����|��������?E�,Oe(�kسg��`q n*"_P%"O� $��&ȉ�f]�mKc>J?xe�ȓx��QG		[6�E&M�.0� ��6�$� `��>O+jM�-�9�⭄�R<��IքE"	1��ÌEY�c%� b��G��	�U| �t��J����&Ƃ������O���d?W����c��5��)􌋘R!�D��  ȣUAR��=�I!�$� y/�𘑢�	���%���!�D�*�Q*U�ć(F8�氄]�Ǔ5ZQ������� I�DG
 �8�⭟���%��|���?��O�2��Q'<3Pn�&�cR"O6%q���$+L��sJ�����"ON(� �?ز ;Ui�%W�t��6"O��+p���+��SRۢA�eB"O���Č!C�h5��aG3G�4Qǚ>���)��
d���lv|�Y�� ��w�@�'�Hq�'���|J~ʕBбS8!iF�k�~U1r�ZJ�<����(�=ؒ�W�{��A�gÛC�<A�,
����X�j�D��c�d�<�bb@)PK���F�"&��g�h�<ÁU��fŸ�OO2&(L�6� yܓr둟�ѷ��Oh4+�+ez���q�\5r��Xp0�F��&�\�)�gy�@��l4�r؞Zd<m�b\�yrF�%1*�trO2R�2,qw�V�y⡟�qh�|)�#M�v��s�.�y���<�:�M�:LWjaj��Y��PxoT.�
�_�W��a
Ԝ��F}REϐ�h���д�Q�$�d9a-¹�����X͟��IRX�\q���=f��K�'��A�聠�1D�@Z���7�rue$X'%��9�"D��9)9jl5R������葃%D�����	'��a�s�H�HW�H�O9O�qEy�͏M��+G�� *~5��	 ��~R����O���O���>��l��k#��B0�Ҵf�\����g�<�a䏅/�mbQ��*Uz�rPF�_�<��R^Tض�)EA�B@�X�<���3>0�Uq�ԫ����@kAj�<�	�7cj��D���ˌ�B�l�d�d���Oپ`X%�=6�ɓLV����kJ���d���`��S�)��# ��q,�Z�.�I�,�6K!�D�?W
��#&KU+L�b�� ���A�!�Z*κأ�,���*Ua'Q�,�!�$�v���ƛS���aGF�6CW!���7�X!��]U'��x���p-qO��G~2˃4�?ys��{�(L�p�ʑJInus��������?E�,O�8 eL�(e0C7uZ�X�"O���c@֜?��2���;\d���"O�X[�ƔM��=�㛻fD��
"O�������+�-����1%�ݲ�
O��eG��f��w�N%(���y�Y���O�|B6퓃Vl�5"g�B���p�����D8`��?�	���*#�^8hӤ5�udX�!�f��;��yw�[�f)*�D�ܕiG*Ňȓq��!@m^�:B� �T�#�<��|���2��'���P%ƀ	�l��	;�(O�L@�C�8��MzԌ��{��R��O�9�3�i>I����'���� ӦK��#7�_�t���3	�'^nLB���8��1�f�,ji&h��'x�1#�?�hTH�!(_0^���'�"��(���v�ߞ^�Dԉ
�'��@v�D�<���(R3nꪬ(J��x���)�)AKT���e(�@]s���8
@�W�&|����?�M>%?����Y��l؆��28A�� &&'D�,�e��M^:9B!ς)?����j#D�� h�y"�R�Ā(��P���1"O����5o�<ѩ&�{8���"O>���N�E?(��g�o
����QH�';����7}D*b�ڄJ����D�e��x��'��'��Y�@�0��,Lp`kC��"RQ���!2D�����?}rʤ!$H9Q?n���;D��a�O�50�e���D
u4x��<D��0�#.�����H�,�6)��<����"ل@c�hi���� �i��ipQ���é4�'3(ܱb�ĳ�\�
�$ႄ1��'a��'(<�*bn�6A8�!�c��/=�E��'�,E�3E5Q�6����
�`c�'t�"g-��A,���o	�-W��	�'�Tm�FJ܊2<v�H�@�'���k
Ǔ�Q�к�n��&�!�F�BM��ɐHR�I�6�.b�'�lu���r���?��OZ](��Z�X��U��B3�Q��$"CT����F�3�ZY�|&��sO�_>\�X��K�;Ǆ����Ԙ
��p���X�2�b(�C)D��c?OFq���3'W�P��g@���\;af��h�'>����|�����'�"�2�"A#o���vB�l��1
�'v��f�K,
��p��Z /p0�I����4����>�Gd!��Є�_,FXbe �ҍz��b��qӮp2g�O��D�<1���?٘O6�- w(W-6���`��=@�x�W�ȟD�U�L�-4zR]��o8���䑶N+�����~ˌ� RKR"j4�՚��F� ���nA��x"��MP�0s��ճ`O��G��92wz�	Ο@E{r�dʵ1�pH�ЁJ ~[v�^���'�|q�%߰��ʘ�9��9ˍ{�#v���$�<ٴ�����!������ �P;(�#�I�C�@�<`?j���<���?��O���k�FNv��� ����B��1�zaZ��^�BNO@Cb��D����p��#���Dt3ԅ��#u��\�\�0����C ������9o���$�Op���wCT�C~p�r�O��,�=i��<)�o��z��q�t�"N�piƆ�t(<�N֭e�DI�Hϣ6���$�-d���R����$�n��)n�\y�	O��5�V?#��qA��}q��D�U�Pn2�'$�mI���P��E@�@�*DDl�|*��@��n�:T�6��`3-���X0�x¤��Q6<��fZr =�=§Pft�t�+a�Ij�>�.�'��� �O��D ڧ�M�b�Y"{�R�a��M�t����*!���%�(�S���p�����	��xҡ>�"��c���(fX��ٳ�Vl��s��@���O	��'�	w�l��v��-׎�(Ԩ�QZ4B�ɛg�`0d��>ydi�0g�%`$B�	�]��XЕb[qJ �	��VV�C�Q.j!�v(Ì;��$�!� IRhC�	��>h��Ծd���b�$��DxJ�'6�"=���C߀n&�T��j5�Bh�c��b�
������OR�O�O���[��]�0޴��Я/e�DM �'�ȵ�Ե߮89�
��b��Y�'��Ds�
�u!��#S�:`�<��'�`IA��zF
�KGJ��RC���'Zr��R��=9�Y���>J��{�.>�yT���ɃD����Ȍ�[�X)9J v~�=H�����?E�,O�Y�'��1fT	���T<�h�U"O�%�G��W������� 8B�"O��ä��5(�y����0�E"OH�@���D����K�]x
O��[�(�h�X�R"[�	f|� Wg1��O�{a�/Z,��@
>m�&X�	�!��J��?Q�N���+�3�$ pP�B�L�,ф�j&��ǿYJ��2�<����ȓ��(jbJ�<;�r�a��T��u��R쬝+�,�.j.n���BB;U-��I�(O.Y��k�/��˰���* �m��"O��z�@  �G4���'��ʓ:�Pg�9r�E{5,��D��?��.Kw���$�'��e��сs"<���LG��VL[��' !�V�t��U��Ί�&�D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  5  �  9  !)  "4  ?  J  "U  w`  Tk  �t  �z  ��  ��  �  E�  ��  �  #�  ��  �  ��  ��  f�  ��  ��  G�  ��  ��  �  �  ��  � � # g 4$ �+ 3  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9�ӄZ���1.*��5�����5	��9���ͺ\4X}�]�=B�=a0T��&�U��8�e�� B�=p�>1{����y於m5c��C�I0d�����̈́ -�\����C�	=ڴ���M$k|$�QT� !��C��2G��l���5[p���C�<�u �
�X��/���C�I>0��[3㔶%��}��j�5 d^C�IvQ�ղaɌ#��I��^@�B�	Z̒���Cv=@T��&_<�B�IK�����,�)f����ס(�B�	�3�ztx�G��J��u��/��C�I�	��,��̚0����F&l�C�&	��M� �FU�<yFb�1�����>Y�B�B��Hɐ� )7�T�u�c�<� CR�*�Ny�tb#"t6��d�d�<�&$�{��4 ��N�i4���(�W�<It��o��13aԬ��<K7h�L�<q��Q�-���34D=@����D�N�<�W���=�����E�v��@R�TH�<���$w�t��4^X���
K�<��mM	a��(F�}�nD��a�J����<A�(N5+FI�'J=���L�C�<q�]�+/���B+����At�X�<��'n/,ds$\�X�x��@�^�<!pj��V�r9�!�!h�:��ee�<)�h�=7��j��o�)�a��a�<9�C�<Ϫ}�W,�(6���R娆[�<1��"��ݱ�#�d���S�T�<Q�'�ޠؓP�%P�L��bK�<�qA���a��]�\;t��F�<��� ~v��`΋4�@���DB�<� ͸�dH�j\/{8����-B����>Q�E�FW�A�`���~�0 mN|�<�1T� �Q�.�VE�P�O�<فn=<���&�*�L1�GGK�<�A�Gx(���21q(����[�<� "�X�'�z�r�I�,Fb�	���`��+���O虺�畵 �P��a�^��0b�"On�����#*JpJ��� E;B�)�"O �s��V���p���+�"�["Od��ŎPG}+6
�qZ0a3��x�)�Ӓ4��6o�r���c���0oD#>i����_5bhzKҤ%Z�Ti���
c���	"N���q��2����/.5���hO�>yi�V:*^�`t�K1N��Dsf�(D�hZ���	_`hd��l�v���AKf�G~��.1�����C��]>��f�?e�R��o̓�P�3U�@�]o�r��x�%����.
�P40-ۃTH*���QȢ���q�\I�OJ�І ��
m�ʅ^"W��J$"O���+���09c`[#�iV��t>qB-@Kdb�:�]�@�b-/D�D�W��T��d�S��4�)��/D��� 	^� ���[%�];`��e�B-D� sd�Vr�d*Ĉ5::ta�!l��C�	5R�p�і�	^��XIW���˨B��6/d��ᣊ�6lB�BNآ�ԙ�ȓF�X�f\��2|!'J�"D����	l�'Gt�C�.@6��-�2I�/��h��'�L�AB>o�B<y�/̕*�`x8�'�2� f��/;(��Ke�
�79��'���!���T`����ڪ����'�h�ڔH�?ӈ�Y�fK�Hp�'�F:�×��@����E���'������R<�CH�.��y��'�X���f��e�X�G��w����'����ȋggԍ�$!Η�.�'��1H�$��"Z��H�U�	x!i�'�r%Z��-�4x�Cc��}��a�'�.�1A��jZQ3s��804�'N������.r��43BD5{*(��'<4��W+�-�L�a�۾[c.Iy�'A��io^|R�)��Y>ʬ��'����F�C�Yi�@�*L�܂�'�	&@�k�T85H]�z8��'����ː�bp.(aDMH-	���3�'mf�
�V�/�x)�p\
N�+�'���Q$��2:w���wH�/Gbt	c�'��B�7	�x�xb���g��a��'�u��i��Ok=�!I�0�zI2�'�#���
���pf��QPz(	�'�d��i5r���p-�^�`��'�:]Õ+�m���K���+��d�	�'.̈b��׺g�v="`aR�R���{�'�j�{��I�?��j׃P,LX(�+�'p��	�	Au��[�E�1z
�'� #��˯7Ü��2�8%��	�'���1�)x
�� rB̭Sy��z�'Լ�8`刣m4�����N#�$��'���p��ɉf�j�� F�6�6��'#�4�v�N�+<N�� � �4s�Pa�'�ri�2)*/w��q@�͐&����'��`����*]���7��v��0�'>� ����/� ���4Č!�'FE��oì�$UkSo�	8��q��'��2hJ.h
S��0@�yC
�'պl�u�T�����"h�.&���	�'M�Q��@AL�ܺ$聆i �
�'F�]��IϭLX)��&m���	�'�f\20��2k�$qb��\�hϞx���� �\CO�0&��@��0�Đju"O �n�/�*<#�j�(v���1r"O����A*h[h"�/��R*mq�"O�i�V̖4����V5Oi0�"Ollr4��S�č�d�� ?��a�'p�'2��'QR�'���'5��'~��K���=k@�3��F6Q���'?B�'r�']B�')��'n�'1�Q�N�Jc�8ô�̽k��m�4�'o��'���'��'U��'���'a��	E��7+�1�aL��h��AxU�'���'���'���%��� ��ß�{�O�r�`钥��#}�$:Q�Oԟ��Iɟ���埔��ß��	ܟ��	ڟ8�b|8� u(Tzw� s�ҟT�	ȟ�I�<�	ԟ@��۟(��Пl9�E͹|�RٓТBH�@�Cϟ��I���	ş�����ß���ݟ��G�#jGr�R*�%�ȴ�2�Aҟt�	���I埐�������ޟ\��ԟ�R�տY�
�k��� s���t��� ��Ɵ���ɟ �I��@��ٟ��I�8Ȗ�+9P�������He��"埌�Iퟔ�	ǟL��ٟ��	ڟL��矴�a�!:zb�p0G�� j��������ßT�I˟��	��	֟��	��rqBܜMsب�g�X}�L���ן���͟���şl�Iڟ��I؟d��՟������|+DY BDٛ}�&�ë�ß���ڟP�Iϟ �	����	4�M���?Y�ԋ]�´R��P�d{���� �rK�I�蕧���d�)� �Ͷ�H�C���To��1�n�h�'�D7�(�����D�O,�I C!���JTH& ���O����R67?��O5��)5��ݮg/n�dC�#l�5�qh���'mbX��D��^�e|�4��������pۼS������OB�?5�����v��57
�h2$/S�d@��"L���?q���ybV�b>=��+YԦ9��:�4�@5\^S$c�R�M��y�E�Od�"��4�z���r��SG�@���s�HTu��<aJ>�u���O��9�C�mF�P�'i�,"���p.*�������Or��s�$�'u��S4,ZRp
s��=�:9��O��H&TE�uz��	��?q���O��q֮ 3ܘx`E@�;"�TY���<y+O���s��K�+�:��CH�b��f���hs�O �	����4�%Y%�e�z��BK1T�z�	<O����O���
;X��7M2?�Ok@�I��}�����"����C�P���I>�,O�i�O��$�O�d�O��qB��oHͱ��ߒ}�b�b�N�<�5T������h�	c�S�� #�gȖ j�L�2�F8*��`)������d�OB�D+��ϔ<a�x{���TF�{2�2�X!�̈́�Bj�ʓ"ʬ��5d�O��I>�-O*��'�13�����6'Tjxb��'����?�'޲n�td��b ~6��q���/�?YA�iX�O�}�'|��'~r�L[Kʘ���;T������.]�)B��i���D���)�ן��������%��` �I(�`��C�QA�.�O�d���#rl�&n5N(��l�O����O�ԧ�i��)$��g)ԾKT�{�([2U�q;P�a�Ip�i>��������u�,T/3.�q�.�)z���$,P,#gt�B�'��'�d�'��O��������ڕ��2d��"��I9���O��d�O��'	�ZH�a�`@��� N-_}p��':���?�����S�D�(6f�d�2Ϙ��H@��ne��cs(�0�N�<�'K���`�30�H1y�!�+#!Ju�,�P@�Iڟ���쟴�)�ey�j��11�Z�B`�a��RzI���C;O��1r�6�S^}r�'�6 �ԁֲ!�(M��ժ�:6�'R���LM����l��iȠJ��~BAA��C2u FL�B�T]ǀ�<,O
��d�CR��)��ՄjJ(��L�A��'�R�'N�	�Ѧ��z%�A2C�
 e�d�Z��)j��	ğ$�b>-�"@���L�Rق�́� 5h`c"�6'�ΓHɜ(�@���$�T�'$�	!w��#1!^'l��9窀�
����dE}2�'��'6��A��<����dC3w=d% C��Xn}��'5Ҕ|���&Dx̙�%[�����c�%��dK�%�����dӠ@&?����O�����ن�;JDL`bb�bF���O����O���4�'�?���О:�\a4 ������I�?1�P��'% 7$�i�)�V"ճA��A��h;�|��sGy�<�	ğ���V��qoZV~R��,_����'X�
J��ѼO�t4�Ũ�+0�a�M>�-O��O��O����O���I�#'Fe���]�z���H�<��V���Iҟ�	j�s�0��,g|�Y0�Lф}���*FΜ-����O&��7����5B�>�s���#�Ik�HҪ{i�i2q�P�I���A�Ʃ�<'�$�'$�耵j��5R��hp�K�yPB�y2�'���'������_��r�O@��P6䲰�f��c������'0����=�?��Z�p��ן�I�Bx�q˄�A5>_ҕ@���)E^���Tצ��'y�|x���?�`Й�t��� ��ATn�|��hn����8B�2OT��Oh���O���O��?!��ς�|ysF�Z
'��d{���T�I��H�O�ś��|bB�
��ѕ'�^�ޱcs�ν��'	rZ�8*��ئ1�''��� ��)N�$�"�!�\��Is�)B�~���/R�'���ԟt�I؟D��>�@U��םj���rUA�2�����ϟ��'"���?��?�(���ʔ��*h�A��	6`IB���8q�O��0�)�釘 ��Q ��y����V�P��	GLV�f��-O�靱�?�AB>��Q�`(��C�'d؅�2,��:���O0���O��)�<�U�i�� P�2b�p=#�d�4T@Ü'���'��6M*�ɑ��D�O���-� y0�!� IJ)��g�Ox���!Yx6-7?�%C�$J��S{y2@��ᢼ�Р���#bkӟ�y"^�p����������I�,�O �0qt�\;��H{4��L�PE)�>	��?����<�1��yg�ʍ!g������#<��� 2�r�''ɧ�O��(�Ĳi��$Lz��q1�!h�у�X�_l�� s�J�'��'o�i>��	';�>D��C�+!���4��6�����џ�I埼�'w���?Y��?Q�-Z��BR-Ҡ������'����?���|m��+��C�Co���@\�'��1�'�����J�gR��#6�	�$�~��'J`���*�pu
!EM�Xd�M���'�b�'r�'Y�>1�	�ºi��A�O
���.Y�	���	���$�<qd�it�O�G�H���R���!�S�\����O��A�0��ڴ����/�.����Ef�2��ߎr�@��.@�-�bQ9H?�d�<���?���?!��?��L�`�0�Z�-��,k4�bW�� ��D�{}�^�,�I@�'^�D�`��؄�v�+挘�%�h�3R^���IA�Ş#p��r��66�B��e�ɲS�B(Ią˶"�� )OLM������?���-�d�<�%�*:�|�`A��F,���U��?1��?I���?ͧ��G}�'V P����!(���c��X�'�Z6�%�����O���O��F�H�D��1CԈэ`��ũ5�L=��6�/?	'�2��i0��ߙ��O*bD	�s�+&� �`�/d����ҟP��۟x�	����R c�gHH�U喳!�j��6 ��?I���?�CX�(�'O�6M.�D�G]�q��
� Z�͂ ,�|�O�$�O�I���6m'?�!�[RV��
�ꎵ^��
"儬�XE�u%�O�XCH>�-O���OJ���O<Y��*Ԝ	Xң>;��e���O����<�V�L������Iq����	ca�~ݸ#�����Dd}"�'1��|ʟY���:F �-)XHU1I��_��a��j�B�S��O��O����͸	��@СK�'D�d�83��O���O����O1���:�6���_�	����V�V��wOX��y�'� t����[�O�����i~`�p��Q�`��e�]q����O�	�Ox�,�X�2ƴ?��'Ap@�W�Iw�<3�lV,���a�'����	ٟ\��ԟ��e��g&<�^�qV�R5��퀄˂2Jf��?����?�K~�!��w�а���OjJ�N6B*�Ab�'��O1�N���l�p��%��X�A%�*���h�3Zn�	�e+�@��'��&���'���'[(dAG������cǨ*VdXY�'}��'�W�0��O6���O��E��}��١2� <r7��h�����OV���O�O�@��A�<!w�	�-�#q|�u����d[�<��$m�a̧Exx�	ߟD! ��=tQ��*��L'E)$q�cڟ��I� �Iߟ0E�t�'���r�P�@���
*�p�K��'Aj���_��?�;C7(�s�f�*3t ��^�����?1���?���M�O
19�冫��0�;�����
�Q(� ���_8ΓO"��|���?���?q��7���\G�t���S@49(O~��'&�	۟(�ZqBMj�y`�퍉	*v����h,�	۟L�	M�)擝`�D�2�%��&CT�"�֕zˈL�'sS��*�6!��O��YI>9.O�xs��,G�z��XA�|�� �O��$�O��O�I�<ѕW� ��? �θ#�*�5p�*p#�#��:@��ɇ�M��R��>���?���a@zq���jJ����J�bt�!�M��O(!�d�Y�(���N�7�"A 8a\�m�G�K0`	��O��$�O��D�O��<��<Q��y�V&�?d\	 E�¾L��������	��4���$Qݦ�$�4Ra��8[:$�Y���3��0��c�	����i>a+" �Ц5�'�T�ա�3����O�=\={�%��@
H-��䓄�$�O�d�Op��ώ\"L� ��0P>�(9�-]�_o����O��l��	ş8�Iӟ��O
�� �-S�c�\qÑg��y��OH�'���'�ɧ���02m&��6���m���|,*S��X+p��6�!?ͧg���It�(
6h���)YRI*��~�J����4����)��by2�d��Xs�K�+p���E5`�����2OR�$�O�yo�_����I���Z�g^�a��e�sD΃#GШ0�Ǆʟ��	_��lf~g�mV��SS�� ����A[>d�b�pQ'I�$Tz �2O���?����?���?A����/渒��ϿdD��U9��r�R���I�����~�s�D����CcЃ1I�1�����įT$�?���ŞS8ԉ�ݴ�yb��L����n���
1(���y���n���ɬ��'��i>��	�x���G�DG��!2�@��8��Ɵ��ꟈ�'*���?9���?��������Ƅ�B�&"X!��';R��?�����7�$�E�7MW��@.
���'���@�b	-XKd���#��pK��'](��C�&:���'F�1�,y��'��'P�'s�>a�ɷ ��b-p����ɠ~��H��&���O���¦}�?�;%��l��O�(*��	��:�~�͓�?����?���M[�O��0�p�	ζS��)���ʷ�via�"JSJHAqO>Q)O���Oj�d�O���O�A	ץZ ��	dc�|t)PN�<�vW������d�	{�s�|p�#�)Hm~�h%�5
9Zu���F����O.��*��	[U04�ËV
�a���1*�*�� �F#>L���c`"aڅ�'v��&�h�'6�A�pqJq `���
��q��'LR�'*�����U�l�O����PZR�
y�H-�f�Y����禍�?Q@Y��	Ay2D:+Q攱��>Md�)F��3xq敃�i�I;��%���O`�$?��@�� ��
AF�I�*X��j������ٟ��	ğ��Ix�'[���VI�<4M0��샯'h�@����?!��6��i>a��$�M{K>��i��U�ѡ�a�	F���4���?���|"����M��O�h��Ď:50e�#��?�Pi�%Z�b��'u�'4�	ݟ��	՟d��	.R`˦�<�k%�Z�G
��I����'hZ��?y���?�*��1Ѷ��(Y�}�  	�q�v��"�����O6���OD�O�S`@p��N�Fv��#Z7C��=���=�i`9?ͧNz��d�2��Y a���h� 
3d�Rpc��?���?��Ş���Aڦ)#tϞt�����DD��|��'�66M>����D�Oxm��F�D�V���a��m�!jd��<�e��M��O��+�:��vh�<ف+ٮ ���
Pl�5D8�@��<!(O��D�O���Ol�$�Onʧ-�@M8��<�ҤSI�~�\�R#Y�(�I���IV�s�P����&����	�Ax�"��5bA����?9L>�|24��*�M�'��Xs��CH�*�Ÿ1�,Y��'�8q:�� 韤S�|�U����ѵ�2c���!Jԑ2E�|��XПd��ןH�	{y���>����?i�A��:���!Owl,Rb�F�[�^���ı>9��?qJ>�3-YJ�N��&�";b�����g~2�M.EyJU�W,���OoHA���7y��^ �ܲBoJ�>��<�������'���'�R�s�yc0(�"A�C+A;V����
G�����O����OHl�n�Ӽ�Q��G�! �/�H�tkeg��<����$T�	c6�,?�T��StL�)��R�z��K�ji�̃�]"�\-2J>�,O����O����O����Oش��NΏD]b(��.�:&���D�<�_����ҟ��IO�s���-X�&�Db�.�Tlju�Ƨ���$�O��$+�󩟾�n5sp��<O�Z�HeM�^O�"P3��	�-�h
`�'.�$�`�'���Q��Ń+��zC��Vk�����'���'�����Z����O��$�3&��Ta�!ąQE�#G	�V�d�צ��?IRU����zyb�+ �a�l��� ��rD9a��i
�ɓ*2����O��!&?��&+��p	�0c��Ep"g	�t���Iן8�IΟX�	�L�	z��:��q�5!$%�FCSC�r��ͻ��?1��.�I]yKwӲ�OL1�苄h���z嫃�2���G4���O��4� �3jmӜ�R� �� �e&1C"��\j��8�eșe��$�����4�,���O����:��ROO�h�R�KR���gn*�d�O��N.�	̟���ȟ��OB�5aWFQ5!"�;�I�@|0��O�i�'�"�'mɧ�IS�s�$`�a�-*��B+R�H6UHv��k!�7M;?ͧ]���V�ɰYZ���%o�N���LȿjY������I���)�py"op���!ϕ �B�2 Ńa�z��?OT�D�O�l�M���H��M�9��a&�ߎ}g��a��l�d�Op��0
`��Ӻh���j��<1�@#kAv�k&��!bj���cV�<�.O����O��D�O��D�O˧b�=ywO� ^�J�I�⚲.��Z���IӟD�	p��Sߛ�wm�V
�Z�ty�!�Y�&H��P��Vß�	w�)��-c�Ul��<Qs��B����b�_�A*�����<!��#����Z�Qy��'2��;/|jUn�} c6�DGr�'�R�'����$�<Q�>��`�β.�v�(���"̾>����?	N>����b��	�d���M�A~�)�L-�� e/�{:�O:�����{s�NW�8nɂ5�Ϋ@�p��#�r���'�"�'0��S��x��Ʃ4�:�{��Z�x����Y�LʪOT�2�f�4��r�Q� �WLC��ͫ�4O����O$���F�7�4?����A���3� `p�"�mҲEGMӃ9޾�a�I �$�<ͧ�?Q���?a���?	���"#����:6����)����R}��'R��'��y��]�a)�5�3�>p|2 I�h["V���?����Şg�ڰ2��C�L��	2�1 J@P��Ć�M��O�(q@�
�~��|�V��c���t�\��֗O��D��m���	ӟ,�	ȟ�Cy��>��/�8�i	�ah�Z',�hN�<�;��&���f}��'Q��'e�@+��	�q!����� P;����M')�6���@B�7�Q>����0Q��C���>�[��Q� �
�I�����韔������j�'>�L�PT쁝��ir3 B�#]�����?��/3�i>1�I1�M�J>	ƣމ,��-$W`.��$.֚���?���|�P��M�O���vBUK:(��0��Q4�0"c#m�Nq��'��'��i>%�I���ɠy���Z�EE��pb�o�b-������'*���?���?�(����d�{x�{C�F�P���)�O��D<�)�V��!2��mK�C�<X����%J�k%�W�pz���q�DLy�O�����$x�'?�I��;T� �� ��#v�s��'u��'X����OB��Mӥ+�H��y��Fޞ"���w���<����?�E�i��O�<�':2뀹gQ�mҐ��$1��XA#߱+32�'�@չѱi��i��Ы�?qA�W���!M�
t�b�]_[��bMi��'��'S��'pR�'��S�n�j=g@ʊ"5�(9�/���D{}�R���	E�Sҟ$�������е�(8#������#^��?Y���4�?a�V0O��I�_:_e�3����Z.vE�v>O��CT�ٱ�?��B>�$�<����?���^0˞|��� Q�������?a��?�����~}��'��'E�M����U����N!j��a���o}��'�R�|R��
j��t"��ɂgL�;E�'��d��;�I8E/�	KH1��M�NH(�g��G�*,�D���ĸWZ����OH���Op�$=���I�t�J|p���ȼ�V�?��^�����l�ܴ���y�H$6t�XC�l(�IX2(�yb�'d�'w�, �i��Iu&�pHD�O����'s�x��� bX���@�i�	ay�O[��'���'��ǭvت�q�eRRj$R�f܁Lm剛����O����O��?ͩ�ҀR$m��I��C8���K"��d�O���?��	^�P���Q+)Cv�h'%('�����bӊ�'�@9 ��O?AN>�.O�e�2�ĨE����c��|B��a��O���OH���O�)�<�$T�8�	�pӔ1sDK.cB�q�ę%"������M��̱>���?��({��#�H��X(ȩ��]2 �h�����.�M3�O���'��������d�w�X�+`��[]�!2��X.,1�'���'���'�B�'h�@CQ��Y�!�	�	�B4R��Ot���O��'V�I"�M�K>Q�$�ɬ9ZW�J�ش17�"���?1��|*%Q<�M�OV()$e0f�ZԂ�$� �	�6�R�8}�C�ML��O���|R���?���P9tŀ��R<谰��:2������?�)Os}��'<��'g哐�XѲa^+�����l�+;�	؟�?�O�l�����1rQ ��2,��tA`��"	��mj�%W'�i>����'h�%� 8��d��2�ځqx��q�%@�����O4�d�O$��i�<�q�i�.��Ň���J��cK@�X'x��'G6-#�I/����OP|��_J�����0����W�<a�(��M{�O�E5���"��<QB�Ԓ<�M��B6P i����<�+O���O����O��O&�'+�H9f酩!��hc`�-��U)�Q��IڟX�IL�ڟ�:���%�O>sj�����$�"e�ׄ���?1���S�'>Ř��4�y�O�QC�l15��D���A=X�<�ϓ }�u��O��O>9-O���Oft����<O����9ʎcP(�O���O<�d�<�eY�l�IڟT�	�eP��`��H'��A�3��|�?!�V�x�	ڟ'�H��L#4�l���3_�@�[�`9?�$��/?X�bܴZ�O+|����?Q�͛]��)�E��B���:A@�?����?9���?I����Ob4 
m"����4�@��ԣ�O� �'���2�M��wT %��פ2���#ʑ!�@D�'�"�'<���?�����ra���4$ڭi�B邦�C�@{4G>��&�L�����',R�'�'0�X��(�_A�Y��Cʡ+����WQ����O��$�O�$)�9O�4���
�E������<%��n�Q}b�'|b�|��D����Ccҵ5�P����/v���i������9�7�Oj�O�O*z�)C)1�4u��,	�K8�I��?���?���|�*O8��'��CK�V�~1��]��yv�Z�?r�v��t��O:���Oz���I�rI �
�(~��� ���{���XxӴ�b�n����?�'?����\ԓ���<�(�K� ��B)��	��D����Iş���M�'9Ů䒲��'{|Xa�H�F�!�+O^���o}ʟ��mZ�I v~�*vȅ�D3����*��/��c����yy�+MO�ƛ� �'� �C�G�?(>���P%Ht����A��?у�:�$�<���?��?a��F�+�~��uF��c�J��Ё��?������EK}"�'���'�)i$^�Q"�0N���̊�'dj�Kj��Ο�	o�)���8-����C����aZ�@S�i{*��,>��L��T�P��|��:{;|u�b+��Cn�``���^�b�'���'���dW����4u����'�!nT�١g� %.�Γ��DYܦ�?��W���I�6@Aٱ��+7gzl�(N�B�	֟�����'Yv��Y�'P$9���|?
9$A�*?,=�����O���O���O^�Ĭ|���O����ռ.�l� ���0����O����O���3�9OX�mzޡ$�=��< c`ȼ(DX�r� ꟼ��A�)�Ӈ�f�o�<$��#
$1�4��>8�nR�<9��N���������4����pfH�t/��N�8���H�>���O��$�O �k���ğ\��ğ�c�
�!�qTL�P�ڴX�x��k@�	��Io�%BJ��!'$��h5���C�6�&�2��L�s)ǍG<��|Rc��O����M��=b1�!/���bu螋Lm0m����?����?���h�>��ʑR����F��,����AدD���dp}U��b�4���y�ᝬ]ol���C="�Feh`��8�y��'�B�'L�J�iK���QIH�`�O�v���I�6#�(9��lB�p���봁@[�|y�O���'�R�'}�֜id��'��|��ľ���,��D�O����O�?Qj�FK0C�Lh����H����D�O��D#��):�q#U�N��u����!UD��s�tӊ�+�if����%�0�'��Ёd�R'T�s&c�+|<��'\B�'�����W���O*�Ĉ5g|�C'gF��NU�*�����P���?�#\���IƟ�]�nvV�Qwi!O�^Ydo�>~p�Ѳ�����'��]��[�?u����d�w�xh#�'%(�[��7L_ ��'#��'0r�'��P�b>���+��jqb	�T��Ο���L0�Or�3�V�|�j�;s���i3I��a,a�-����'F�������ʛ6���Z�ܹe��� C��R!p��J�T�&�S�O��O���|���?���c��+D'�0j|�)�E�XlA���?�)Ov�'��I���Oj��	��?'�q�bͤ<*@J�O���'���'
ɧ�	�< �D'�"ư�C5`Q'L�j� ʚ^=��xb���5�R�FV�	K��$8����QJ>���Ĭ�����˟��	�P�)��hy��tӎ$�.I���Y!��%$��P>O����O0-mD�1@��ɟ����| z�"��MN���i����I>x�f�l�C~��^��������߹l��a�u��5X����IޱQ��ĸ<��?��?Q���?i/���b��,�����$��
�m@}R�'#��'��O"��q��́*�!�̆=uI���,��y�Z���Oh�O1��q�fӚ�=|����a �A�td����;�`�I�F@%��O�O���?���c��1�"	�l�fd��j�$X�����?)���?�)O�u�'���'��A�v@���m�0�2��K�O���'�����G��@{��S%<�DQh���Y'�ɧJN�E��XV��Y$?e���'��}�I�|(N��RHS:�M@ei
�5r��Iڟ�����I\�Oj�Ϗt%0@b��\�r�ڑ��	�b�>1��?9P�i�O�.ŌN疴��*'�ns�AN���d�O�ʓR�\Y�ڴ��Ć1<�L��'L�Z�:��L3H�ӥ(�Xh( �<��<)���?����?y��?�0!�[���Q����~��p;4�N2��d_v}2�'��'��O��B<0�:�F�>q�M�a/�p�8��?����S�'t��t!ɏ*_-���6���~�~�x�`϶��h�/O��*�"��?��7�d�<��.
Z�����A�;���tnX��?)��?9���?ͧ���Bz}r�'8���q���br��-�j}���'�&6M �	����OR�Xk�!ÇcE808�D����ѡJ �Mk�OPdx2NW�r�'�i���A�+�-��-C���"�.�$>O`���O��D�O����O��?�Q�N�4��S���y�*��ܟ��	����O�ʓ!�V�|,�#5a� Ǿ
�����ǋ6\��'����D�Ќ]o�V���J��(����ꂋ��Tz��k��b�O^�O
��|"���?��"
ٹ�K=?|pa� P	 ��U��?A+Ob��'���' 2P>��󠖳([���F�K�Z���9?�"]���I��('��b�6�)U�R
%C(��P��%�<�;�m	��2aA1��R~�O)rq�	�%�'����
�+7����j�o��;2�'���'�����O��Ɋ�M+��'7�x���)� x��hL�<Y*OD�o�V�,��I�(��0!X`�J�"�9�4RcΆzy��ɡ3S�����E,�d/HqybG�
Ov�:�Fҳ8�l|���4�y�T�(�I��D����,�	�0�O��y�c�+;Ζ�8��1������>i��?I����<�b��y��.j\�5{�� 1E3�=@��"���'�ɧ�O]��IQ�i��� �����:U̜H�#H���^��v=O^���l��?���%�$�<�'�?y����v���*�X�,�����^��?1���?������h}b�'|��'����`�e]� 邮��U���2��R}��'��O"|���Z0t��ܡ|�t�2����P��o�:}#5EV��n�bğиr�G .u��V�F$c#�T�t��ߟ`�	ܟ �����D�t�'���D�N�f!��OY�.w�\bu�'� ��?���0ɛ��4�l��Ծ#�h��@�E�"|T���9O����OH��Š6-4?)�&����)^*b���V%�#_��A�D�zL��J>q.O��O<���Ob���O��S��X������5h�!򓌾<	Q������(�	~�s���5���VE��&@��~��5B	1��$�O���6��)0d����V[{lٲ!�>$L`	y5�no��-}|����'���&���'�x퉂GQ8 �53�R01��'4��'������V�X�O��s>�ˆO�gW���Fh��Ao�����?�3^������	�B1V��qIF�C�����I6�8;���Ӧ	�'.&�1���?u�}�������3��x�\��
�H	�U͓�?a���?a���?���ON���p,�"B'���-�FX���'���'�����æ�&��K`հ6�vDq���s¬H��(���H�'��ta��iD���T6V��-N�N��- P�(:��*Y,��	�P�Oy2�'G��'mr!۽Sb&h�͙
����N d�'��I4��D�O����O��'cg�ͣ@�$GZ�(x�l�2Eh!�'t���?1���S��-	K_�+�ڙqx��)��TFݒȰ4�N5�6��擏:v�$/�ɮ�ĐH���3|���+����Gy��D�O����Oj��<ɳ�i����W�B�쑪Ǌ+xUb�'�r�']N7M$��)���O�I�R�$~i�ԏM"�(uE�<yu�T!�M��O"U�A��
 ��<�Fo��w^ڵ
*�PInH��l�*]��8 �$_�n��Щ�e�?�r�J�\v�J�(�Lq�QCo�$I����gjѫ��y��៘.���
�`�_䔽�
��T'a}�J_����t*�';�f�f�?|���ī�C�Z鄄GB^�Q�Ď�W��P��(�-'���de�+T��Ud�6J߮���C#��Y*�ᅲr)���l��5'�@�1J��1���a� ^��8�2A)����Q₼f�xBe,�u>��3�e�f;�Ѥ�] R�Nh�I��M���?��?	dV��'[�A����.IZP6`1�SG@7��ͺ�(����~��s�X�B}@�i��[�~.-�Ÿi�'HR�'��	�0�	ɟ��) �p#BZ��������_�Z�m�[�ɧ;U���K|j���?Y�5ܘmI`$*P*�k��]Sjn$�#�ilB�'���ߟ��I՟8&���hm��̫Sp�� Ƌ(=q��-@���K>y���?!������IoJ�`�ͫQ�bE2m�$ú7�I}bX��	a�I���	�]��Tx�#�k��(5-%X�ޜa��	E�	韬��ן'?��'?���Kd��%*|� �J'v6h`l�������h&�����<9��IL?��nr ���@'cY�#��C}�'L2�'L��y�OH"��3R�Z|��jK/V�X���KG�6m�O�O��D�O�e9aN�O��'�bD��-�"p��+�G-	R�`˹��I󟼗'�"]>��	쟠�I<H�.�SቮL_ryy�jô���0H<���?',�������{�6�P��ƞd2ZX����7�f_���Iß,����<�Iޟ���5��@'d���E�,���h��M���?)���!����O��|� �ʸta]�1Ɇ�c*e0ٴ�?i��i���'��'��듵�ĕ���p��f�	^"���C��8@�l�0����I^��Y�'�?9����~���$�1*hu:����j����'2�'����>�(O��ħ�@E�8}�B��D�f�v�J�&�ɝw��'�P��ȟ��I�>�\lE�[W�|���ܛq�d���4�?���+s��]yB�'tɧ5�%�%�Ĥ[�l��1�����섺����[� �O����OP�$$�(�N���B���.<^aQ"���M3�Y���'�R�|��'��� �X��1�*5��$x��� /��|��'�'��OǊ�,}�6�W%� 6h�8'��9�`6�<������?����V���'8��e�E�y`�r�δ-0Y�O^���O���G�S��ħ �����Ɨ4,8̋PHPk���B��i���|�^���ϟ짟����g�J� x{(��/�T[�i���'N�ʟ��K|���?��
@r�D&	�|,��	���@��'�ȕ'OR�'b��yZwP~|�6͈.8��a�B`�#��h��4��$�Om���i�O2�d�Q~2��"7bj	���1�P��P���MS,O����O��&>'?7��pl\LxC�	-:ɰ6���w��	Ο��	��I�䔧�	�G-�,(��W4RaQp ��^.��'@\l���Sצ5��)T%~"��2ǏW2k����imb�'�b�'��)�N�!AJ��&�:����^	q1d�QDn���O6��~Z���~��F��}�F�N�?2��%��8�M����?�/O��O^�O�@XāP��"Q��#v�4�:��|�ɥ9�b���iy��O� � �2@�*7�2D�#gL*QƜ��T�iU�	ڟ���w��?��'n�,���f�ԩp��!/m�a�4:�ܤ�<Y���d�<��O5Fb��0sy����ˀ-I�ߴ�?�����'��V���{ӊ��Ӎ��L��n�,mY|��`�x��'��ly�[>	�ɮ^������ P��O	<��e�ش��'XBZ����$0�dÍ}Wl�3����v�"�ҳ|���'�Q������'�?���C�	V�/��	�g��/f���c����Ŗ'-��'v��'���yZc6��HA�O�2GjԈ���r��Xx�O�ʓ�?����?���?)O�Δ{@h�!�,�%8�dR�Ȫu�v�'��I���"<%>}�W`�;	D���^�Jq�AdO}��DVȦy�	ܟ���џhI<�'�� RaO�@֙R0D\㶍�E�i�B�''��'��J��'�[mr�yQ��9+NT4YU�?|7M�O���O
��Zo�)��'^0q���\���b .J�PF�U�ݴ�?�H>�[?�I�h�I�t�&��6 P	C=���C����M{��?a�P���'U�Q���i�Y
��H3-� Y����0�ܴ(S�n����S�$�<���?!����$��S��F�L�`C+��{a����i�L�����O:˓�?����?A֦�H�ـBc_�	|6-
6Οcy�X��?���?����?�J~r��i�
�ӆ��J�^dI�'Jq�j�.n���d�O4�$�O��$�<���\9��ϧ��Rv$��R�Z5�p��w���P[�P�Iɟ�IFy��'��꧈?Yv�e)8g��2�dځ�Q!vX��4�?)(O��O��dW�v�0}�
w����_��>E���M���?a)O���E�D�'��' (TbT�X%�X��t�_�P��2�J�>	��?��;����9OX���g��-Bv)�T[�} Q�P�o��6M�<��:����'�b�'Ҩ�>��-�L)��KE��k���&N.m�ԟ��� fE����9O��>i9d�W�V��YH���7��t�0�g��$���M�	���	۟�ʯO�˓��T�CP<6��)�)�9N}:|��i��T��O<���O�r����l��o��H��̥e��7�O����Oz�d�~}�_�p�	P?�2��#��@��S?o��R�m����%���#�p���?����?��oY	2#��2��E P\ċV)Ÿ"��V�'��o�>i*O��d�<a��KP&DX��<2Q�Gx�r )�C}��y�S�l����T�}� ��AI��Č�?.be��æ���Onʓ�?�/Ol��O��D�v�>�:���7G���9�B�۶�#�d�O:���O蒟f��'Y6��*fe�1���Z��F�tf`�o�syB�''�����I��d�o�֘�Gf��
�� #�T��&a;�6��O0�d�O��D�<	�6���̟�� 0ഠ��( ,Yp���
,6-�OD��?���?��G�<)����F�ЍU�̽��-�T��	�Ύ���������'O�~���?y��K7����ꑘU�1Q�D2=d��vT�`���<�I(��	ǟ$�'���ǜ����� ��V� �`�	F 39��'YB�'�>7��O0�$�O��������ݨ
"�9j�EP�5ұ*��iE�'��^��'��i>A��� XVHÏ'iL�)��ݥE�(���i��ImӬ��Oh�$�O����O����O���	�;F�!k�IĐ~��m��LT���a���{y�^��3?�'�?�AC/DDYk�+'"�W�;E雖�'b�'�"G�>i(O��$��T�s(��Rd�<�p�;-X�� �>1+O�d�ם�����˟ʂ�Oi��q�h�%Gl�����L��M����?q�X��'~�W��i�y�7��3^�}Ƀ��H�R��u��>��R�<y��?����?9�����$2�)�����,�2r��2�i>듿��O��?!���?٣��
��hՆ��PĐ���,��l����'���'���'��i>�ȝO'��*�-c<�XJd��:e��	޴����O���?i��?�vX�<�U�(Z*YhP��&T��PjBfό#��	͟|��؟�	T�$tӘ���O�h9�������G(	�O�R�Fj�즱�I֟ ��Uy��'�F9ۖT����a꫆�7���)݂%.A�i��'"��'�ge�^�$�O�D�O���T`�F��WBy�bѦ%��Sy�'U|���T�����ܴ+��лw���<�D�ς(�hn^y"�'�6��O����O$�$�B}Zw*�,7��-6x��օ�(�%��4�?���Xn����?A*O`�>qh��o��� `��
�j�"qz�6�$ۦ��I��0��ޟ�S�� ���h0i�o�X-"6Y�5��TX�B��MD'�2�����y��'��`�	!C���ɥ����,�mvӰ���O���OF��'��I����R�Qq@��V�����Yk2q�'��	$?U���|����?��|T~�����&�
�{0a[�N{N��i1��'� 6��O��d�O��D���O�P�o<7�����Ki�*=�X� x��/?��?����?�.O���q�ҹX3*H�'�
����)e��A�>9*OV��<1��?Q�y���OY�,QDE���"{�Y�F�<�*O����O��D+�	��|� &ױw�|��V*�Q˶%̦Ŗ'�B\�����@�Ɉ�
�ɬcK���%��8�*yjD	�\�½c�4�?���?����4��8�O���7� �]"�&^<L�P�;����`O=!�iE�X� �I����8P����~���X"6Y�%�G�7!R0 "ᐼ�M����?+O���l���'��'�b�2.h�N��uK��2'�m��>���?1��)�� ���9Ov�S/u�TI�e�*N�pF��Om.7-�O����O�oϟ��	֟0�	�?���U�0s�W�hn�q+4Ia�0c�Op�D��2��$�O���|�N?�ɰ�
yLb�-��?ުT׋h��������������܉M<�������X#e^�r��Ѹ_Sq�i�����'M�'3�f�d����"=�HIc2�� �M���3�M;���?q���?�1���OL�Ij�^]ʐm_2!"�����E~c�X�v�:�	ğ�����zU�;iݢ�����I�� ����Ms���?����O��OkL�~� S7H�t�fQ�Ї\�k��	�Yl�	Fy��'J��'�W:xU���=���)��6�X�m���?i���䓱?a�e(����*a��e��L@r0�#3�D�<.O
�$�O4�$8���|���GPm<�
���}9K@g}��'E�Y����Ɵ�Ɂ8�z�Ɏ ���W��WX��1ϖ�o���ON�D�OJ�$�d��%�ħq���±$��4Y�I���:@z@�iY��|��'X�i�o�"�>Y�5D�-9���:m��}1���ۦa�	����'B�:���O����5qCdl2-\�h}�Yp�I*{�N�&���ӟ8��!�̟�'���'o��m	�ǣc|���n=L:�nyy��'�^6mJh���'�b�%?��0��薫B�'�hׁO�%�	��`K�ҟ�%�b?5*�a��#`L�y�b�/3�D��i�4��X������<��ޟ�0M<Q��S�tϚ�'�K%�^�8FL�r�i~��3�'��'���$׽c�����4t�4)��(h��!n���������	���'��Od!�Q�F/V�6x�G�ͽj$8h8�i=�'*��r��O��'�����.h�E�˗4�d���6T6��OH��]�Iş�	w�i��q�"�.����hM
M��@����>��(ѵ�?y,O^�d�O���1�td()r�I����=e�|Ec��.�M��x2�'���|"�'��/\���� ��7 J�H�#(������'��I��I��&?�I�O�J���u>]�����B�ȮOv���O��Ot���O��`-���x& \�u,i3��T :�9�>���?��p7�OEJ��s#(֐! Ġ�k�	��	���Ʀ�G{_�8�Iw��E��,huHZInlE��ΐp�ZH�q��R����4��S�(��7/���@����	YO(ə�Td�
���+�2���ro�^�n�+��z}�p�����H6o���`(�{P	��i�r����a�*����N�$l�M�����r�`��ǅ�Bx�a��Wrt ���%�Ȉ�ć7d1a1�AV��J㌋VPD!0��2.��DAuCٙ^�����&��xА|C�jIZ+��I�H� oCZ�)F��8:����AܗB��\P^��d��BB�p�1�@-\T�Ղ���T�a6ĝ�� �ʡg�]m@p�F��@B�6��O��$�O��)�ͨ��Y�M���Q��}m\u��Ğ
�\�uo6L ��G�g��xi��&B�f�6y
O� �j�z�-�z�I�W���W��|���b7��%ʵE֊��D��S(R��+i�O�)&ړ�� ƺ5,�bg� �a����z �I�I�9dԨ�i"��I�6�'7V"=�O��Ƀe�>e�v�_����C`E�S̨p� ��M���?!����Ol��|>�3�HA>V1��tMV�4V"��"��0I�X�	Z��q(��Ux�kU�Y�ML$��X"8�$x��וY3H���#�_3F�C�[x����C֋z�0�$�3F��%�O$���ON�=!��8pN�lA�n!�6����y� �;3
4i�Ui�'c�-X�W��'������":%�']R痯�Z9P G�$DD#�
9!rZ����ͧ~a�l����"�y�W�O
� &�
EAĩ�f��&"��Ӗ�'{��XTė)��l��h��t��F�)~�0!v/;�LCF�3O�=�t�'F^�"��ånJ*��g�fv�6�/�IB��0�p'�)L �J�@7&U݁4
Of�o�:�R�Y2��(�1p oʌX��_yR`Љ2bꓮ?yN~�����xҲ&B0�$۴$ȑu>��;��?���,y$^�)��/3�^�S��^>����]�u8$�W-�-9�lzCk9}�JW�5������!D�ڣ~�"�S�e�J!�`E��:���T�$JH$�'o�>m���B?PwJ�?��ĩ�9ئC䉪:Od�� &R6�$��b�8����Ċy�'��0{S	Fx�R�*�(q��	%H�>����?q��V�|����?q���d�#Re E��MG 5fH���"C:�#�"ޯ��D�4=��#�|RhR�L���ZUو�z0��B	 2��塖*Qv}�fT�#%��}&��I���m�5�g��	����џ$�'"ɫ��|���(^Hn�k��Õh�L�@��s=!��N�EB$HÕe�8�>���X0/�	��HO��wy
� �l���Y�����mM$���
��=�qo�����͟4�'�"�'V���SM��pH��y�ʱ���ʩf@���Љ,�����X)Ԭ;�d7Z��Uؐ�̪W�t��v��C�����1�az"��!j��vj�f�j���l��5�(}#���?���i�V�H�	ZyRV���G�L>.�rX��e�$�@U��>D�H�0����4�&�Sw�.�Pt̓�M�ıi��I�|�n��p�I������BWX@ʰ�@�e
�y�	my�'I�?����������O�u9�'\� ��A�w䆪!2hP`e�'��T�E� �bX�'JL�S��A�R��a�Q�B��IǓ�J��	ɟ��	ҟ�8a�N�`���3v�B�(3j�(�My��'I�O>�/N3�@Ia�.yX����;0!�ā��%�W ĉX("�3���6�6�x��򟘔'��4j��'��'��s��ɠ/�J�����2R���w��X���O�d�9ow�d>�|�'�vUj�B.W1j��R4(��O�(�k4�S�'d�|�إ���0 �b�<i����O�e@&�'���'�2�iI%D�Z� ��D.�����r�yB�'��y��!��M+Ӈ����T"�0<)`�	0Uٴ�A��ǰ5�D�2$�XS�[�O���O<y��1�����O��ı<Q5),m�JR�M@�`�d؛��܂�`�OPi�*��1��'ҜM;ahD�7��t`.�"r^,�#U*T���q�X��v��|Ҭɲ)ܺ@Srf~�0�`���q�B�'e2)fk��,O��W�C���6�\���I���)�@C�	|��c��'�ic����6��[���h�O���S���D�4=��
�H�Qk�m�$���M���?Y����D�O4�du>}��ƴW���[�F�6����G �5ФB�	%`��d�u����]3���hn�i��&�x�u,� ZW�����s�͉V&V	I����;�ObIҭI�U(�lf�ޞ<\y8�"O>6��z.�+�,Լ��	&��C�bx���Ұiw��'p�P��<�^�� l<#/�$���'�����I�|
4���('����1,��è�.d��E��:O>�y�D���2d	�s� lׇ.��x2�ː�?�J>�	>*�����ʛ67]�|딎v�<q�$
h���-�t�L�!�b�o<��ioL�`DJ�:1"E��L�����yBg̺G����?�K~���S�x�i�� l�}[��Z�v������?��#�*�v��I a�@����Ķ��|j���,��)*%���@%�1�O�D� #s�9K7��3=8"-#A�R���P�qǢA�'�f9�b���#��eQ6�>ID�O���7ڧ�?�`�
ȺL�2cOZe�T�sG�R�<y&/��\.���a͓Ŝ�:��V�����٭J��n�<@*�)ʛ=��n�ҟ ��֟g k>�Iʟ���Ty��:F�� S�l��	!VR(�1OX���':ڑ�l�I�Dd���t�z袏{�#Y&��<�	B�v�!%�V�)Z
E<�?q�O�5R�����?����?Q�)�%Q���f�X/|'� 6��x"mԒU̜�1�ON*�teH��H9���@c�����'/�Ɏi�>��T����^ j�Aԫ&��12��*�M����?�����O|�$r>U�ЕU�NAxgA
V5��Щ��
��X$�Yx����T�{?��Y�LD*w�)c�/�/}?���ևEx����'K8���zbϓ�	r��uѝL�^���O��D�O��?!����Qe�iP�#*�4 ��Ӣ�y��@o��0�CO]zm�F��'��6�O��vdu5T?��I�V-�=�6����Ѻ�צ5kĩ��GyR�'��<��CJ�l�"E����B?�cᗞ_ �b�oX>6�r���Oq8�@I���V�@�`O��~rى6�Bj��E)q#�mI��ڣ�p<1��ҟD�	ByrH�/A1�ƪ�<\������Ԙ'��{��CO�~�s�V�M
��1*��x|�ԝ03@�M�b��dB#t���9Oxʓl/���3�i���'�O���#o���Iv)�!Ulac`.D&W1��'���'�1O�3?��-N�s���si��I�ެ�]�	3���?�Km+w�T�qo �EN4ҁ�-}rc� �?Y�y���� .j��3��y;�����^&�y��/G��,����tH��"��C0�0<s�ɲze�-a��D�Y�T�7�B�)� h���F5n1)�҄s��xd"O�=�e[�1�F #�$�r�rK�"O���5&١J	Fܲ�@IhZ(�Y�"O��ag��t�d����.k��(�"O���).X0Ѻ��Y�:d	�"O��Y��
i��84�� �2��a*O ؠ�+A'���$��:GX*��'�Ь�u∍z����S�T�)�T-p�'�y����,oph����o��=��''n��f���Z�,3�e��J�	�'�8��J<��c�b�Y��'�zY���2��'p���'tB`�@�,:���S���i�
��
�'wb�R �,x8�W�Kf�
 ��'���Č�?[D�{w�P�d�:�	�'��M���(�P��w�Z�v�"�'5p�z�яu��U�'B�JF��z�'N"9��_� ؙ�Vìz���'�$�'e �E�\�(�J�wuB��'�n	�w	C^%��`ɾu�ͻ	�'*��'ʐ�7Z���ۂ�A�'R��Q���� ��2����'�&!�CG�6F���'�]�M� tz�'���5唫V�z��4>�qb�'�j<���j7񡢄K
ir��'5D=ɇ��u�b锂s��q�ʓ7��ʂ�H	wK�����|6��ȓ7 �퀑��& �gz�`{�'`$��!�~�(PkA�8kIx���'���� S�bj�{ �5�����'<H!���4�,�ワa�B���'JBXK�n�R.�ٙ��I�z��'�iQ ���,)b�L?��|r�'��͡���� P�L�	�&tZ�'Nf��*�+����Sm
6vf%�
�'�޹v�Ho҄Z&DV�zD�Di
�'GzZt�Z��D��"Mp[��+	�'����GB�pU<<b�	I�aT���'}ĸ��iK0����?l�]¡"Oh�2��"w2a��ֶn����g"O�1c�%: 0q&DΚ4�I�"O(����C�[kR �M��t�&x��"O�]�1M�$뢀`V�;F���g"OZ����0!��KrLE3�N]�U"ORE@�@	:J0�8��m�\ĸg"OΌs��r�$�P�������c�"O��Z�"���	adLZ�d\0�q"O�t���1.�B�2��D�7e0�8�'1δ��ⵟ�bQ�:�1�%d����Zs�#D�X��kN��"hkRi?82�80�!7�7by�"k/�"�J�1aaH�Z$R]�!h�C�Ly�ȓx�ԁ;�� � \Sƫ��=�¹��I�w�)�=E���)��&�׹8&p*���2ys�(�ȓ6P0i�'ҋ)e~�1(]+h0X�u�Nlis�1�O��agLYj���� dyn��e�'���zQ�i���U�P�T��JߛN^�� ��'D�(aF�+Vb9	��݄K>�0(c;D�|��(��3(��	-;-qd�U�:D�� �O�1�4��'Ț/-<���7D�T�q����Pjf˙�\Ys7D�d��9��0,Z2P��dh�l/D���.*[	� 5J����۠�-D�8!���W�����c���#�O,D� (gnHY/�U�@c�I��,�q�%D�� ��8���I�;�8��0�'��RRP��A���)��4�̯hp��h$D���`�N�bq�VK�q��!�`	8�$�,  )1�'K��eW���S��)VI���݆�&��%��`X$n �e�
�y�b�L����"~�n������KL{  :��Z�T��5�ȓapF5r늫,"�\W�I�M0�g0���&�;�O���.�)$޲8�QO�6VP�+��'"v����OA?ye	-{��bԨ�?�Pa���\�<�E���^(IAծ�<Wr�=� �X�'��u��NK�OAH�h�9qj���B��5
��8	�'��ju	Q�BvTx)��&�b��u�[���=E��'�I:G�W��]�VlJ3s�9�'$���M�S*D�y�,�=�(%�M(~]��9�JT�wH2y�׆B2Pay"��'>q�혃e�$W�laK%	_��0<��g�<l$�`bK
	x��V��=?�p�q�Y�=�$�0�N¿kv���k9�t����$���(E2_�hS�J;?�')@� 6Ӣ���N46�1��ן�>)��UF�A�%�m����8D��� ��?z2ܐ��ʕ��p1�BU�Op���#�	-\�j�@b>Yʔ�>)Ba�qX1�ł�	t��`�͔k��|1��1��h���N�yy�tʄ���-�T�4D�ՙ�O\��H�؆AŠ�p<��a�Qi� �w-J6?L�t@Q��U�'׼y��HD�p��|���{�P���'��㥥��t���
�cL$P�F�P(<�Ak�3?s��ga�*�:���I[��8�7�	>�f�P������Ec&?�|r�eP�}��r�Z��dh�eЩ�yb͗�$��5���-96�a�X>GV|�J��H�kX���(cG�8�O؊��kSl�$��s���HBm�2�Iᑦ�X�~ڌB�����j�)��}�� sQv�xC��'x(�0��7�z2m��w�.}��I6=�E�u�A4VN�d�B�>I��?�M�-GQX8c�m�3x$��S�]/*����:w�>t�pm&h�4$��|(<Q7cN��@E������4��@]V}"Zl����IDj���5/['�~���#��h^����3:7�t�I�y"��B$�\"'A��u���p!�� O�#@*�2���+y�y��ęZ�	i�$��!�1;�EX L?�uYSj��f�b.ЮG�6ՋЩ7^��K�֐��;�dC�H*q�IߚDn�5�O��p<�'K�M|F��d.ˁ(c�e���GO�'�6��B��l���ۓi��^������#?�̰q�(Y6RUZ1�a_,Z<��'G♋#�^	�^��D6|�Y�O���3�,��=���X3�$�)E+`�q���(7��?ڬa�];3����"O���ɚ�v���w�ȯ`I�\k�����h�b�09�7-��+�2�>�J�Hhᦞ�Nձ2�z>4u�!��rW�\ v��xK�D���P���2��bD��$h@�R��.e��+�a?=r�Ɗ#mԂ���b�3Q� @�ቃu�h���U���p��_�AC�%���S�΄R��u1�_���$�&( QC�h�-T��0�0�ـT���(��cPi��A)ʤ��*���ɕ��2��'A��|�F��u%���!�d�*4@Z�'�~�I��JײpNvЪF����c�i�Z�X����''���T-I�	}D�ib��ڎoFnq��OT,K�aŦh��!(��Jx����aU�Vm�J�@a���~bc��Lq���dZ�DF��H�(ԕ:iч[Tax2��e�zD���>ݠ6�S!b��a9�fW�HA0�P�U/c^��'m���C�M�XD�6�'t�A���C�!д�[DHX�O�<A�aQ�d��������xJi�?OJUpPĬp$�`!kʔ~M�쩳�$4���P���֬WD�����1+L �R��|��<�c���w��bf�xT��A�V��[�'c����
�G�,x�S�D����M#PW����*���~Zw��yPÒ>�Z�1�O:�� �8�����G�z�~u{P�'�p?�<*W!��C�5�	Ô9;��HG#�<<�t�r�O���eUZ1��S��ӵ��O��ABj�9r 4���-��@�"Q(�|ˇ�Ĳg��`\5�0� �d�P�Q�{�2�"G�
��n�@�,��?9���=���cE�C4`�Ƞhc�ܮCY�	ӷ��.eA��v6���',(}�T>�]�&�:���.Y���١b7Rh�B�C��1��͌u����'�Ȕ���2�@+?9�O��-�j�'���s�掵3=�.O�3�N�NحzC�ձ/�rl2��'-�|��k�����Y� ,I5� 7�x������/B���4�
q!u��I����*Ĺ*�,�?�4D�y��e ��ј������ܓ�h^��]���[�,\�0L>�&Y4��q��-"���d� ��`�M�)��?9�JK��9��A�q��E �#,�U���'�D"��ȼ� c(cG
�2,��*�N�J��Z�'s@9V G�!�\U�s
F�H$�A�ݴ{P���SƘ���@b�iV-7 �Fyr	Ќ;Ю��WΈ�F�A`�aF���>�ҌjAa�_\��C�ȁI��I+J���&�P�M��n��F"=ᥪ^�P��+m�:���4�(�RQ'_	Ë��8@x�O�*x�?1և�<fB pH�S$?���!"��#���a"���>sCޟ~U�����
F(; c��q�����en�ދ>{Z8��j�=To� d�dcQ���3������A��� �.pB2Ϋ~��A��a�y����W�'�����	�I�C�/Z��x�z�BK~����oV���ȕ�wш��#�2���F�C�����,>l�z�N�w+hd{�B؛(D�OPijqI�MaaJ����$ڂ�!@�O�i� C�_�4%��!Z(4����=<���%Z	g�\1��_���ȃ)ݢ�r&��2wc���˓b�z%z6R�D�$E:��R2=���)�G�'� $J�C"O���æɍ %��
)����E`Z\��Q`H<Q��ھ[�t��"B�5�x������O~T�O�H����A�F���n8F7q��ׁ�"�r@��.F��}B��Vրap��l
)i�/�26��-��#�1R󤠟���dI^A���փJ�K�ў,�0��
� �2�ȑ��ŢW$9�O�%YTi\#aφ jsOY�n$lU1�썰h�L��d�vw��
���-�5�A�j� �Ʃ3"E~f��9\	@QK�'	�N��O�Ȱ��ϕBe�4)�i��R�\e@	�'y���%�z�CA��5qfmb�O��9�l*z��7c������Q̎&���E�af�HZ�"O��۠Ě�__��x��@�Z�j�PE�M��I7C5jH�1Jy�3�	�I`�<K!�$^>\|��E�I��C�>uR�16��6��Ij"7!QrB�ɍA��鱀�8
������nw�B�	&vR���G�E����` �ͮ
Z�B�I�?vP����ӌ+��u���'�FC�ɵ_z ��ԈQ�m���BrJN�%T8C��\����a�<8v�"`̟�*��C�ɧ �a��U!it�@䑾q��C�ɫ.�6�Oɭ)bM2�OQkʹC�I	>^l��,��a�Bf�7�C�	nAn��G� 0@����ZC�	AF�=���#I�,�?� E�g�<��I�,'}h}�v!�r��ȉ�i|�<Ye��<l��,)#�C�B��Z$�}�<���C�`�W���9���B�I�Yκa2R��~�v�e���C䉨.��\����\��Ac E�!9`C�[���KF�R�:��HB�Sf�>C�I����BsK�"ʎ!'��8� C䉽�Y2�K�"zvn �9c�,B�I�M���7iߵDNm�ׄ��X��C�-\R:����Ӏ9�����M+v��C�*:����w�3]� [�ʃ)D�C�Ƀ�ʕ �׊t���rb�9U��B�BS>DZbMI�������0&��B�ɢ 8[cJA
�J0c׫]�T@bB�9����<� 2�XzC�I|� eeY9O��A�D6RC�I�%?�`v��q2���n"r�`B�ɀO�6�@�x�کRP��p��B�	�x^&���V)p@�5���(B�	����˄�čzA$A�RA:<�C䉏X*je�5bb��3c�,7Q(ن�H[��!hI�b�N����ܑS�؆ȓ}���a�E.J�[���I%I�<�3�zΜ<y��$�tT�s�Fh�<cś�HZ�{#�N}VDbB��Y�<� ٙ�g	����),z�-q"O�j�������b�Ãg�\;"O�DRlM�vxvQX�F҇`亼��"O������gt�Y1E��(mq"O0��ҮAw�"��k�R�
%"O^�0G�RITɪ�C"u�D��"O�8b�A��)ބ��a�pn��k%"O��;`ƏDl�x[t@��*_���r"O����#��pH E"	�,Fx��"O�TB5nۖl�f�!`�"6�l�%"O<�uG͘2��gE�o� k�"Od��G�)��TC�!�kR)qA"O��j���"U��!��U&"�&��@"Ol��P��9 C"t)kV:s��K�"O�]2�e�6b��L���6sn�e�"O��3��/�l��(�	=�,���"O@<c�J ~�6��w�.�T a"O =A�e0lT����n�^�x�"O����"��j��T����%7p�´"O� �3��)CY�����<>`.tӡ"O���KЙk$8HU�
_Y	c"Or4������je�V�t���"O�顴G�8@DY�f�WW���q�"O��#�n	c�:�s�!*� ���'D�+4�ߔ'L�%IE%<x��'��X�rf�PT��U-H�/�%�'p��(c�A��*/��3
�'f:���_E�cV[�~I�q[�'3� pg��h��U�v�1e�N���'��!tN\f�s$�*},�	�'����PiT7��L�E��Q����'���sk �BQ�5eЈ^���Q�'���zUڀ9-H�/]�T��m �'h���W�����ᓑM_�~PRh��'���L�{�pA��c��
�С�'��]���XU��	!�M��q*�'jR�z��ѻu����'�V�⠀�'�<�/N�zUCG�)v����'Z����	�o�2��-po\�9�'�X��넾��(�k�o�*�:�'<6$����t�&Y�#c�r$L���'nK��!�2���"U��0�S�c�n�<��bUXJ��>X��MC� j�<A� f����f(� ,c�U�Ld�<�#��95@B�Y�����(��ǛK�<!a�%m�^��g�o�BD��H�<#�
�}�z�ie�_��VQ�Q�k�<��3ǖ��נ�*��Itg�k�<�Rf_.a`� �>8�E��{�<����m��	��.���L�<� Ș7����&&Ke걚�N�E�<)t �Bg�8j�
��r�*:�&���|�l�t�bd�h��D�A�%LM�ȓl[}�oƋ[w05���D�-h
F}���81�|(I%��l�����ì4c8B�	�|(�S3�q�682Q��C��`]"�ǿj��,���UG��C�	e�e 0��(��j��}�C�I11z���V�c�܅��+�v��C�ɻ	V�0�ŗ(�������2��B�	�-�E������� ֩Ʒe�B�	0�%�B	=Y>��h�=;u$C�	�DFdA�g�r݂%��g�
S'�C�I�g���2MЁv�@�i ��&A�C�)� �hqe AJf� ��	8+�~�Z�"O���6i�]����qIA#0��y�"OnX8�	8��"JOCL!q�"O�`Y��Hjxp��H�y�E��"O�UQ!����Z��'��d�(�V[��D{��)��3�ex�J�lsΉi��2�!�DǼl�2A��+T�A��2;�!򤔄.qİ)T&ڍAZNa{VH��J�!��9H�9���CcxР�U�V	J1!�Ě�d�~���X�����Fp�!�$H�  �a#J&��J"n{!�$�[���Q�.,�=(F���!�d�;�t%uF�%�b�#7/��@�f4G{���'̴�������m_�8�@�Q�.D� Ȧ��`R���� .p�TM+D�ࡁG
�$&<3⩞8I��=��+D�̰0�����@�0��e	r�@�`'D�x�4c�&e!މ��� D(f�lG�<�g �m<�ź��T�Bv�г��}X�<�O��9"��:SԢ��B&ȶk���*%"O�0��gA@��Z>o-T�3�"OXxp��ۇj.f"5�'����"O �0���8xJ5�W�G�0�A�2"OfẶ �!�.Qk��1#s� T"OP��I�%� �{���WI���"O�mX��\�|0X��I��|�2"O@U���0R��*�$L�"Onɂ%�a$�ջ�ʏ�6��z@"O����?sX*踤
̾Y����e"O2�Z�@
#%��rԩLTu�yA$"O�0+�dW�a��lh���X��"Oz��F㝞o׶�Z�ꏢ]���(�"O+o��]碡ځb���b9�%Ch�<�$#�	@����h�0̞�@u.K�<��/�xք��&� ��F�G�<��̓�t#�=⣇�C�$�i�Z�<�2m�4� ]��f� )�c��{}B�
_��H�0��A��|@r���c����"Ot��Fy��=}��A"O���������Q���8:z���"O@ًîe	��Jb���~I¡�t"Od1�'F�P�T�a����p1����"O�Y�� ɚjrvx"��-a��{�"O�	4)K&.�~���E�C&��"O(���
kb�!��2�"Ou@�A� J�Э@�fD	���1"O�	��d?I��=Zg&��ml<r&"O<9 6��60W�Ɉ��΄t>�Y�"O`|�#�"A~��ŉ��6�TA�%�Im����D?ڦ!q�
<4�yI�+u�!�E�d���H $ �3�B��!�d��]���(�n�x��pQ#�L�!�d	-rU	p��	��պb�K&!�dҧ|�pX2���`����%��i
!�D�\�A��c�����g�	X�!��f4��[���>o�֕XvDɕp!�� >b ���%�`:6�b%d�X�!�fa@�k7��3&�����!��ט��B*�6L����F�[#L�!�Ē�I�.�j�lϖU���a�7H�!�DY�n����P�$�Tpb�oԅ{!�J80 ���p-�(�u� �D�ȓ3�f�8�힓X8�z�"Ӎ rņ�|�I�^6TH�8u��KO���S�? �՚G�2��� �|��eɓ"O�U��o]�""�!�di��LYd"O�mruN���-��(�!{�.���"O�!��݄0/
�8�K�n`B�:�"O(9���x]ʀ�E�!I��S"OhA{���$U>]2r��wGjĪ�"OP��$Fj��P�^�tȈ��"Ov]�b� �>�` B-R�J��56S��
�k�
� D���R�i�F�&:�܀���}pr�
?�:�R�Ӛ�I��"O����#׋�\��b�t
҂��#�S��-H�|��r�ۥ;���to��)�!��zF����W!��a%��{���6�S�O��1�i�!��
���	8�.���'5������+�z�0Í��2J����t'���of�'~%1D�N���0�[5T�r���'D&�i�a/}_4 )c	�h@��'� aBM?Q�( �g�	�8�'7VT�G�E�3}�! �-���t��'�b-a4!ŷ3�" �1y~|���'T��vF�	^�@ĚҪ ���	�'��t)�NA�	�~ �!�Q+��x
�'�81i��p�ы�
 �P�'y�hE.	*d���`h�z�D�
�']蔰���T��`�����l�<�
�'<0��祜a#��!)ܝ/?6L@
�'�N�Y4劢+{8!��*
'4b�s	�'liB*5���:�޺%�]��'O<T��,��b�����$�r�
�'NЈ�D�SÐ����[�+��+	�'l�[����g0*0�䯈�'����	�'�,TA�鏍Qe2��S�E7�DL	�'�R�+B�E k����aä	 ��:�'1�}1��}+VX+r�X�K>nh��'+l\�F����}��k %S����
�'FLha*�4����WIk�P�	�']���CI�$��+�i��!��'�2 �ɟ1��獔�d�t@��'�!Äc��2��	�� ��(�'�4�RPB�3}V!zu�ҁ,��'�H#�
�]V�����ӆr^��k�'Lr�&�l����]����'�L�C஁�pC�Y���"?;�`�'T|@[���"_��QI�$Q1� x+�'N�1��S<��r��,����'�]�`�� f��x��
B16k���'K�I��"��RK�)>0N��' �C�k&��@���?EO�1S�'e�	�eaA��%�M�'my�D.Mq�<��H�%�y�Š\����a��o�<���$S'@q�%��T�ȥE�@�<DnA�8���ʢ�Y���[x�<Ѧ�U�lܹy�NU�6� UHy�<A�oW�9,�r�QwP$[�jQt�<���Z!*\y��IO�'�,�R3�H�<ц�U�?�n����&Y]��XB�<!���-��5R/�<D�49���V�<	��Ղ0�1��-��D�V`���k�<�ᓅT��iV#�1�rͩL�L�<A�� dl�GgǊ�d�y���K�<Q@��n�,iG��?����t��K�<�q"M
UW � �,�-I�L�T�D�<���E�
�QJæA�.X�gkRZ�<�%��3���Z����^�$ J�ϏX�<� P��FB[�f�
�!��I/d2]�%"Ov�zD��U0vb��
�\\.���"O�(b����T���(�4IV �"O�1B苶'ʤ=����8E����"O
����P�͠���yC��xc"O��+ &�W��PsU�E8�=´"O
-���aEH�;� 2��8[�!�ds� �"�d���3ȑw�!���d��BE0k� Š�j��"O���Ҏ��{]�ಗǀ�e�p��"O�!bshs�Q�`�^�[�4�PQ"O ���Q�x�6|9סF
]����"O���$��r)�Kda"��q�"O��F�W��������,�<�v"O&�cř���pWE^���y�"O`�A�K��DNj�`d@K��0�"O(��W��	\�4Y*#���B�����"O����Y J9rHf���|�"OȻ"�ӀQ�؍�����o�bQ�S"Oz,��A�25���P��9���"�"O:�������ը�^�"�0�"O���h��Q��Vf�A
u"O�qaI��0�V�B�[~���"O:uR�	�7;2܁2e�I��Ep�"O���TL�$,6�+�i	8\�z"OL a�U�a�șK��I=58y�B"O�i��fq�p�ҩO�)���w"O� ҅��~���ñf�^"2)�d"O�h���R�h�����(4�j�"OV�P�M�4(�@��&�?`ղ�"On�C��ߺR����������"OV��B�o���eO�"=�c"Oе���P�&�y��(�(�,r�"O5�떋FS$��#��Ăǜ#!�!�1� Yb�M�F~p5J�yU!���T:$�A=N�� hE	*N!�
/|3p�[��D U5�u)t$D�x�!�DYez<��!H��9�D('����!�D�=T���'��6t���⃕Y!�$[9�X�J���	sq���6�ƌv !�D�SX)�If2���֦ӻR!��U�'�h4��I߄y��x;�+-[&!�d�%;��1�g��;~������
<0h!�$N��ެ�c�B$�����0p]!�$չOw�iS��Hlt�	�C��.!h!��S	5ՂP�viH��4��#.�!�$C'c��(A�(ޣGN�q��"�!�Յn�@{�F�S/��y2���-�!�$�;{��&�K�>q&��bㅈy!�O�8�L���'�yi�$���^n!��)B�nL�\�wyX]ؑ�ٷl!�$T��(�����f(QP�K�!�^/+dV���n�a0��I�� C�	x*�Zw�A���)�/ɘ8@C�I�Bs�)�� �-	��{$Z&a�C�I�8(�� �@��$Ȱu��W
��B�	�O��ePdA�1~�Ƞ�C�(#xB�I0x� �@c���~� �1�A8S�HB�ɨS������$=��uk��!�$B�	*���'�<��is0���sB�I��T=��o��@�CNŸ6�B�*P_D 0��ERf�sI�ΚC��5?�<X�j��V[���@�*G@pC�	&2,�W�B��	#���o��C�)� 4�T)��)�DѲ�\&K&`�ha"OFD�$3da0e3�H��{21!�"O�A�2O�5KO.
B�6+@t��""O8\PħI-Q��Mڳ�R 	@B"OԔ �\$oze1q�)X���"O�6��11hňa�F5"��iq"Ot� �&ʒs�h��EC�7����"Oh��'+;P�ٚ�DL�0	�3�"O,�z��̬w�\�ף��c�V�K�"O̘�(\�2���4$ͦ�lu �"Oȭr�o\�x&	K�Ψs�`|`�"Ol�%�X�c���9rO@�}���R"O����g0LӴ������{�"OT�ZScQ11&kK9>�8dP%"Oƭ��m�#uZ�@�����[�y2�]$�<MI �ɰQ&\�X��	�y��A`z��S`� f���"a� �yR������4�2p}����^��yB/�O�.��Sc�37��� �_��y���<x�Ș�C�[Ē�S3�Ă�y��/O`<h�+�I9Br�OG��y�`P�
H��;�jF�L
��bD���yB�5#�(�@#�ўp�BhC&���yd�0x�����!ih���y��]9&����S�K|�=��B�yr-�1 �I'`t��L�y�G̽To�� 7EO�24
|TW��y�m'V44��Tʸ)v����y�,(��	y�
�, ώ����y2'J��l���V'e2��#��*�yb$�N!����S��(��Ĉ�yϘ|��!1��I�ѲR)8�y�J�ks�pb�-Ҵ@���AI��y�Ţ/��d;2Iݎ(^}s�(�y����!锹	��5�L��'��y���g*�U���,^���P��5�PyR��TQ��nΪc�Ac��X�<)�)��j���F�=X\�@3� OW�<���&u�5�S���\�����$�W�<y��r8$<�e�ߛl>�e#�i}�<��C�Q��]�#�-|�L1C#��C�<�c�Q���b�m�(l�J�Fz�<q�g��l�;a �	�Le�7�Cy�<A�'��G		6�EҴ�;��y�<Q`�2Md�|b ��t_��+�O�P�<�T��70�d(s�� [)��8 6B�ɺ����tOC�BM�\��5%n2B�	�T  � ̊�-t!���t;B�	�vW,��׍3(��a"qƤB�I��vx�J��/����nu��C�I�35vai����Z�4�c���B䉵����@�>�B���dM8w�B�	�*Vz-���I�'���`��Q4�B�	�$ܖ��A̳�L�Xq� $�B�;J�@����I�=�"h�����Dj�B�	X	l�{���d�[׀�(QN�B�	 Zv� c<�������C�<aZ%�v�;mA�m�DM���B��"�X�H�R>^a�]�
L�C� H��#�]�ux��k���-{fC�I�]��@�U�r}ҙ�lطH��B�	�`0�0��%����f�.HEBB�Ʌ(8��	�(�܌[�',dHB�	�~�d)���"Gָ�6��(1	�C�)� I�p#QA��(_-�䍛�"O�9ە CY �C�fƟ;����"O^����A�\�8�c@�a��;C"O��XT�Îu��a��(@�P[��qa"O�@Pc�\�t�d���v^=��"O�`�H����H�1N��s%"Oֹ���R�jI�-���E���"O$M�ʉ$ ���ԈY�ni����"O�d�rHJ�p��r'�7�b�D'�S��(K���c"	,a|e�H�.b!� o����FP
M�4��(@�M!��
������Zڦ���۟8H!�d�%~�Q!&��Z$Y�Ǒ2)!�F�S0]�r��/Tp��GD=~!��Z�_
����cѺH�
mC����!�$Ky�~M0�	�#�t�9ƭ[��!��K"1�h�! �ٵw�!�gȩ1�!� D,�c���x{t�qTA]��O���ĉ����v�6IpL1����vk!�O�4�v<�g��'B�0	Hw#]�nL!�΅�L	�E� T�M��Ꮗc:!�*7��PFaH.:�H)  8WHO��4-$7�4�@�_��`�"OP``���&P)��q,���"O&����2fX+w!�:N���"OV�aǪ٥c.��#�/�>!:^���"O�٩����lH~u a�  :5�"O�-Q��@�F�� �7���By[0"O>es��L,U��!T;_����B"O�ey��ˋ:(*�@7� =�t}���'�ў"~����(����d�t��QR���>�O��ä�'���g��/a�x��"O��a��M`DiWnW �F��"O蝁sA�?
l���.K���@�P"OB0�ѵ+܀V��%�����"O��1�Ϝ�� �MҬ,�6`gOf���'�4�]���K)@�a  +D��Q2ķ��Ty5�գ%L��[�%D��x�
�$n��Yc��yQ�BD�"D�,ȅ�*%�>5" �<+f�P��&D��p�i�jxM�S��5)�`�Q/D�@Д����3,c�l��1K,D�P٤�Ȕ�^�b�QsTT��&4��� hF/���� �.EB�50�L�^yB��`�'E�*0�������l}8h��
�'>%0����J���Uf��e������hO?�@���x��Qd�!bU2�ʰ�Gv�<@Ε3'���14HG�>��UB��t�<�#T���i
�z��H�"Y)�!���0K���2�1p�T ��o�4/�ў,�?�͟"���n��;,�;2�э�4�[`"OI ���=L�$ ��,��UbU"O�v'ŧ~L`�Z�풪a�0��g�d0LO�9`Ҡ�9�꽲�Ln|f�@�"Ob<����^_Z�*T�LC�q�"O�I(�	�| �`�I=y5���"O��{���]�*�V�P�ֱ�'"Oj*���U	�#DE�ع�`"O�Xp�_	5�`]� ��(|
B�'X�$лk�|��2͛�<�6��-��'fў�>IP�H�7i˴h�bm
�{�ę��
;D��r@%@�0\�f%�����AE�7D���$'432��3E"���F7D�ѦA�|$����L�Y�0���A5D�� ��"ș�mi ���� H���!��|��'{Đs ��>�p����0ԙ�'�g�^0Z�P�m5zaX��
�'�`�"�e�
!�5 �K7Z�P�X�'��¥�4?��pFF!U����
�' b)Ѷ��ERAR���S�ɸ�'���c��5�M���Q�a�X���'e�x�#��'D`Q���.�h�3	�'�=�w�p��ɀd`�. ߒ�Y�'T��	��S�|3�XԡU����{��D+���
 :Axl�A�_e4��E"O,�8��\ f����
2�a�"O�X�"�"B���0A(p�؉"O�պ�B�m�� ��.�Խ�1�	X>�y���K��!B�y�pQ�"D��dHG#f3\�2���/<���K#��0<�fǂt�"CqdW Sn�R�B�'B�'-1�@����W��I�0+��z���x"OD�(��$�\-3`˝�x��Iy�"O���j'��d��0Xx�b�"O����S�k�N��*�L:	R�"O�Ũ�J�A"fq��1I6 �r�'�IU~ҥ�&����f�+�x�)禅��y�皤qLdPz#��|9��+V;�y�MO !�vA#L��Q�F�yR�B�;7�7[��J����y2�Zy��bB 2�`%���y�(�Z�x#��2��X���/��=��y�ѷ]SRi� ��v.䈀ʘ�y��'�N��ƣ�0v�����4���'thA���JQ��U��m�6F!��'�`���C�"�xqx��ځA粬��'�R ����x>��3@	�=� �I�'?�IW��l\p��#&	.���'������D�5j@p���-GD�C���'6�,�F@�DD8�D�t��
�'%�K0iS�bQ.0ɥJ� P�'s�])�[�d����t<4�
�'Af�I�,^	*�t��d��w'>H
�'1D�k�hY�g~2���W��<�(	�'��3�D01��)0�Ϋv�rMQ�'��p�gi�7Fܹ6�s����	�'q�h�s%͢o�>4����}.���	�'���E��|Q(�!7Bq4Q��$7���|*r�T�S7��jÆ
&)�!
E�H�<�D(%h���`ª͹4U(��R|�<AC.Ӳls\�����K���l�<y�C��5����'�#�4���R�<ͨ �2]���W,�� ��V�<)��O�3-N��'
?l���Q�Zџ4D{����ʤ��
����� "��*�?���igL��zԁ�@�&@�u"�PD�O��D"�g?�� F\�4J��Vrb�l�<!QLQ��s��!H5*��`�<)(3~�\y�s��1v(�@�<�'k�sKA����H�Rԡ1��<�gm��^��Lz�#ȕsҸE�C�w�<駦��aX��k�d�)H1��w�<9�c�>qZ:|��N�\�BU��e�g�<qWe�/���r�%B�\���2g�<I����ǭC J@h�d�ˮrU��Q�z���
H���`��yԌ��l
b��0���Q�� dH�$UЅ�Iٟ��'��%��/��E.�t��:Kp=3��� :	aӈK"2gN��B�]>�T�"O�d2�.�z���(�?��t��"O`�󈅬^�@
��F�'y�l�"O��#	qox��1h0�A"O-A1���h)�*]-��{�"O�|�'�+���kg�S�)t����'�!��5}m�d@SF�X��u�P�ʛAJ!���E�JPq�i']ج����tߡ�$�#ZQ[s����>L$��<#��C�I�Z-�!�OV����
Ɔ��C���Pq&�:�* �0,�3$�C�I�$�M�R����X� ÆEnC�	I��:#��f���6���|�O����8��H�È4I�`p�� 05Y!���'��9CT�X�p�h��OE�eO�Ih��(�����L'D���j�@&O�Z�����<LO6�˒�n{^�B$�H�@q��3w"Or��OZ�=�y��ܝo�T�u"Oh1Q����\LZ�䒱<R����"O|q�.ҕ�����A�j�vș��|R�)J��4�Ì�BUR�����8j�B�	�"sZТ�_�k�����ɜ>(+rB�	>=�j��̴f��p����1��N�b ��®&'𜸋g�T�j !���fV�����<G�6(���L�!�D˘u��ʲ"[�6-�{�j/2!�d��T�8��o	�"�&iC�]�}��'�d�>n����޴h����,!�	$*�b3��K�e��}b����񄚦*��*�$��`�|���L>q��$5?��H�$�]�%�Y/=l��D��h�<�1dZ�@����F�ͳg�>��wɐb�<a
�5��J
��$8��`�bx�xExR��P����@��|u$\;voT���=����dU	^��0�F���YHpL�3�!�]�8u(ffE�'t�	˵J�F�!��?G���iC���qH�J��ވB9�'ga|BLѯB�v����Ϛ �-91�@��y"H�f5ld��[6%�<�@�
��y���3��d�,G��a��X�y�n˥���s���2O^�[wn���y�D�c,-��]�1^��ڶ���yBl��"Ӏ�����?��}�����yrc�	!!���զ��aٔzSjT��y�/��v��!݂Zl��Qm·�y�F#�8���WЌxA�G��y2��A�,|��h֧~;���p≍�yҩ�/@��5��bZ�K_0պ7�ճ��>��O\m'Û�%b(�uF��ܒ��"O@yt�_���)C,.�P��"O� �� ^�6W�s4�uZ��"OlY�6h�`��a�Q6f�ۆ"OF����P�ri���r蔇} "q�"O��À	H?a��d�h�P���"O@E���h���y���:|�����'���(�CD޴z�T �W#��]���#?D���Ϋ_/�ݓ��3�R壧+?D����T�X����w���`�8D��2d���j�A�-)I�xQ�8T�P��f[�{ErD�"#C'e^4��"O��rg�V'�Dܹ��5\J R�"O�U���1.x���$h�jdR�"O������>��M�Y�.4�P"O�T�A�3?$Ph�'ݐ	ɾ���"O� 4@�+M�y�E�A(SH-Qq"Ox5`ㄆ�c���r C0D�Yu"O,�(%Ȧ.��, ඉ�"O��'^#*��ؘ#��B�p�P�"O$�����'�(�{�����l��'�ў"~�f��>@C�tp��w>T���� �y��
���4C6��X���c�h�)�y��A�	Q(�Qb ����n�"�y��N���0�V)I6�指�yҦ��uO�hP��GeH���,��y��\?�����<Jk�9C��ֶ���hOq�R|��."�>d�$�#�|��|�)����0�G�M�E�񏃈K�C�	�U6�̛��mFp���0��C�	�j�p�W�(ٲ��qU ��$�hD{��4_��(�%��L���ɤB[!�y2�ɭ����F 9�]7JT�y��?�l*�)փ2ü��&c��ybdΘ_� ���n�75��	�DF����0>�K�{J��B-׆<��Rr$	^�<-=N��膕*h�m�`Dl�B䉠n�Q�mٮy���;E����lC�I�G{pArv�|�Y!!bK��5D��c o�*K��3�N���d��/D��3��G�6����-�J.��
8D���-�m#F<��MӸxeL-qi7D��b��O�h���#��<a�i�	7D����M5LEp� ���e����6��9�S�'n�$�� ޘU�Ll[���;MZrm��k�.U��j�<F�����Y:F�|a�ȓ&}f9�����1p��/���ȓ~�Z!q�v0A����!�ȓ_y%Y��;p����U:΀хȓ*�.Hۦ(^fɈ�0Vm�	U:� �ȓw���N�.d<@�N�0w%�1��Ig�'�b��W ���
�y��׿`�6�эr�)��NR�,�-B	`ltD������yg�,�d��U���\1dapuj  �yT�i(����� \�0�$+���y��E&D8C�ֽ F䠣��y��>Hv$�v͘�s���It�V��y��"k�4lc��T*r1���C$�?��?�'��0��1F��ЖN�)z���
�'@�|A@áԨ�5a��J��b
�'Me��l��.��աd�	�+��ؙ	�'�fpy6d�#E?�\kc��&�~�2���yR�Ո~U���Dͷ�sp��yBa 8#8q���A���1�B��(�yR퍮0T��L���B����Չ�yrh�1�*����`�abܒ�yR��M�i��㍭ќ����y�d��^$�e��	���`j��Y��y��0M����GF*��ѵ���y���`�㴥F�Db2���F��y2]�x��0atJڅE���悿�y��ا&�HHB1Ƃ16d�z��Y2�yb��;UHA��L�+{^�ۇ`Τ��'�az���M�p�j 
Y�4R�r�E��y")^�mq2Ĉ�e"���.E��y>AF�d� b8�$�rfZ��yr�	&5��-� d
��
�m�0�?�
�'Qu�u�ΰ�B�'��ap*y��'H0Ex ���R�P�/��^��J>����)B�?N|�e(_:>A�`e�!IJ!�� ڔ�a§�̨����}��5��"O�q�ԁN%0���C۰s����S"O�1X!�^"�,P�C�X*r���"O���e��x�言d�<6�؉A"O�PÂ&�,H�L�HƆU�Q��5Hp"O�4����E񲁐UF@�x�d��G��5�S�i[�J 9���, O�����%ў��ӣe�B�8�
�*tШ��R�B�	�:����o.r���GߨE8B��%q9�y���
�%�Z4��F�&�T��p�d@���?\?X�)E�Đ*G�!i�I7D��sV�.�92c�ě�b5�V`)D��c�Q�$dM�@X�$U��+3D��� ��GD�uK��U���q��2D�p�4�B<ʥ�����U�!Z�!�G�}V*� 3H�4l�ܐ��̦_~!��8G_�� �$�(����	3?~��W��(� 1��U2�!�Ɗ�X��5��V������\d]�lP�VP�ɨ��'p�B�I�9�$:�/ͫU��eH��X�a^����;�	&8w����5d���Α�Z��B��;r�\9��(ܾ�i
�.�4:�B��=Y�b)�W��?L:h�Zv	��4�xB�%�ti@ulϲ
$ 3f�ږS�\B�I�j'v�P E[q�މJ"���2����0� �0D
)�|A���/澸8�&!D��X�P�Czԙf�la�b=D�T8t@�Yb<I�Î�.�@�aF¹<1��品e ����F4�����g^�-�bC��;R�b�ҀfQ��a{��ې[ؖB�I8�~ۤ�*O��C1���A�:B䉴` ���Q&�#�V�Q�#Y2o��C�	�J�qS�)_##޹{�n~!��E��L�
"bX e���y���:Ro!�$ŉoR��RN_/(�$��UFPP!��	�G���r,��-�����sI!�dX�O�N8�&Ĝ�gl�뵌A]P!��۽5�f�ь=���,��7�!�d��&Ut��㌋b�H|q��;m�Ib��Թ��Ӏ�i���.0�u��H8D�t�E0�n��C�����Sk*D��`w�Y�
��'�&�|\�!�Ą�ZeƉ	��
�@��Y���\/!U!�䍆iy2)C�����c�m��LO!����y���
�Jp0�W��$E!�$ȃ*!ؠ�'Xh����N�4C!�ׇm�U����jNP|zw�d8!��Q� mf̓�瀻_�Z�	'�^�!򤏙l�]��If�x��!��2!��$?�Z�L��)��#�]�I!�$�$�Z�{�Fz���:1!�dv�%Ac��P���S0�Z�`�}"[��be�3g6`�%��{���"O4{�*Մd�t��̶
\�m"O��.�p�ƀs��P�:�j��%�'���G!8e: Fۍ#�x@
�+Kw�B�	�:�X�0@		�_��'�W2zZB�	�tR�
�N\ @K�o�B�!�B��C��c���υ>n�C�	�\򰱓W�����A2��H4{:ڣ=��'i(�\� -"�SM��z�,�����X�A	BGڔ�Q�f��=K �kc��FR�3(�7'8���ȓ'� 
pd@8��u��%^(9o�U��S�? �\*(2k�j�"Ŏ�Z��Q��"O2��
U���H�MB*T��K�"OD����D�m�4X0��:QE<���"OLUPO�O�r0#F-U$:�}R "O�ISU ��w����V��!94�#3"O��ӣ�NW�t��,ڰA(�B�"O�� ��K���ӱf�n=2C"O6�0�gpvl���L�'N�ų"OP�Y���)>�dyT�6QO�SS�'S�D� hIC$	a>p�rH!�F�CcҘ��j��#��Т�"Ot����,�����*�9_�J�"OP؋T)��F�qK#fP��b�"O�zdIM�J!��0�F�X>�|S�"O �sǤ�}�N��P��t��$]�!�d�e�t�����&|kl�
@�9u���i>Gx2K�+ Z=b��
*�V�Ӕ�]��hO����O8lآ��g%�8';�ȑ�ОO!�dD�J�t�����(�
Xb�&��!�$�>n\��8�@��$�~u��ܢ\�!��(E&�*���@M�����9s�!��$�d 8�	�7(�k�e}�!�)L����5
Ր���A!�D	�2��0���&�X�bξ!2!�Dδ2�4@b	t��D)�?'!�d_�[T��!DK,J���Ƅ��!���Lʄ��B2>$���ϒK!�D�5<�(�taʿ&h�w��!��� 
�(D�aHU�D�ґ// "!򤉟T-^��G,PK�Z�+²@!�ЁG���%KY"�r끋_!�*h��İˀC��#a�^!�䁌_���N�5����E-7Z!�D�ӊ4A���\6�I(�e��T'!�d 8u������X)�,1��x�!�Ě�N�蠛a쁛9B�3R�^�!�!��ڗg~=8�C�,0�y��,�J�!�$K=6��4�be�0v��!ֻJ!��$l��UW���i+��c��Ӏ!���@o���ȃ�/+
��%!��\-t������(�L��"�4x�!��sj��!���++��a�� �~�!�5��
��t��e�I�B�B�I ;	��3���8M��E;qG��mvC�	2����/�&J\v�STlۖ�NC�	�R�� 頩-�Z�2���9:C�ɶY�hY����d���,F��B�	++����fA
���ÔCQ�
q�B�	?a� I�-	Kx��%@�;�ZB�I� j��cc�ɬe�nH�q�B3�B�ɦA��A��4f�|���)���FB��3]�=�˒�Py$)D�B#X��B�	�+ӌ|S�K-a�3�L�:��B�I0�H�5� �^�|h�
]�M.vB�FX�	��H�ĢF�ݴ_�6B�Ʌ=DJX � O�˾�	0.]�(:�B�I�u�|�gi�"H�Eΐ���B�I'SfR��B`ߤ�x�����K��B�	�!)H i D	T{1�J ߖB��1��,;W+�������1vB�I�^���33M�4nm� `�!5/PB䉩0qj�B )�R��z-˺JmB䉫7т�ɗ���8��u�h��B�	[�.���IY�s�)21&�y
� Πp� o���a,Q���{�"O>��@.T�hz�Ś�L��O��
�"O8��&j���f@&aF5]L�"Oȭ���"h���[⏋�.��q�A"Of��ʇO9��H�.�;k�>�PE"O
�C��yc*HR�K�K����"O�=��n��k��++Q�ah��@"O�D2��6�b�D�ROj��r"O ��F��"������H����"OB!r
4�@-���Jl9�͑2"O��K��^�l���� �D��"O��񄆍�<�Vp0 \Ϻ�!g"O>�{�e��B\��@�9b�� �2"OqI�2����0�;� �`r"Oڤ�f�K�Bc{�����.��!�$O56F!)��s��8��c� v!�$[?<��e���O#"L%��B��oo!�$�%;J��%/��0c,ĪU!�䃞9��I#E��l��q�A�f?!�ă�l�Lm��E��k���;��&"!�D��`0ֱ�ʋ颅�@IJ(!�d�~ޤ=��nV�1�IX�	��Uy!����s�Z��sJ�k�`�i��?np!򤔊���Ce"�h���'68_!�B�][�LS�`�\��A��^�!�G�9�x@J��,���ӤS�.�!�D�,�j�����qB�����!�I�x�Z8�S�vc$%[�G�@�!��UB���IJ*���'��	}!�Ḏ"�	c��Ěe�~"gf�2!�`��FH� 93V�Z媘6W
!�$�OL�iU��21|P %�@!�dH`�X@qP)ݒS$b����G�!��*flJ��fL"?	��[@�<u�!��X�
o��7-�\��@s5�ݺ�!�D�PCh*���(�v9�a�à_p!�1yQj��1�-0�TMr�"&_!�DT�Jh ��@{�F)
�N�8U$!�d�]�>�*�g�.:+����X!�D��~ɢ��Ņ#1rq��`�>P!򄞽(��t�߬#����x�!�d�C�D�oVRAq{T��$�!�@J!���E8<>�Ѵ ěd�!��,*�]�4�'LV��p���)W!���) "��6G��&RusF�F�j�!�H2����)I�P��y�-�=L�!�D���y�u�ӟ����_�s�!�$�"<q��	��=kn�
�#C�h�!��1:�Ҭ}k�)!(ך$�!�d�)EڠP�J́wg��=�!�䎠K����1���SsƵ�FR%�!�D�R|�p��%�Wfa���<!�D�+@�B���_�
Q�����!�d��+JE�#�R��d�/�b�!�$Z�:�1Ţ��!{v�0�$�d !�D�?x0Q�'�:B͎)`BdʇA!���!���7�<��C��!��Hl�e�`Ҩe��-�q���!�Da����@��D�ো&?�!�d�b*���I�UlP�kGeQH!��Z�&l�Q��6y� 9�'Ì@b!�G6����G%�a�,SZI!��~�X��E,�Av���M�y=!���,(n�ոv�Z<'�t�P��k��OX�=��� �={ 
ظ�B�Aƫ��7�J�"Oz�Y���(&/�X��ٴ�k2"OF<�F �a$X�p�i��Y�b"O�@q�@=؊	��H�:G�����"O��!Ӫ^G���1c	�]uFxp"O� �
3k�h�rf˱X(1
"O�Á[P��A�T�k��2�"O)1&KF(�NI;6�[6XN@Iб"O"\���ޱ-,��tU2l�DQ��"O�=KS�\�U���%���̦��0"O���$ΌE�����V�M����"O�$��.*7��3gV�@��3�"O���M]%�V� �f�z/��3"Oxi�&n[�t؃�E72�έi2"Ot48��� �V��E�E�&��P�w"O\Tkr8��Hǩ^�Qw���"O�X��i�e�v���E�kaȝ1e"O }8��/@D���[�fй3"O4���B��SCR1�l`"OB�Bq!��{{�)`G�f�����"Oj��\��B��>��E��H��l��'�ў�>9�v`�/�x9K2U�� �m/D��J3mT�>��h"`��5�P�h3D�h��L�M��@��gt�(0�%D���G@�<�XyBc��&`:��"D�d�D�>J.T8�G�!v����4H6D��aU�ɧ	PtI�na�	�qg6D�<�elAR�ɔρ%Y9�ݳrN0D�h¶�ӿ~\�eʑ	^�F��$D��Ni���������'6��C�	�$D���%�̥c�E� #�C�ɉ)(
�kU%�'F�!{A��Pn�C�	�D�Υf���>	v U�X3�PC䉹?*b���ٵj$��刔5�C䉋{�4!7,��JA����y�C�*b<�\��Å+'7:@bAZ K��C�"<��	�j��*m����'��C䉭u�<�G��S�$�I���40x~C�ɏ�fqk�	I�Lv��W#[m(B�I���H �D���&G��TB��=V���q��I�~���#p.�4[�B�I�<ԘXD'ފ���$��8��C��-c�����	ɽ6��	0����4C�ɍ,N~%yV+U�ʼ�"���NB4C�I�
����U���&�J��FAу:+`C�I�4�a�cT�6�(X�'�=)�`C�I�|��D�@���9��;�fɷ�2C�%FI��醇�֍�Js.C�I�r��0�e��2;�����~)��D{J?��2�J�wK��BOڄix�i�v/4D�hB')����F�14����.D� �@�2;����H��mǈ���++D�|�S�^�[��ɓw��-@�X�`��'D� C3��6 ���#�+)�
��R&'D��񅒒5���Ǐ�t҈�%�1D�9I5�0�;�!L.e��4���0T��y�F�%v�r$$�($"#"O@\�a%W�<j��v#��:�	�Q"O��1�(�X���a��T�R��U�#"O�x3AfL�nR�q��B��Q�G"Ol�ؠ!��,��iCp%=%Ot���"O���V(R�@��<����k�|bc"O1bwn�+�q`$�0q��E:�"Oz�+F!թyY�T�g�Ie2h��"O� J\���ՀsuD����@e: ��"O8EA!aW?B���V@')�L�1"O4�&ûi����3����4��"OHA����V�F�L?^����"O���GmO�}��I�B#Ğ,x��2 "O�0S"���D��T`R��(��%��"O�l+�/��{SPYe�)-���d"O:[3-�.L�
�p��N�Z<��3W"O6�a��BHZRϔ�5H��G"OX3AL�,Gw��#ӍZ�d2j�&"OV * (P1�&4�i��Z~�|��"O���T?���z��4%����"Ov��1�\j~�Ï_m�H�u"O�T�!Ί�]�0}(P�v|\��b"OlLj��ؓM�DȂ�K9=x-�"O��XǋZ?$�B�`H/q*Zp{�"O��GШ�Ѫ�Nu
�j�"O�
a�),�n�ѣ�0h���I�"O��/�
1"���F<��0�+!���!ۜœ@ϛ�n$�Xу�'-@!��7��]��d\l(��19!�ė�e"L�`��+�<��)!�Y	F�|��Po�m�`P �(D�w !��?WW�ա�d�G芩��(�_�!�Z<Q5ū�X��^0�T�ѥa�!�Ě0��=��Kլ%ְPk%i���Py�D[�H7`ŐH�a"�ٳC ��y���
^���s���40tzQPC T?�y��'����ո9������y���	���
ڷ�(�R�1�yR�N!Vo�Ӈb��qSV��r\��y�&�\t4���W g)�*/���yҌB}X����R�H"��{���?�y�%�(g�,��I�@�$u[�d4�y���}�7�7?ƄI��[>�yR��)s掄z�J�;�V9Â�ߍ�y��H9�Xck��N�c"�&�y� R�}/� ���(��!��k&�y��""�R�[��bh>mJ6�%�y�M7,S�H�#US ����1�!��ФZ�XT:v!¶6�F�i��H�ko!��%(�8��щԏw��u3��;mP!�D�.Tj@���b�@0$Y4È.!�$�Xb6(Z��HL��bB�PQ!�$H�[n"�uIA� ������8h!�䊃c~�e��F�#�:��ӊ>0!��y���!�c�{� ��EG�!�B9�%G��0{�9ׁБ:�!�䃡Y�\�#�/"la�E ��!�D�.)���z���}v���6%�!��T4x��B��r:E�I��!�d�W�&I!d�=v�P�JÏ���!�d�z�z���(D�X�|y���2-�!�䆽}z�T`����c���E�N0Ag!�đ=[E����(L�� ��B3J!�dZ�B-(�� �0�g���7J!��>@Q��`�A�$��"��
F�!��Y�6QJ�G�;ȃ���$-!�$��
�( �H��;Y���w���!�D�$n֒ ����')>����h�2}�!��j��)y���C�fm�(�:T�!��T�Qe��Gj��{�f�)�!�=TՌ|@vE#Z	�=���R��!�
�!)X�똁{Rݪ��/-�!�� �`�F�W���/V�Z����"O8�!��t��1s��ׯ���e"O��ұ؁Xr��,<Ǿ���"O�E��$�L"��Q�ڶ\Ÿ�"O��Ҕ�ݍ�:D�B��?A
�E��"O2�ʥ���J��XrW �3��h�"O�	���~Q�WOҹ]��,A�"O�p�Pk6V2�D�6� �3ऩ�"O��Qr�ק �1!g�'�4�g"O��It�S�( c�G�H�iG"O��8T��b���Y5�V>,>�Z�"O�H��Ŏ?3�\��ւ&/m�#"O԰�ĭ 1�֕���|�,�"O��Z�J�1�&T�1�]�Q�L��B"O8DZ1#�->�8�S��+����V"O����	B	��X h�54t�d��"O�p�scúe7t���͞e���"O� �#
T�@���pt���3\LU �"O��БȌ�^#�a�g�/�^�E"O�j�@��a�@����VǞ�""O|ݢ�`�i����@��Zs"O8-�aBGN��y�q,_�F�"O txA�t"��s�_3d(82'"O����GɫJP�TK�?��0��"ODQrWÝ�gE�AE�Έ3��19�"OF��`�Y�nL�JqA�#2TZ��d"O��B!Y�=.�0[��8-c��pV"O�M��9G�P�ӴA��\&��a"O�͓��S6e�ti7�.h����"OR$(�L	6 ��`@��5�=F"O8yB���Ё����2�k�"O��bc$ʹ,�@l����)�. �R"O��PѬ�+I�P�f�Tz����"O����HS�dT�1��L�0��U�5"O�S��	�h;ĥ����s��-�c"O6͘�I�?s60�3�#h�ƙa""OکC���_3
=�v�A�w��]��"Ojы'-�	~�p2�K�#;8�R�"On����L	-xâ@��/�8�"O�MPCF��S`�Q��$M�LV��"O��f��9�*�DT�>n�x s"O���L�ha�- �{����"O��ڕΓ�I��۔Ε�g�e�p"O��BL�	��8p�I!N����"O��Scd	0n�
���J=p�`"O��
���Tf��"�"Od,�0!�$d^�	��/H���`�f"O�8�#*��T�|��n��ii&�[""O���:j�P1c�*�:��"O}�1�J�"~05b�,��$*�W"O�%�+,&���eJ��Av��T"O���ǂ�;������
�.q�u)�"O`���c�	gy�8���0c���2"O�أIQ.g����IzK`�k "Ol��팷.Kp�	��\&x����p"O�թ�#�,wF��P�	x/����"O�-I�������C�y�`�_��y�ўYlX�!܂ql�x ���!�yB�O�8ü�°L�z��s���y�o�"�cV�B%p{b [�L��yr�I�5N	����n���C�y��J�NĢm9A&�'$�Ȗo�>�y�^%�:��P(�j��%���yb�cʮ��̔�\�"\X� �y
� 6X�djˮS��}(��A�KY��c�"O��Ƅ�>4���b�	�n�a� "O�9ZUk��hcd�`�9t�8�P�"Oh�H&I�0k&��B�ʔd�I"O�-
4�4^��(�@�Y���#�"O&�hC��4��=����a(��'"O.�I�g�� ��7hߩ9�D�"O����B�)f
z�(�F�!|,���"O*(r�o]�:��,:�� #I&,JS"O
!�r,S�>�����e@�fj}@�"O��)ӴS3���Sd�pbjd��"O8���	:��0��R7��1"O~(3��$yFH0c\�G5мC@"Oh��fzQ�,��z2��5"O9!4)enh��@!�z%<�
�"O��	�E�֐�!"�1��\�"O�<�* ��a8��8l� RB"O��(����^8F Z�-|�MA�"O��A����pk|�XbEļv�a	"Olm�3�L�1��l�s��2gt�ܸ�"ORհ�[�C�p�1���B�����"O؀��%i�I���	�r���"O^!c�k%[����g�S�ι��"O�(��	����%��I�le�\�U"OP�kEL�a��a��ͅlQ��C�"O$1�rGCR��Ԇ�1�:��"O�I��8&P�yj��žz�x�7�?D��rD�L	6H"ID��p��HC#>D���o�-%'�LA'������9D�ȣ��Q+��tѢ�ÜQ���7D�z�'ۊ����r녔g^����4D��QåK�hB�zC��-А ��4D�0��A!r6:��Ӌ�.sIXH1�0D����%߄d^,%��E/�
�HSH*D��(Ӫ�A��Jt6%O:e�'D�܈𪌙�n(�0 ̙.�����1D�P���0=m���i�!-��g�/D��j�jĚG�ٺdb��R��h�:D� �G*�su��*\�wD� �9D�pk���&�����TBx�;S-D����2%?�m��))lb�
-D�� 5	g���ՃCA#&x �i-D�(k%�%*�0���I����@)D�<s��'e��t8Ą�$,Qa��;D�,�&CG�e��P�/��x �y7D�8�S�C�E�D��$Q��1�R�6D����A
'��q�ȌjX4y!��3D� �w����� �#�L�o���f6D�P�r',Ev�Z��˨63�ճ�M3D��`��
�>>6�	3�
�|ћ�a-D�x[�{���YB�	x^9p�+D��Q�MI}׊�J��J�d����(D��
f`@���̱��U<*+p�&D�ĩ�67+
80�Ӛ	��
��'D�\k��%h��h��Q�f��<��2D� В�X�J�l��h�)u����+D��1���`�b�鑏8=2�)	$M/D��QBɯ3�l����F%�ah6�,��p<9�#�Q�4P$o�� �`�R�S���?�!A�3��y�U*�CO`!ȐCR�<�%!_�z:>�6
P7kV�C$�L̓�hO1��l{`�˱.�4ű��23�j�
�"OR��"��gEĈ`O�=V�8����t8�|��E�n6�l+WG ��Y�j.D�� �i�KG�-/l\�s��$��a��'��'���r@�ߪ���K@oi�)!�'��l��f�h�*ЄSrB����:�S��d�V��9A���M�@�A���.�y�ω(By�� �]�1~~��#��yR�:a��ASe��7/>�K��ֳ�y"h��tr��?@�TcR돳��;�O�L��R�:��@i�&Ġu5N}!�x^��yCe&�S���*D�ĠT%0(HQ*��[7��?I�'!\�����xR��#bA��E�\}!��7���"~��@	&U�m���l�1�NW��y�e�?�XD��#Bъez@
����<y
�3�d��D�B"N�C��K�QВ��<:�����P���*�G�/AX���ȓZ�N�{���&���z���w�ԹEz��'����peY�LS(���.��/3p�1���	p���*��9���k�JU���1�S�Op����G2��]��E�u��h��I}���I�7!c�4�#I �P΢���5f��d���	7�I?qؐZ�	R38Ő h�# D����e�>����T1#�>��*�O�}�'ٛ��s�h�� �ݭC}"��TN��y��dMF�CIM+���#�ގ�y�A�|��`cT��n���BVd���y�=|8� (Ҕa�<����N��y�i�l2e8���'EM�\؆$��y򃚵#�	 a6�����I'�ybKD���1�Ƭ��;:t���'1�yr'�u��%�S�L�+����Pŝ>��D>�O(`zPc�>�|�js�hc�h@'�'�	�n�<ӆ
�DZ�8�:k3�C�I3kP�C�B��f����#<���?U� Kת�"(���Z����k8D�|0���w�D��栞�~�L�2�<Q����K�aA��+����ˎ�!C�z��I��ؿ*����P�
a0C�I�l�2��2�M�/�|��f�#7i:C�I�!��]q�LY�GD4�QE��%��'�a}�eEl<�����P�쐪3�ƕv]��=�~"1K�>QȜ�%�  ��㍾-t�!F�n�<���<h�����j-b\��-�y�����(On�0f��4�FFf�`�f�)Em$�Ұ<4�>�Qj��|��$������v�U��E{���'��mg/J�w����`-��M:C�I� Z��p�	[#��DJ�&[���x���Ox�=�OD���A��ex}h��^s|(��s*��;�`��$ H�J��K�sl��O@���\w:(� ���9h���A���0���Fz�<�Za��ئ�����隋���x "O��pƭV`��Q�)կ3��	��S�'��>��- _���@F�9�p�ٱ
�
��B�	�Z�=����"7e�H )C�z��ד�?�TNS�-�x�R������UI����<�]9R�R0�JC�qsEE�<%�2 �4�q.ĴzP�e#�gVCX��Gyr���c����j��$��en��p>�N<!�lIr�j	�D�Ù���b#Mc�<A��_�<�8�{�&��LA�����\�<��M�3�&��#��~��� �Z�	|��J�<I���]�Ba��n,�O@�H�q��,�<��#Fѩ���ȓm,
�+ηKe�!˖��#�% )ړ�0|B��H�����i��U��Y��J�<�D��2�4��Px��9�Rl�<� ̔P�hC)����#�>[�ʸ��Oj)�Ɨ+�m��6ڐ��|[��_�<Ac�Q$`#�i7��' �
�k��@�<���	�FzHxr�L�!~[~u;�e�V�<iS$Ɩ\ ܡ�d��i{�,OR��hO1�(!@j^#*`0��(�1a�U�r"O�,�E��&ިT���U0PF���"Oڍ;Å�s�6��D,ȻT/���"O��7��0���kE67�"8Pc"O���	!
�̰�)D~����"O4Ȱ��U=T,�����O��l�"O����@s��T� �	> �#��IT>i8tDG�e����Oڲ;DHV��yR�\�d"�iB���4���Oʵ�y2��/UZM8��ϐ;ʤ�R�D���y2
�p�`<(����: �t���L�yB�d�8AH�=I�������yDB%�Ѡ���!AIh�����'��zr���X0�fF�fgj�;U����O��~�Ӏ3�j��������&ԕ:�!�Dӵl��@����=L�"93V���R�!�dC�W�N�z�D�����X�!�$K\��@Y��j��
e�Ǿ�!�� �D���j������E�9t!�b��]H��^7D'8|j��FU�!�$"g
�AJ�����i� j16�!��O*X�����Pa:�jդ�h�d"OV��u�I��J+#��XA�'lў�S:Ŝ0���R.�|R�*D��д�J7*ɤ �R��(�h��A-'D�\JQn) ����X6y�B$�d%D�d�q뇼��m��@�o$x� �$D��+�� �2&i�	 �� F� OH��ē7H���$�ҸV�����
	�w�BYZ��?Y��
R(sbgO�f�����5<��-Gxb�)���)x��P�ŪW�t��ΟW��D{�P�,V,q�1��*Tv�l����."�C�)Fxc��Q*a�&��R��ٶ�ՠ�yB"U*V��C�eZ!JwdI3Q����~�kI����0,�+W��'�Qtz(��r�5D�8Zt�W�%�����P8���gC D�<񵧃�L���G�M-;ȁ��O;D�(Q
йzu�Ђ�l�!\`�;s�9D�h
���:�ڡ�"IJ�č��9��D؞P�LM�X4�O-\����w���=E�d�i��sT���	�8LxlHW/����'����ӦO%Y�ّă�K��3�'�kE�[��&�>@θ��
�'.�@�.��Z$�/5$#
�'���Rb	ѓF��J� �.vgH�	�'O�sd́���4�Fe��2 C�'�����C�d򆀑{�I+�'޼�U$�3O��bȕkn4D��'�P��^�X�z�N��/���[�'1�Œ�b��M�B��TCH�-�p�'��h�Č�wJFQ9��U�:uB�'����.W#k��C�D[�r�c�'��؄�ʓo���rC�=�����'֤xz��ʨOp�5 2�DBx�i)�'���%!��T�l)���Ż7�^���'Y$��	Ȼt��D8�ɹF����'�� a��
�8XČE�E
� b�'rr���D�G� �$]����'1����Ib��|8�f��g��=�
��� ܝ;��:�*d��J�F'P�p"O���&����Lk�%��&��w"O8}��ˏc��s6�	�8�$�r"O��`��8��E� ]�V�)g"O6���O�ߎ�B ��9er廃"O����%L����`�::H�`A�"O�X�jT2�b��c��3_ ��'"O�P�s�J�KoH�m�8��R�"OA��LX2V�Fݰւ�/�ɱ"O���b*^�L�.�3�h�8�)�"O�5B�Kկ4��5�t  e�R�bF"Ot�j�����BRE��M�}��"O����
Q40�{�	�E�BxD"O��6$�'ƊJ��V�g� �a�"O.��%�V?<�p�d����Mj"O����%��0�\%�RfS����"O� �s앛Yg�����)�AC"O�x�A�G(��斢%T��`"OB��@���a�ꉠ���?���"O
�
��!AP`�fƍ� ���z�"O�4ɴA��
H���$ h�؜s"O
�xD�ڻv�Ne
W�aP���"O���4%Q�ФJ'��rF�MH�<A3ȁ
�6��C�.J ��g�I�<A��t�"I����;��Tz�@KC�<���H�z�q�V�F�[$��)�/P}�<q�����F�p��01����M�<�U��s���F��S�5��]Zf}3��N�h[�-C%!Z���`�M�Q�TqA��[	>B ��G,D�8ő�#rY גZ�>�HÆ&D�|��B;8��*Q��K�P��J)D�pS�K��9�dl*kP���0D���aF@��ը��Q�4���" 
1D����M�J���8��C@i�h"g�"D��"�]��z�f���jp�!D�̒ס��}� ��E�8];���A<D�˔*�HnX���mZ�p��8B��0D�$�0����&��Gخ^�9�$D��i�5�����*١?T���#&D�8�
�Y��5��W�*QnDAS�)D��R���'$}-��FH�$\���'D��)�@93�f
�C�-|&"a7D�P�ǉ�>[�B1k�
-e�
ЙƄ(D�4:�C,;WPt����u��k��&D�p��,��(���f�;]Z�ۤ(D����JC0%ӱ��;)_<Q ��#D��%�{���A��G�F^*\�`�;D��X�D�}H�[u�ŹM� �y��9D�X�D��\J���6-�/D��v� D��aO �4��S!Jj1�lh��<D����K�2;~�cP��b�� O;D�0(��5 ��K���F/�1���;D��˱!E�%�\bP�ު�bYB7�'D�p��BI�� y�	6�؊ OB�	FH��*ݻ{N�9�䄕���B�	!d� ��#G���zu��Q7��D�	�2�b��4����fR`t!��J�d�28:�#�0afX8�� 2!�L�8NУ�i�:�0yХ@vp!�䕮6\��t�	�4<&���<i!�Ċ�y��uz�	�@�nm��G�=l!�Ā�_"AhC�ʃXh����}*!��	+-��Aۇᆀ?SX�U��Y-!�$��lHaf	ΕB��x6+V�~�!�� ^d��nK}��@��c$|��a�"O���-ͻY*�#���?��m{�"O��8 D��N���Д��
Z"�R""OD (�&N1|¬P�D�Ǯ1KJh�"Oj�9�K^41�"�pR���R�3""O��;��W�(r��ZjN�w�B�`"OR��'����Rv��'�z��u"O0��1����2�Ԭ�"O"��`�\�(���Y��K���"Ol�C��Á'V���
�@�A�"O��ǉ@�_#2�+���7 �"O)"�CA �Q���;Z�0�"Obx)T%.p!^��S������"Oi)Ƈ5m���bh%��PS"O���C��5X�����W���k0"O�	��ע��¤�1_�=+�"O$�y�
2*M. (Vb�'w�<1��"O�a�7CxW��5�J�����"O�$	�����3J�r�<Q�"O��$ D"G"�\ȅ��vM�R�"O(��(Ӏ����Fb�f=����"O-�Fl�E���hR�.Iv Bf"O4�B`�,بM"B�DQo:�*t"O���ӫ��`x���g�&*���)T"Ov9J�P�/l&����ţW�T|��"O��i����1�@�23�Ic��h5"O�I�Eҕ
'L\x�%�<f��J"O�T�iF�1(L鳃R�u��{�"O���`�y)���⃷#��@S�"O�y8խ�S�� 8�!.}��`i0"O�҃�-�,Z���)��d�x��;S�1�=�~J�d��)�r����ыE�8s!COj�<1S*�!��
��؄@M�8����"2� �'���i-C=ĘϘ'6,����0��ti5/�8��3��v�hT0�܍B���ˆ�5���:��
 j{��l 8Vv݄���(逡�a��g�<IS�@M$���>��n�*c�5Q�j�5
�LJ��V�j%K�b�~����LJAX�"թW� ��=y���O��
W�%�eZEP������O,@P�S�+�L���T�N#r�Q<��z6�&J2�bYæ9z��[=A�⤇�ɪE�ؼ`�O��	]�Y�g��|'��jg�@5���۴x�J��b(z�K�j�,��G���<�B�"*����ݦ/�9�gCOS��Ы�ɔq髧��of$=2���70ft������a��Ңq�YqS�F.�K_>Z���61�'��ጇN��,��N_�^2�EF{	�"B�h�A�?;����cW�p�0���kL:��pO��5eN�)4]�	����(��u`* ��O�##f
�I�D��CE�?}�mP��'c���TJՙ?_L��a'Y`��<s�f��K���܋`�C:s�pI�h	�&1yC��ڼ�.\���o�()�OV���. %b޸���V�hc�@C��(�`���L�|������B��S�4� D�u��'� ��6���1Gݨs�B�S�O5�����I�4���"�[5䐍�����y�������J ���+/�4)�HIIN.ɱ�U6턵�'7.%�Ĕ?}(Wa�3O��%A�/�t(�RF!ړ�A�2� �n=# i�%���1PA�,J�a�5G �հ�#�-�[F�o'P{,O(�H������	�
j�:�鐀t��b6���9QB����Q�) 		"`_tʳe�	 ~�
�I��u�1�n5�VH�s���CmP�pЁ�DN2i� Ii���*9��|�lSuI�1X�kK.�$������]�&ii��ނ��L���ӛ}��D�M?u�ҥ]�5� =�'D���I��g�h]��(��s.�9�
��x������[��PEX(h6��6QT�=!��]aq�!b�P{u�i!�'��y��J�����J@)0��[bDr5¹!v����O^0E0y�P���Nƹ5�h�@���TlHx� � )�6�Ap�܈+ɸ)k �ŶqO�=�"ێ��O���qA_�[�Zq�3�����8��OX���*K��2y(�gYLo�� /�K���	��t��%)���x�& a�Q4l��yb��*������(�\��I�=㐠JpQ	<�:��-��=�n�[I?E�%%�)y�I�Lq0l���H�1 Bɫ�L�s{��D����p �&�/[0���bK�"u��8!��<j��5���-��5�V�8���I<|ʑzw�_ulҜ��#FP����T�R�4�{���5�M��ڃ?{�� H(p��Qm�K�L�L+��A�K�!�dT�Lt��8pM�+S]8�c*u��ɠV���!z��1=H3��4�ӮOI6�J�+�}	 EX�DҜC�ZC�I,�X1ؒ�Zr��(�m�o͊�'�v���GQ�k�zd�p���n≉g��	��ŗm���xMOK������d��ٻ�g\hd��J��>��4b`b�q�U��F�� O�.�Д���$���D@�=@R��#f�j��@���j��_2���ca�2)<�C����0!F &y\��4)��)r|���Y)W�Q&O�ҧ(�HQ�tbK�� �!P+V6J�$��F"O���@�\�(�6�P�&�^��0)�Y�䈬N �� Ӂ2��$ЉyV�QyTO�(&����"��P�}\(`�$� Ʃ8f�R�
|�2�˃�mF�u��	cG�scƙ�:`�=j҉ ����?9Cl�d�䘩׈�'�&�j�O��DB��sIs9��-(D�`jA��W8l�1#%^e+ ���h"?�C�
=�^H�A��N(�蹋�)�"y���r�[]��
� �30!�Lɼd��J�m�n�C����z^����,�'c~���I<�ѹ���|n'x଑c5m��uᬀ�g���yr� �F�~�����?�|�Q&����?yD*�8Yvz���7lO� r��Z��^`jGE�,Tl��q�'V�Ђ�E: �(n��C�.��4C�����6ND�&��B�h_��`��V'�����,&��������2ܪL���ӛk RD��͈�*s�Q�wK`B�	W�$�!^+DJ��Ŏ7ADtI5�Ix��H��D��'����D	C�Fi$� �76Ly��'yy�2 �<Q���#�ҵ=�X���+~�C�_�<�(���܁�*HJ�ݔ@
Y[�e�T�{�@Ѵ&Y��pu������D��X-����+,n��4D�����):?��v��0��q�N6#l��z�)�h�n��TL�"e�� f�A�Q�aY�"Op��P�J�2hp���@w0,
G.�
ݹ����O�#Ȉ�Ey�T��oB��j1"O}z��V	V9z2]�}��%z�"O�0�2��Zc.���$��P��\�v"O�wnB�@x�2ǉ�1;��"O���!mM
�䓢Ǐ����"O�+���u���
FF�%Q��*�"O��S�%�l`�I��G�0�d,�7"OP:7��E�LA�p��`�~l��"O&u�@%��i�0衤Ր�a�"Ov8��m�����c\�r��]�f"O��u�M�
	6�bg��s���Z�"O�582.�/s�ujvLH5u� [�"O(T�R��;�"q( ���ײ�y��W�RNxY򴏌�V���S��=�yBh�@{�8�7�Ż{�
9h��&�y�/&��ݩ�@́j�*�Y��	�y�/
6�b`�[�1yp(Qn��y�/���I�" �>��U��;�y��Dl���	�?d�@�	�DH+�y� .�:Xe�@�e�uH��޾�y�aАn�`�£lE3 ŐAL^�y҈��q�D}�	U���Y�K��yR�Nk(���Z&rp3�aɋ�y�[��(! <K�X�����y�΍�\�h+�l�� I�0/��y��^2>|����ͺ	r��@���y/��tl|��e�݈
�� ��2�yҮT�Va=J�AȑJ��)p  ��y�7[��}z#�
�%��:�y"��d[zX��K�x���Ÿ�yB�O-� p�W,r~�	ӑ���y��_�5[���FU�m�(̝�y
� \%�-�=p����a�?z%0�"O���@k=Dp��@��Z�j���"O^x�cNo-��fe��f��E"O�$�4�ݣC��xb�D[�x|",��"OX�H�J?aW�PS��X�c1"O�	b�MI$K�PQ	"e��tU(l{"O�9Q�` �h���MO�=�$"O
(*4�&\gH��NJ�Ղ�"O�E!�	#��it,Ё-X��R"O�uÀ*�9V�t��`�� a��	g"On!i�M�.ќ|�u%\.eT���0"O�u���2 6��'Wucʄ��"ON�샿vl�zTo�<WPtt��"O�rF
T��t�^,Pxx4`"O��r(�[�(aN��'Zt}�u"O�A$h�� h�,���9m�6�� "O���E՟#�<�0�}����P"O���wA��/(�x��ݑj�|PQ�"O���Űw]��iB�'N 0�"O��pm��:��Q,d���&"OR�ZC拿6uL i�`٘|�X�y0"O&��1�B�;����ca�8�����"Ob��'�G�R����1��*F"O��3&��(~5TԠū��|�%�v"O�\��B%7�s��H&a��W"O�gD]�2\x1��
�h����q"O4Jb��4�������.�t5�"Ob�BdʒP��R�c�8��""O��:��A�>o���U�S�R\���"O�Ti7�U/��J"���T pH��"O��Q�H
egZ*C	S�$�hY��"O&u��	�>�0��`�r	�(""O���0k��(�L�+!�T�X"O�2���.B����+�2^�Y�"O&]���Dds�K�J��@�"OH���R�pZ���Rߊ�#"O�I��@*F���z�iB����"O&EK�M�hW��;��H;$�{2"O�(h%JN2[�D�"U���5z�"Oi�qH�?7��+DG*6��1"Ov�{�ƚ�{�>p`�H��S�2�K�"O��k􈅡j��}+�	[)M�r�zU"O�L�Q���<x03�\�wӢA$"O,C�`�.�:Y��EW�fozx��"OP��"S**ȱ;���)Wh���"ON)�)����X�����	5�p�"Oh]J�D�.b1J@�O�5�+�y�<�5��)��D:,C�}R�!�5mw�<Qԯ��p��XU��A�D]�0eCF�<iE� �3i��7�H�Z�"j�B�<�G��R%n�z��YP޵:`�}�<a3MCq��ɀ�nS	U�$T���TQ�<��ʀ#��WO�p������GR�<��d�;yW
��-E�ܖs�`@N�<QD���]�<�y�F*:(��9%�FB�<Q�M7f��xʵ���9���Я�D�<�C長[�D8��(ם(nT<��	X�<rb$��)F,J`�Dي�/�s�<!�H�R�ݫ�"�3e(� ��]R�<��"�[=��'���P6��9 �p�<A��& ��jS�^^|a끅m�<ɷf��
��S��n#:�B�i�<�@�
��A�I%RK�Qׯn�<Ag�J�N��is6G�'����U�d�<� f�@5���K� s.ۛH< ��"OV *�h�'Sp���/Q�Oj���"O���!�!F�^YeCZ-����*OH�@2+V)#8%��'_�24R4�
�'a�̣���Z���X� ^�+êp�	�'�$�y"L��F8(�Q6(���A	�'��|�� ,I	1M�WzA��'�6p�5�W�&Gn�sf$A����'D6�g~�t9#/��w�Bٰ�'�^�2��3\�z�c#@G�Z1y�'
�<0���DYcϊf}�q*
�'6t�C �|o��R�X_d<`��'� �2hA'��`��l�=Q|�){	�'pF��j�w �P6�P�_�~!��'�T`�%
�\0��5��WA4���'��2��ÐI�:q�dǂÔ���'R���a����I$ċ�����',�|&�T}s�-C�{����'2��
��Lit��1m��lI�'�q{S&]�a����X8>��'_�eǟ�|����#�	i
�8R�'uX�Z�'Y�Y����k��di�'`�\;FeU�{J��ف �`lЂ	�'`2!R�a� k(	�p#Չ@�L�S	�'��Cʋ�5EV��cfEC��:�'U��&�&:�!�5�?�e�'$�[�h�-?����EV�ܡ�'��(�C�<:t6�c�M�v�S�'n��3U�6I@:Q���<90���'i`��.�c��12	|*�݊
�'��%�mM�\�8�!�� /�P�
�'�����o�;�r��c�V���Z
�'�8�bf#��p��"R
y�\���'
N��OۼN0�Qf�i�!��'�x-�F�\�t�
� ��q5^���'� ��Q��� ��@��m(�аr�'�
,ҡ��*6��aD�\�b���'WL�
���0��	���!C���M��^�{Ò\���՞bXC�ɀj�p�1�E?D<8cU �6��B�I�e�� DFʴx� �&e�&
f�,H,�2��'f�>�I�_?4)a��\�3�8���f�>p;�B�	)!$�Z��ݿ|�!�'��!"?�6�\���۷2�O~��%��94h����?3ۤ�W*[0T��cÖ�d+��d��,��<)��� ��ya��ŔBe� �k�M�<g �_�X�ɤfu��ZȀlZ7�����鍥*�& %<� ta�O�E`N?���<�4�D�������#\O(��W"_-8�6Y� ���:�D��B��@H��{T�3<߼5:'�U�->dY,O�t۶<�3}��֝gT��A�O�4�T P��8�'(0gM�x���b��B��f����q����las([�F����鈺]��@��0>�B#B�8��A��e�n�	PG�)/8:t��lQ ��;�@˧140b��.3�H�'h�I�6 �r��&�r���1
�'��x��j�6T�Ƥ��*� l��m�f��&}��P#�9�"0�6�\n��|�/Ot��`@;�aK޺\$���L�c�xT��Fr��8+�+~�qF�F�{�t���:N��h@�	D,=�tH�I
�}���Y�`��a%/�q��Q�1&�r��� �Nb�	�=Q� %4����O�2j��t�IX�f��T��!� 9b)�l��x�!��I�����'A^�	�mœ^�Bxz��.1$�͒r��X ѕ�D&4�0�CBX���W+�д��댉��$��J�%����T��-�P&��L)!�dB�š�)f��$Ql�"�V� !�2D�L��`.����4��7�T<��+�|�c��8��@���D�|���w�|���ط
��x%��ۣK�"qN��f�8V͌d�PNQ"!p�kBTX���=�#
,�Y.҈�%�� ]�%p�B7LҖ�E}M�[�FQ���B̧p�RA�c���W��s����t��S�? .�Y�-�458������Xv�O���a�Q�s�|�N��}���ѭ?�n<�5-Y�͚Ԋ�j�<y�]S��i�CCX�	N�LS%�f�Ć�{�X�&��0<)D���J��+�4���qň\8�,��#��q���
�;�&��)_!8�"]:%���>�3�\�6����'1x=p�䐃s9���ɱ0@ �Op@U�ǒac>��VI-׃@kܧ'�|
�K]Kl�B�\lɄȓ	�tHT�֒?Z<�y���E�����O�����3m���%�IM��ē`6�P����H܈Ȑ+�,��I�b0�PHͦ�.�i#�"e�,��f�[$���?�v�ϼ7�����H(Bl�A�'��x��I6{(�$>��0մtv���J{3*���:D�x��#ӰoS|�p�dݟP6�VC�<��#őspZ�@ ;}��	�x�9q C�p�qR �y�!��(�6a{"GN9*̒��v+*��O�1փ�"�X��qO����-~�pZ3�V49 �YQ1�'��4�̸D����m��@0v@�8!ؤT�h؟dj��>ieʕ ���@�X$���;�r���'�T�� �s�,[#���Ԡ+ff%��"�	���\4�y���B���b�O���6舀���<o4� LP�R��r�1ڧ
�I[¥���X��]-
���ȓM�dI�O�	e'�P�b�/S���Č��(�@f�'-��"5��^�g�	�I"��;aO��F��AE��
jB�I;#c�}˲��3��m�0Ba� ��ܶ/�^#�ا��=��#��F��
1���2�i�}���8#/-5���릳i��|��(	�0�`�ߞSe�	�	�'��Ig1=��A�g�CB�`�Bȃ� ��#�N~�O�|Y	 �X�|�Fl�a?�q��',tU1�/�9c|���K_4X&R������*$�c�'}�<#fڇ��[d%"K����'0D���MF���ܡڶ:�������O`�`�OO9�}�ۓ>��.[�ިzvi�0����ɪf�z��w��?���C8 ���
�GB:f���cU�y�Ƣs�y���!S#ԠI�%���O��S����G�}���,S�N0��N(r({��N�<�#EN�l���8��U�7B�=S�Lqс�v�S��?rAٍ
���x�R##��q�Ҡ�j�<)�M�p0q铀V�g��0�%)Gm�<���+a�~����~0����@d�<Q�N�-I>���o�0~V��RA]�<�qB�
U�Z�E�RT��D	Q��T�<���ݞf<��ZǏ�s����D�<I���X���A����2�B�<��b֔x{�eH�
�*=�(i��q�<�u_q�4mr!.�'_�y��
m�<a��_�:��T�� *#LcS�b�<qf, �;\��C��`��fK�V�<)� �4~�T�c��T�)�Ҙ`)�D�<�$�כ<34ش�S	z6��"�X|�<qV�ͅ��U� p�E`]s�<AT��&w�R���etNN���e�{�<)�4oP�ݩ���uL�[DDr�<Q�GN�\��в�é'�VX�2�Jl�<���<Z�t��V�32��n�<ab=2�>�0���+I�6|a���k�<ɕD��Z�����h�-�VA�a�<Yj�m	"�[��̞,g(|1�T�<yAh̙6���`�9�bY�rL�W�<��b�1"kr!�?;Ӷ��Q�<��c��4�w@��(�z��φU�<��M>q-���� ؍�P ���S�<9����YСC�O/3�E(1��w�<it�E�*�Nɪ��A�̉��@�p�<��e�,��L���<0z�z�&o�<� "�!ST<@QϜ!op�͈U"OL, ̊�(db�!0MU#X҈{�"O��*G�B��P�mN	 .��"O}���B� ����m�(u"O�P�� �bX !Q�B>�p��"O�4xQ듶B�y�8$U�"O�UK@萤RP��¡�J(n&���"O&�yd�4\rYqUZ�,U�ɋ�"O������q�R`Ք@؅)�"Od�[q�Gc��a�J߬UH�8�"Ot��\l���r6��K�^�#�"O����Z�'@>0q��U�wv��"O�l�7�A�N��P�3eg$`*b"O�$��mǾ`�
3փE>V��"Ob!R�m�=,��\1��ߋs�88�U"O�	���I��Db����x���5"Ovd*��R�w;����R�<�6x�C"O�ݳ ��&�n�cH�ki��Xc"OM����8$59�fɱDA��@�"Of4` �_�^�Ҩ���>l7��R�"Od�T.X|�X�صy"�Ls�"O`h��i�G�N��#nك: ��N�<��dÑ��m�L�:
�1 e�B�<	n�h��= #�W� �DQ�lK�<y�h��%/6����qj��@�G�<��q �)G'	�3�LMA�<�bЬBv�$�#Ļ)Y����l�A�<�g!V�o1��[%�
�KiB�R���A�<����go��0"Iޮ>����Jy�<1)N=#�69P��96f�҄�s�<	G�̣0s�<�Q���j�f]��s�<���
\�RAR`E�9)��q���e�<i�#ήDkH�!�K-u���c#�c�<�cbܯ=M�Y���0U4,���-D���vaW�݆�N�9�n��z��B�	i+��R� �?.�P�`�1�L�FBJ�r l���&	������n�f��e��{Y��M	jW!�d]4nP	:�쁖af(0Q�&�7tO!�E�b���Xt(N�H��P*���qc!�۰Z�������Ƞ1@�NY98W!�G�P!E�F�t��B�+��P!�䘻n�t�q�M�Ts���'�+J��z�՝��a�p����!��A��_�SԪ���H���iUs�>��'^�Gbl4V�V��kn��������O�XIe���hC�H[<<�5C���V�$�o��$h��)��	b�S�,���R�#Lo������&GK�5[�'�qZ���%�>)z2�Ory�+�.�  ��I��Y�X;��>�J����\�������<E��Ǝ�-w��8fE�B:�h �A Un��2G��aR�- ��<E���X�5�͑i�6K>܉�SFLm��zS ����0�a��.҈y x����ŐԂ�� A�*��'� ?�EI�4�q������0�\0O����,c�^���O��m��&n)>|�.�M�O����B��a�r-�mY�	��A	�+�� � .[�Uc�i������M�O]��Ww�My��A,cC*5!R��
T�0�Z5g{Ӕ-�%�H�$@�r����H���J�,���S͔
�Z����]����ri�	3�D�$����S�RNh٨�@��/�0����S:%<д��L�ɦvNp��g�)�$N�9� 򁉀�7�P9Pw(����5�X)p7�����	 ���������5_����婌SJ��Ѓ����/F.Ma��rE�`xݥ���OwV�3c���%�Ԩ�Be�uY�F�S~r)Q�-�����|��i�z�j�W�*X?\$��b9z7�$�<r�t���C%|O� ��Q�8��4b�;8E�\`c"OR!e��������3v:�Q��"O���w   ��   �	  �  �  �  �'  1  �;  �F  R  C]  ,h  %t  `  ��  u�  C�  ��  Q�  b�  9�  }�  ��  �  C�  ��  ��  +�  l�  ��  b�  � -	 t � ; �" ) H/ �5 �; iB �H *O �U g\ �b m %u g{ �� \� � )� m� ��  x�y�C˸��%�RhO5d��p��'l�I�By��@0�'�F��L��|�t���pd��46��-zw�G$�`�	�A��{g�cY�.rA��͇A�BY�G����u�蕦f`�T��V3�$��06��	��d�<x�-c��3d�v=Y�	9mC�����UF}s��^t��֝CB���M�FH�z�e����В.Xe\�����.2H¥В&|ت�)Z��7��	�:���Ot���O.���4r���Z�*�X�#d�څ'P8��O���O
˓����O���O����\�Q�x�tc�#2&���O
��5�$��o2�d��6����?R%�Ȇo ��;�'Y�b�F����d�<�Ф�dAvZ�`�*r��1�Kǟ|���X:�8P�@&ϣ\@u�O9)"0�_#{�(�h�e���������~?�A�!�O$���O��D�Oʓ�?���D��#�$�J��߂��1x�k���?���i)�7m����K�Od�nZ<�?�ߴC��	/+��%+���/����EI�����$4�j8Z�"X�E�ʔ���LR�R`�'������8ݞ�hr�� &M�f��OZ�=E�T��1u��Vh;l�H���jy�	c���r5��.!�r����Թ\�Vi��'�Ij̧öp���ƕ��4b���<N�$��f����!�� \2�@Y0f�C'=2i���<���K�}�8pn��2�@�	,hP�1�.�3H�\hV��?=t��	^y��'��<�J(J�'1O~QhW�Z;1(
��0�T�*�V`��'�IDyB��;:����FU`Id@^��0<��������a~
�8b���F �@O�I��V$�?).O�=�}j�E�:D7�EЧ��9E@v��\��4���]+t�6�}صi�(�[�0��IK��HD��G���O��aB �^�
BĔ�n�nU�Q�'T2�'l�A �Ѧb� d��bJx��4	�'k�TH+C8�Q1��G��| �'}T��7I��B6��Q�*@��z�'jb�p�ًa*؝����%V�ș��$t�O�@L ���/�:�Y��	�N����~�&�Gx�O^��'��l=�8z���q��U���иs��B�ɶ:*�PQ��P�1zܘK"��HP�B䉽�J�����6��(�0�\��xB�I4X0�`�ġL���w�31B��/Vz��T�o���U�<��˓-Z���|�P��+N���K�&	*"�܁����#=z���O��Oq�� S������HI�+L%~9��"OtA C)	�f*T�pe� *ꐈ�"O��3d!����`GR8E��zV"O��fZ�4g^� d�S���y�"O���GnǢ7{lb�*��%��`�Ғ|�6���6q�T��4�?y��PDpL0�@�e f�Bb��:�h-9����O���d>)q��UѦ�<q�eZ4z�@�X�O�8�����OF��:$�c��}��`�s�,D�����'� ����c����Ԧqxڴ�?����dٞ��"�� r!�6��9���OR⟢|���E�|�8�@gL��R@�U�	{��Lh�L�\�Iv���fO�|��i�	Ay2 ��RS�т��9O��D!?��$R��M�@@�)c�����OL�xG�/3�qO>5�g�i��`r�N�(q�d�P�8?Ѷ-Q8gK�"|�U�����A��6�t�k�o�j~bÖ%�?Q���'��O��eW.�)�ޕ�H)_$�@J>���0=饭����c�j�Mڝ5��L�'���}�7���V,���M"?��H����Mcvm��?���_n%{�'�"���?y/Od`S�k٦6N��y���9�B$ya�$�I�!ۤ���W�/z���߱G�q��#�;1O�����'9�y�`�Uk"Й���lY�\������QR[r��'Y�	�����K:u�0�������U0�J��Җ%R֡��$+���'�h#=ͧ�?�+O�0F�ΊE4PIF�	>[r����GO��$�O��$�O\�O�'�EH���159���)��eW���cIW<q@�(1��(�ɖ�Jqz� ��ہ������2��8���C�4����lO���ܛ�.Oٟ B�bϐ�{�J�4H�X٥�7Yѐ��il�dq�DC#S�����5Wt
&�Tiߴ��wuN���^�4�����<C����^�q@<����wy��']�'ζ�A�-٤m9��1�'�� �I��@#b���h�ԘlGFU�q�'Tʭj�*�.�"�:�l^Jhlsw������\��h	{�B)e.�Ebs�`8��$�O��l���"΢!.��� ;8 �G�ny2�'4�OQ>Ep�퍽E�:Ex�k6=�8s�5�O��l�>r5J�S�Y�����͖]ㄘ�	{y)R"t7˽`F��D�|J�'�T�V��y�&�u��=��lF<�?��;���D	���T��?�/���'>2��xUNM"h�0Q�C<,���-1?)o�v�ބ�NW�. &p��a�O�b(YO~c�@3>���[��1H	JE�V~���/�?I�a���'�>`�θ�,��Ǡֳ1h���&-�$�O����� k@���a��&�z�џP�4�?L>�i��Ɲ�a��Oj�U��Z���-lk��'J��s�O,��'n�U�����'h��q��� W�hp��l�j̓v���D��8"l �b[D���+[�1O:T`��,D���=r��T ����	r~�쟩�?i����?!�Oe�d�քB�R	��K�	G01��t�'~v�B�fQa�	7*��.O�Ez�O�╟����W�M{0Yb��nw��{�L�<9��7�?����S�''7�u��̯8Y
��/R�s,�Ćȓ1�Ȕ��.�cW��!"�.�e�ȓhR� cEP�I�=�Q�D�W�L��f��u��OF�g�RgeK*p��ȓ<-� saY�=�]1��M�I�Ό$��ʍ�D���DO�\��=*���`@^4qL�|R�',��f�� ������B��@w̨�����*�c�A'o�s�r؇ȓV�\�'�7x �%��-�E��QR0��G/�<�V�8�
Hn����	��?� ��s�dС y�\Y�o`�'�}��)��f� ;�m�:�\%���[�A�����O���dWlS\d�W��"	�:�#�lm!�l�2��ҡ�@�FY���E��$܂Cr����/ gl�E蓬֢�yR�'`���C�'F2�BYj����O~<E�D�V|�.%�mZ�
vEbC	W�?9��M����'u�@@�H�Cm%B��®,���L-D�0q��1ȥq�
���`�ж#/D�,g+ܦ0��`��v���a'D��p2d�):I�1�L? �Jh�7�$D��H�J^�E�6 �a�:��c�<!w�)�'orNY��AD�!�X�/�1ne�'f�y���'��|��a�g�	0��� C��kSn��y2�˄m)�9`����j��Q �yr ��E�t=Z�c��JH²h�3�y�j�VÚ�S�ĐDIquʞ�y��	3�r�b4�P|Z�!%�K;�����pi6J�� +^�:\�e��� MV������|�'���#�t��!�!`���_�5��`�ȓ�؀#ӮT�d���X w�$\��3Z���A���SG���UO�m���ȓr/�Tz�⒋^JR�ѦX��I�?Isպ?� ����?c( ��SnV]�'�,Ṋ�Iݹ jh;��F+w��q�u)�P�(���OH���HlEj���,��4jtgX�}�!�D�j�7(Ў�&�p���Te!�$˃n�5 "#��Qz�|�JC!��ٳb�
d�D���[b���+�>;џ�я�I��	.�5CPd^Rt�F�C�b.�P�O�I�O|��6?��jy�!mW�����X�I� B�ɗ�<5Z`�K�<�鰡D�M�*C�I�eb)Y�9.� �RR�&i��B䉞~a��$��D���ABgR�WO�B�	($��y�bN
� ���,Rx�rʓV���|�r��(R�4��.��ak��shFMy��k�B�'%ɧ�O�E*�d�4�>�k�9;D��	��� �TI7�I�M+H���D�5.84E��"O��c2�RC!�˼j I"O�|9V��
��=�׃�~
�X�"O�a��L�bW�T���)G�mP�I��O����OD<�@�"�ұ�e�0;��t���'~�'����>���i�������De�<��-ߐa��xS���6��x��F�b�<�#º@ǲhfNG2@D.�K�d�_�<�!��	_�Q��I�T�4$#���f���Q�Z@��:���*rN�bƠ�0dy��E{2hɯ���vm��`C^��*e�#8�4����O���+�O�l�"�(ItI���4~U��"Oҁ ���(ؤ陻{r�J�"O^ �ÅE��m�0��S�   r"OʭJ�++6L �4G��H�������h�(��T�Ͽ0{�(+Ѡ%���)��'����4�����O,�1������.%��IT�ф+)h�����`��
S����S |F$�ȓΊ�`%�ݼl�(��we�?hn���ȓ')R� �X����n�>8 y��Hsн�Ш��H�\T�c��w��Ֆ'9�"=E�t�štGt�`���e(�DK ň���d
4!̖�$�OΓOq�n��`dB9��=�g\�n�8s�"O��JnD:�j���
�Z� �p�"O��0%F��s��XF��s�Ꙛ�"O��$#	��8I���	P� }��"O���M�O)�����'Űtz �|�)������U�XuI��.f�Yb�3W�l`��A������O^Y���6��`k��$�Vs"O6�K'��U&BT)�C
;�~4ʗ"O֕ã��$��qQ��Ҭ���hS"O��Ў�8nTѤW�-tq���'4��ĕTS�P�2�T����{ ��H�ўH���*�')/03eO)�\�ɐ~ �lj��?
�&���SgG���ԩ�ͻ�U��on�=q�#�j��@q��68_\����.	cWʄ~+2	�Q�B�Z�(̈́ȓ8�V�7��3�t٘�e��mfB�DB�#�':�� �"�]0���/���ɍS�&"<�'�?����DC	a�=赁�
u=6$��(��!�Dɥ6��XD����HƁy�!�$��6�%{�j��KHXSTĂR�!�DG	�`cNeF8j�,���!�K�A��`��¡A
�q@K�ko�Ɍ�HOQ>��
��11L��/A
u8��2l�<�֬��?�����Sܧ�&���I�8�l�+���v�6܄�~i�ma��#�xɫ�$��v��لȓ_�0�G�ˮ�"�kF)�=�Ni�ȓe�h���%�M ��B��
K$ԇ�H��	!���ˬ�2���1��e'�j��$'53�䓋VF��$��bu�(�Ҏ��?b�|��'_��.x��&!��[Ɯ���-_�E#bp��v$��P�n�.N��F�,��ȓ0ќ��q�٤#�K�a��AN����������	�U��T���RY��h��I��?I��PiJ�����X9~ƭ�r��s�'1��ˋ�		aӪ4�w�Z�fN�l9�mό�����O����աN5*���)՟GAD5�Ј�~�!�	0]�0E%��
e5�!��$�o!����2|�'�ʏ8Sr�B��D1s8!��V�1]���B�>Jl)U��)џ����L�wh��ӕ��X]�S͟lr�G��O�	�Oz�8?Yխ)�t��S�ђ}�Z�f�N�<�6�gTީ��7z%"���K�<� ,�E�׊�(25�`o^m�P"O�� �	Ĳ2Y�Ũc%�[W�H�P"O�x+A�)��Pт[H�C�X�(0���S(\J� $D'�.���D:aK˓rc�����?�L>�}��C�q�@E��cK		J��!�� b�<��̡z�4y	�"��v�)v��^�<���͋e�b����T=89�taY�<Q�IA+7*��c�6w��Ty��[�<	��ُdc����G�6M��l�~�I���OX����O���$@$EHN�-^�N���'r�'O���>Q��IN�m����v��q��~�<���Z7}�$F�sq&� ���<i�D��W PIWb��hn�Ҕ�e�<9�eG�R1 -SE(
�Q��9�eO�g������`,@(�}ihU{`�,(h(F{R�ܧ�"�a%����! ��h�p��AA�O��D?�O�s��@.B��Y;�n��E���(�"O��Q&���yQo�_�@�a"O�h�7N\_�$!w�Ĉavn���"OPAE�QY����5��k��ɶ�h�Bu	�Cq���ț[]L@Ӌ\#�?	VXN����'�����Xs�1L��p��%+I��� �$D�,q�cD��=�B���T��4D�h@�J�,����n\=�T�z�m1D�����E8AFF}YEJ�4`�t�J1D��R��a��D2WےU>|`)�<���)�';@@��2C��M�*e8�m�6'&^��'ȘP��'��|����Y�+����BE�r�D�2`T��y�����n%�vπ# Z�4�̚�y�Ǝ�[C�h!mu�q�G���y�)�0N-B�[s�[5�V��
�y�	
P 8�#Ϩ<��}��`G.��C4����G̨�+FK7sj�C�E��0Z�U��'�Od�O��$!�3}���Ah�H��Ҹ!�������y�疷N`��]E
�h���4u�B�}1�A��k�^��0BM$9E�C䉟N�z �ЀØ$(�Cv��v���V���p0,G�U�8�b	�����A�h�x"~��JX;4���'�	n.mZ��Ԇ�?A���0?��P"K�UbrE�e�8�j��I@�<	`�"p!�q���~9Ь���|�<���|TqB�#:{)��2E��^�<��
�E021t�E�r��1�ӣ�o�'��}z�(��t-\� 4lF9�|����ƟĲ -*��|����?y�O0"@ �� �"�5o@l�:�"O�ȷ��UŐ�y� �;rX{�"O�䳁�D�;� �E`´.˂�8"OHţ�'.� ˔��%_��Q�"O����GU%K�`����V9X2hL #V� y���S�2*�)�ᑕD�6JEaɩJy��8�������?9J>�}�.X
GG�ٶI#T"�a�c^V�<A����6�X�Cv�M#�D����
R�<aH�A���A���&�P�<��b�1'L���G�& �ӄ��J�< �ݷ
 ni4���2�=��]�I��O�	���OV��� -�r�
�JG�zQA��'��'����>�C�~E��:D-G�q�T�r�[�<Y��K/4%�eA� �~V�� �#�r�<�F�ő��ʴ ي�L���k�<�����Z�pS��D+���a�L�d���Y��n���+۱j���N�<.�iF{R��䈟�,�d��>����D@<�|�*u(�O<�$(�OT�s���#r枽˱.ԡ6;�Z"O�9�F�Ѥ&�6|:�m�_	���"O� �Iz�޿�xyB�A�"O���A�J L�,	S�I�Z�����Ɋ�h��E*�-�f���4Fi�.�A#�'!�ݒ��4�l�d�O�=i������%k�2���\s���ȓwn��3�)�h7��#�,��*���JV�J5D,"$XP��N�~1��v�8� �n�$���r-�Rע	��%����s�*��qĜ����'T�#=E�$�����!�	8P�� ���+��˓X��9��?�O>�}���̨`�p�����t5��37�t�<�cH8X-`\e�_�*=$�#a�o�<!"�$i��U�k0e]��bNQh�<�rhU�
n��cBHA�g�F��oFh�<�5���z\�R�o�RE�����h����O:����O֤q�EJ`�1U��:?4����'N�'>���>�AFW>!���@��Y�CZ��H�"�_�<	�M�\R0<7���v.� ��u�<�1��)rj�c.�?�,��1��J�<ASKԑE�<���:6�H'b�O����]��)�L������bչT0��D{2���ڈ���$���)*v��b��'�Խ�¬�OZ�d%�O���+��]����Q�&��"O�HRMR O8�$å�0nŘ�b"O�]8Cl�ԕ�B��33����g"O�Y�V��`Pc�j��P������h�0Ek���+#~�Ac�Id��Q�'�@���4�D���O���M�R(���\8@�S*(��I.  Wǖ�TB\˄'_����!
t!�s�p��ȌV��`�ȓN~(9҅G<6/vЫҏ��x�"L���U��%&`eZ���͝}/>Q�'g~"=E�tAMk �7�]^��X���v��>II��q�ҡ�MS����?!��~�*����х0��xˑN�3o~t�/O����O|�d-;Mnwc�+"��8���1���S6�T%`�(�`@�fn
1�#>Qԩ_�2@T��@K�;�$�	�Ī?���.�8ɂ(A�Y�R� �Ѷ$8�w������h�|�W��#�j\��C��"��R)�ky�'�a|MNvR"�#��D�M�a9�����>�Y�ȱ���	5�`�G"E.�x��5��<iWL�P�&�Yv����O��J-rz���@'�M����}�"�M2 d�X0��Ӽ~۔��6n��=b�I�'�d;��
D<: (��Y
!��Γk��9'�Ǚa���	�qYШD�Dd݌��A��� �n��1��y򩱟\��h~J~��OpM:��$-�;q��-{&Z4��"O�Y�p�37������R�khh[��5�ȟ�F��RP��#n�/��XU�"n�Z���O ��P�Ȧ�����	dy��'��H������řD'���CX�\�(r��O�؇$��UH��'�?#<��D�9	�~ܐ`�#��@ ��4	$&$��� Et�P�l�7@.���Ory�cZ li���}/�������8�N�O:���Or�lΧSuPP�f�q�4�H�ソۂń�v����KIe*�Z����	��i��5�HO��O��4�"�X�D��X*��G(�8N�Hyp�K�7N�6$�� ���'���ӟ �I�|b��U$n��8!�� b�T��"/�73ޘ����� ",�	��۱�ay"F�X-��@�NKU�
�2`�7h0e��*��@q�l͝e���$�U;����42|�B�+FI�,�&g��S42�'$�O��}�"H�/r�X�ـ�������yR)ȫZ&`@%F����3R�����ꦱ��E�iS>u���I*��]"RHfQI��A�D�(�|��'���'�P���'�X�Š�O�ԨB�'̢��L�Qsh�X�HW*H�*�
�'���P�I��|��:��M��'��"��ζ,h��-����$:��>�[��B���6/�R�+���R�<��� �I+x��#<ͧ�?q@C@��*b��4e�qX��W8�?�	�',P��7G��uw���U�
.5QF�#
�'�I���4��HB�&���.�y
� J\H�S�(�y�B�"Ds��2"O|�9f�6�|-@�k\�-Z@x��	����ؐg�5
L iQ�Zl�Ѳ#�1�O��	�O��� �$��6O�0 Î��
�H�B3'�D��B䉄@G(��`�~:��A��2R�lB�Ɋ
����d�?�
h9�O�{�^B�)z�ܘ�ą�h���3��V I&B䉘#P)��)�s����� #���J}����PEKQ�� r昬���"&! �H�O��ې��O(�d0��S&G``��vdߘG'z�S�Ee�C䉭Y]y'
?ѐ�<P�B䉴$��T�-�&ݴ���/J:�C�Ɍ'o��K�	+U�	������C�I�u@y��Pa/��)�����=��O�I;�?OL�
�~�T��g�Fh� OM+I�*�{rfNg�	��I�n0��(*�i>��S.J8uf�5��m�0m��ȕ@;�R	�h�"ʧ\r�!�OP->�d=rso�Q��DG|�@�?9����'=�V��D�Ȗ-�HZ4�"؀����?����)�	��"������kB�:�l����ey�f&�νHŊ�8<(I��e��D�O����O��?��'`H����h԰�RF�k�d�y��?��r�Dx�B�!�@+`Z ���W���'���xb�ĻJ���+C�Z�� �xd�X_v�4�'>,�	�_vjӧ�9O\��*݈r6��&�S$��8�AƄ\|��I��| ʱ�O�'>�[G��+V(9W&���~�kr �u��'T��<��<ɶ�٤n_q���F�"H90�3w����O�!�O�ea4�>)�U?�'��lY��$�Ϲ|���!j�OV�f�>��N�O��)��/�,�hH�&��&�*%�'�bȊN�LqJ�x�!	9}��d����	U�Ae��E�I7�UؔQ�����/}�?�'_����!�XJ��i�
��t���O<�RB�>��y�&����6Vվ8�!�G�y�@�,!�@YkU��<Q�@�u~�e�G�O���  �E.)�n��E��Т�l��	.u�,�S��'" %��'�Ρ[�/�C�0	���J(�.-�������_9`ip]�R��+q�Hm��`�y�!�D��pL�i!L3Yj�ʥ��f�&�'Hb[��0����'��iY��0�lA�!����*8p�~X��4�?�H>��U?c��s�Vuc�> :�%	�K�a��Js�x��)�S�x_v@�2%2�-���V�Ay(B�	�"A�����:r�t�:����W(
B�	�X�he0aF׈u=b]�SDT�S�C��p�x�
F ��C�2�����B�	� "�����,6�$i@�Ф?�pC�	�z������0�Rk̂a�XC�	8|�h�(�.K��Ԫ_�)�8C�	b������9�	3��<�C�ɉ)(�p�D�2�Y��-��c�*C䉌sK)�3O�*O����b�4#?Q���?���?���&��t"%G�2j����N/ME�����i��'\��' ��'1�'���'*�d�1&a
2��D�ؕh��h��o�$���OF�$�O���OF���O����O�%Cf	�R�tj��Y�P��� ��צ��	��4�������͟<�Iߟ��	��� �:G��I����B�����9ڴ�?���?I��?���?���?9��L��Mb�DV�'�\�g.�"'��@1�ig��'���'3��'q�'pb�'}�pz-V�h~�9c�j�<G�=���c�����OV�D�O,���O����O��d�O�Śp��q�j:W��F���ʦ��ӟ����`�	����˟���ٟ��>K�R�§ؓd׮	!%���M���?y���?����?����?Q���?�d�ߚ"'�廖�Ke��������'R��'Mr�'���'�b�'���D$z �����2 zR%�5�6�6M�Op���Ol�$�ON���O����Ox��6�:�k��i!r���
���n������t��ߟ,��ٟ������	�s�6@�7��]����S֪��A�ݴ�?���?q���?1��?Y���?q��0��̪����IH<y��&��n��4�S�i2��ڟ��'�?�A�L"�^�/��6A2E}�R�,�	i�'H���:OZ�X�"�Dr������E.��S�'h5ON���@&~$�ٴ�~�� k�!��jބ����C
�?a�'������hO��n��	C,T@��á��,����O2���ᱟ���"� ��
��>~?�a�ӕzY|����D�L}��'R9Obʧi[�)@ �!&9��K��0�D��'��Ń&@c�O�)�?	��o�֬E;f�`��r�^��v��<�+O\��(�g?�R�����$B�E ����Qϟ���O��S�&�4��I���y����'JՍ��!`�b�O����O~�d�-$^�7�*?��O�	}�� ��S�Bw��;͖;u԰�#�2ړ�?�,Onc>u�e�ȹ"�tu�!lS.��ԉl�<��T�ؕ'Vb���""\����ơ'��9ǁz���'t��'��0�'qg�����U�Lcp�
�D�7;���{a��Zm�'z��柰چ�|�^�db"��>`e��`��#k̈��K���2�O\�D_�h^ 1�5e�)�lHP��¦��?UP�,�Iڦ���^5|TZ�k mjh����PM��:��U��?���=�d�����D���a)�(Z���0�v�B�$��D�O���O���O��9§'���G�[$H`�j����X��?��W��	zy�+e�Xc��H�(�2�p���^'B$Ap��O�Iޟ m��?���%\�9�'�|LKT�N�9􄰅gT�G��X��_�����[y�'��)泟0���=c�Xe����(H��9�����O����O��Jv���4N'����}�2�'�"��?	���S�)ы�:)�GJ@R
��S�ӤW�)��u���J�<q�'b����B�ɱ%�2��3�	<�L����J�(�����?!�GȤ~��p�A������D��ڟ�x�4��'2�1�\Q�8���C ?WH�=;.�*$��7��Ǧ%@�ڦ��'�<԰""��?);��?��刐"b�hd�@'�"N4r�
�O��?���?���?������1Nd���p�Iv���$`�_����?���?�M~Γ���;OzX��R�� }0��*�P�֎gӂYnZ��ē��'\ �8�4�~�()�nI��h�F�4�{�E�,�?���c�����;����4��N@�]�d R�b��~IrBݗ"B����Op�D�Ot˓���������0qƈ kD��X9_G�s�Is�Sm��ȟ���{�d�8�� &��Ҕ@��+��61�'�.�R�(�(9��V���*t���y�t����	����Wʆ�wL�����O���O����O�}��'��IPFЧ(����a眢
}����5�	̟P����MK��O)�����F�>�P9qT� D�
��'�l6��צݴvc�X��4��$��A���'pZ���a��W�tUHu�@�)��w(���<	��?����?����?�fa��_ع����3~�x�X�m��Fz}��'���'�O��(olb]�'��l��x�r�I	��9��F�l��0%�b>�C�m�>5T�H�@� |��@aM�.R�E.?����6,(��������D�9" ���5ꎅ���E�I�~�N�d�O����O��$�O.ʓ����<�!�A��T!��
�� ��<9�4��'r��?���y�ƛ8�0Y��'�!C�0����ܒl����a�'��%[aMw�O�S=8<8|��ʎ�an���͐�2l��'���'���'{�����-�d�ш#�t�� צ;t˓�?�PS���'.���D�{[^-!Ǩ�5!W�������'�'�2�G�a���4OX����� 0+�m^�ǥ�V�<�j��ӏ�~�|�Y��S̟��	��"Q+hA�IDf�8X���6��ٟ$��Ty�>Q��?y����I�"�"��3� R�B0���$t�	�����O�6�d�)���	D�0�F+oy葚�̉a5��sg��p�RE�O&�`M>ye$��t�y2��W�9v8)6H���?���?a��?	L~�)OBY�I)[�L�Cމ����Ƨ�|����<�ֲi$�O���'�R"��Z0$�Ċ��Cc��{AB�ws��'�JQ@��i!�iݝ�4�_bɟ:q1'�Z?'+�I��o��~�Y�'1������П��I̟���k�D!��ܨA���mפ2��GD��ʟx��Ꟍ&?}�I+�M{�'�tT9ԪϺl4h=B!aO�AL��pƺi�X7m�M�k�*dG�l�J?�W�U�'���H�t"��)Ej��tyr&JUr��_�Jy��'�bd<ObD{���+N�1`קڑ.�r�'b�'`�ɍ����O���O(@�B�7S�藊 ���n׶}��O���'
B�'
�'�h���Ȍ)�,@[�ziAC��.���[���a"�}�h��|�G��̓M� ��&��Z�N�#�ˌ�\f	�I�����	v�O��䍄P蠹2&ת�"Ԧ��	���>���?�$�i��O$�	�q�d1��*�"z�p9`�ɞCJ�DZ�aZ�4{����&��&>Ob��#L����'s�	�#L;dH����	-�D�B>��<���?����?����?�s��>C&��R�'�]�&A���C���D�J}"�'���'���~"��cG	KB'P�>�X�� �
u��I��	E�i>5�	ӟ��kպcD�L���B�I�5���n'�$lZR~�??����䓋�d��(�"���� q��ؘ����j���O�$�OF���OL���W���H�? > ��ܺr��k$&�o�6��>O�7- �ɔ��D�O��|���2��FP�Q�3־<�Ի�o��!�7�+?�S/?l���|��w�JDk�l�
U�0u"%�\�7)����?����?����?������TM�8`���ᶌYu�~x���'���'�8듷�D{��c�h�gi�LХ�%��NJ ����,��O����OZ�{��x�8�6ڮY�	
 ���h�fr�u�,m���OD�O���|����?��-��R2���XX,Hf,DR��z���?A/OL�'t��'�Ґ?]R��)*���D׏$g�Mڠ�<y�T�@��4l��F�/�~�DjȢY��D�����,�F�X7L���i��� �����O HM>�ㄋ8�p�넷�|�Q�%N?���D�OD�d�OV�$<�ɰ<	��'ި��rɆ!G҄�#��$?X������Ϧ��?�#S�x�޴>�.��F�W��P�J
,�<pr��i97�܂ZEf7�$?���M�U��	+�P>�X�gh��Ql@����z��^���ޟ(�I�t�	џ��O~��c�?B��;�fS^�9B�R���	�����K�s��2�4�y��<�>���@٬p������?���Y�'�O�u��i:�$N�.�$Qa�N 	,�ш ��v��L�&� ��Ɏ��'��i>��I>{5p�Ã¬v���8|�]�Iޟ����T�'Yf��?����?��,��FX��#UlF�4�"�B�(��'�Lꓶ?!��0~�'����D��BF�<x��A��T��\��S做xP)�	3?ͧ=�����y旼�Q�B���7n��#����?i��?����?!��Iv��
A�,(����c�ʷg' r��O���'R"�'�v7;�I�?a$��^
v�SuN�P3�	�P�������ڟ��	9=���md~Zw]�5�pܟ�����V�6E&hR"�*c�/�$�<���?Q��?����?�х֒]��0�a�� 6FM��d���D�u}r�'O�':�ON��0 �$��{D�����9{`˓�?	ݴ"<ɧ�L�6��4'�	���X��݆vqDa���s�2?A'2��$Y�����@��J|YE�~���Y]��I���')�'�B�'F�S��O���G�U}�=J�`�?1hR�rc  GU*��঩�?��X�$���t��k������xA�#��;k�*��cNP�I�'����?��}B�wJL��/#
�����r�Ա���?����?a��?����Ȍ(bH�!
D��uM�<.?n�B��'�b�'���?�� /�v�䒯C��t؄��8�&�H�E���L<���?��� �fx�ߴ��$�%r�R���`��D���n�^�0�Q"É�?�1j4��<�'�?1��?gl�cA��2�cuh�"�����?y����F}��'n��'e�S�/� l	sjG�{TC�	�W$���I���m��S���\o,q���M~�(��;����$��$YR��'+�D̉៘2��|R��Z0`1(����:���/@R"�'&��'C����X�����.z��آ���[�ba�C��[Xm��O~��i3�O&��'۸6͟�A����sE ^��]�F��#�
�n���MS����MS�O��we����N|���ތ4�~��dE�c����m��Д'�B�'�b�'&��'��	V��y�k��PM��D�0E�H��'���'���'�7�p��qUj�[~�k�I��jU�����O���6��/�)ٿr2�7ͨ���4 ÷$�2qf�d>�����O4|{�/W�~�|�[��SΟ��&��2v`B��� ����T�r��؟x��䟜��iy⋷>)��?y��MG�m�OK85X��J��Cs��p��ȯ>ᖿi*6��j�	�Dv:�i�&�*CU�qp�̗+�ɖ'�=Gd;e�8K�����ܟ,K4;O�7��Vt��auF� �N�S�'���'o��'S�>%�&+Z "ҋ�N�\0"�a�'����	)����<y�i��OH�	4m����W��	S��d.Ip�D�O\�D�O
�@ ep�B�D���S�ǧ~��ŀbR���+,��@��b[l�Ijy�'"��'���'��'g���� A��������XG�	+��$�O���O���D��&�RݛFb�+N�̰娋4@�n��'�b�'Vɧ�d�'	2K�*m��	�Ap���w�ӌ'y଑D"��M3�O�䱰�V��~"�|[�2�mU�Zm&��cI/i����Õ����Iޟ\�I���Iiyrá>��QS�) ���x
l�S�iVF��tJ�S �&��UC}��',">O�\�#��F���a� r��}W�2_�6����O�<4�Q>]ϻ@�R�I���w"Y��O͚\�E�	ݟ����$�I�X�	B�Owj����L.�%�
�1`�����?��`��	]y2idӆc�8����\ҙ�7��$������)���O����O���2�z�Z�"�Hu�&�ĉ��rEB7 ���:g�F��k�	sy�O ��'��܎z��d��kʈH��4r��܆E�2�'��	���O,�D�OV�''
�X��ǘ8�`�rEC[
<�'h�ꓚ?y����S��\$���ÁT�9�"�CDۖJ�ȽA-R�9#�֗�T�7H�$3���;@=�ɃA���P�B�4T���O
���O��8�i�<���� 4��+�<�e7F�4z>"|h�'��1O>6�'�	���O�[�O@�9܀��/v�Q��O�$��L�Z7�#?Y���0�&c?�c�ʒ +��)b�hW�+ D�{'�O.��?���?a���?	����)ڏ��K�C]]�]2B�e듞?Y���?iJ~R�'��V4O6L ��\߆���n��[�,ݘ�LcӼ�lڵ����4t��ٴ�~,'qX��q_:o��<c�F2�?9��S�4���ȳ����4�����	f�
�C��|��Zӯő����O����O��L��	�����ٟ�J�ɖ� � HY��I5�ܚ��DW�^>����lZ7��Db(�7&��}�~su�E�o��P�'�����猖4��eK�O�)��?���j���qE]!�I)�bɠ��@���O���O�D�O�}z�'M�l�sË<[�,8Q�d]3��@�/g�IR~�iV�OR�Ɋ�iO��`s��:?�zPz�̋?�\�$�ʦ�Jߴ��k�k������D�ّ~+����<�2�іG�@L{�B�p�&��2�|�R��������ޟ�����`2�j��,�9��	��)�~e���Z_y�F�>����?Q���'�?i薮u��d�ec� }��Lpw��35��Iޟ���z�)�S�?T��2�DN�ך�JD�-�R|���#F��k[
�p0n�O���O>Y(O�%3 ˓i�y��^ߎ��df�O��$�On���Ox���<�D[��̓S+v��G�G��:�r3%�!�|���>�M���>9��?�'I ��t*�oM�䘵��(��|z�mJ��M��O�������t��D0�j�����-F}�����EM2��b�'�2�'2�'�B�'l>�:��;���	BaN�B��$[��Ob���O��',�'��6m*�I$|b8���c=aH�u�)�,��O��$�O��ĎM�7�(?�;Kb&}q�T=Q�Fx�7f!_�L9a���~��|R]���	̟��������S�W;�<�TJ׼(a�:�ɟ��	Pyr�>I���?����I�t��|Ia�dr�%)��8�I���D�Ԧa�4Ig����1X�I�]��5k��?"�B�T@^�9����������:+t����:GK6��g$�	���⷏��,�p\��������E�{yr��O�eq@��&@2��N�<H���'G��ަ��?�vW���ߴc���x����e�6��4Ƽ	 �i\7M���6�&?�� ���=�	°ڐ5�v��0��X�6�V8S��]�������I�����矔�O��i�
b�:1�§O�NV(#Z��	֟P��q�s�X��4�~r��=`�1���8$������\��\�I[�Ie�S)Ȩ�o�z?I��$�����1h��uB"ߟDb �ˑO���3�Ĩ<ͧ�?)T� 83M��6$�E� =x�	β�?Y��?9����dAG}B�';��'#�ss�]A�� �$L�#�5�DC~}r�}ӎ0m�2�ē�r���K�W�H�c&�A�$ �z+OV��e�בX2 �Ә��("����<�&@Bb5vuR��O
�0�`FIȟ$����@��џ�E��6O��Ef�(w�9уBܭV�>��%�'G6듕�Vަ�?��'"�hѳ�"� ��hT�G5LD��H��?a��d����B0⛦?O����2�����u'�3hp����@(v�11�$����$�O8���O��d�Oj��X>\�f@2�\"���0 ��cz��b���ğh��ϟ�'?�	�m�i���R�ND�9cǟ>1"���O�pnZ�M�W�x���.�I��ݠ5��c�Q`�ы=��c�H���ԣ:{��#�����O�˓)onP � T�v�,��9*�)uN�Οt����T��ޟ���ryRk�>��g�f`�cN�43n �y4�Ɏ2f�ً�;�&���y}��'����On��& ���˅Vk��3��MD��搟�If�T���D�Iu��r 쌖);���s�Hp@��O����O:���O��D�OT#|�CǗ2Y���K�v����V�����ǟ��Oʓٛ�$�!�t|���+�}���۾(�'���'#��F�ϛ������Ǧh�tu)�&�	�
�r�/Na���V�ON�OB��|���?��?]Ҽ��&щc�.�T�Ȳd4!B��?!/O�Q�'�R�'��?9kQ����x���L���7 �<	2]�,�	֟�$��O�*(�P/ �O�X53A,4���Pi��1k@p�޴����ܨ�'��'lp	���0"�.��WdNOx MxT�'�r�'?��'��O�	/�?Y�/�%r�Cu
�?j�����P�	�<��4��'����?��ʎ-_4��1�Ă"iF�t0���?��T�h@ܴ�yR�'�h��@IE�9Ol��	),�θ��MX�=N4"��O�ʓ�?	��?����?����	�!+��,�rBH�<H M*# ����D�ON�?)(�4�y�T�>n�����ŭKԞd��H�)�?�����?a���?�%���MK�'}43S��O��c2	4�Z�3��'DN����y?O>�-O�I�O 4����&^�H���0X�����OL��O �$�<1�\�������I�$�A�,V.^�L�v�[�9]�8�?q�W��Jش<���L:�'F&�A2C/7O^@�ȗ�Fl���O�q+ @�R��):Đ����5�҈��<1�JF�x�d�B`D��R�`�B�@Tǟ���`��矤E��2O� �����Vj
`j��
&��	B��'<���?��d����d��~���eF{��DA�%Z�3��i�3��Of1l�8�M���i�P��Q�iW�ɵm���˔�O2���cӐj�B�[��.t�#tK�Iny��'q�'�b�'B���3�2I�9��<S�Ã�L���,��D�O��D�O*�?uh����:l`єcm�L�f-��� �<���AsӨm%�b>%�����C.V8���
�〈��jTe=&|:��Ayb�Q\������'_�*��a�*�������F�F��<���8�	ǟ��	�'<���?QGo�=��,�u��R.���n�6�?ჺi��O��'�^6-�����p�^�RPM�
>T��@�ꖰ ]���c\��1�'��be��?A���4���D���NT"	�!-Sbqzg�'e��'���'q��'�>Z�nG"|~M:s��z��0��Or���Oy�'���'�<70�I1h���ԊH�EFد �R�O��D�OT��H]n��i�񋱋ҩoș ��7ؘ�b��E�*�������D�O����O���D�Z.����J�6sۆ�PĈ�"T��D�O��3���� ��ҟ�O�L��"R�!�$]��#ټ�<�H-O���'���'9ɧ���=j�`��Բ3���C��4D9��F��	��7�Rry�O~�D���>O���& �J�<�`�k]+e!̕����?���?1������$�ǟ����"-j�1�����IQı�gk�O����O��oZx�8����Mk���e"f����5Yn ��蒟*��dӢ��ubf��f R��*�d �Ο
T�a �50���0A���d�n�Pr�'�I՟T�	��	�L�	f�D� V�0�GQ�ř����8���П�����\%?��	��M��'Gd+1H�6L�)+���.#=�e�i7�S�I�?u��?�a�n��̓l<aU��0�yz��йVH��8�Th8�0��O�3M>�(ON�$�O���"�+���#@|�����O��O����<95R���'2(ӂ3K ��� �W����ɔ�q��O.��'R�i_ēO�0Bc*\[��)��z�xų�'�� �2Q�A���>���៞D���x� �/������u����v)�P8�$�O��d�O(��'�'�y2+)h��Q#腚0���b#h^$�?�[���'v|7>�I�?��ak� 
���Q)��7�t�@�!L��	쟌���3�XnZ�<	�Yo�鲐 �~����;&���r���)\{��@fTW�iy��'���'�b�'E��C<f�޼x�	��i��,�F�P6�I.����Oj�d�O$��h�I$+�aP��@9|�A�K>-�>p�'��7�LԦi�O<�|��BٖY�
��go:]�b��0p������O~"��a��9�I��'��	�lR�I��ӻ9�8���A�D�^���џ(�Iϟ��I쟘�'���?���J�rhb���1��xVI��yһif�O<��'�f6�������K��س�l�*3kz*��F�CU�I�E��U�'�97��?�}ڞw�8�ʥ�F 2���(T��_tT���?���?A���?y����,�
�/�a8���$]'�|����'�2�'jr듿��{��b��1�NH�(e��7�K�����.O[���Ţݴ�° ���Mk�'�B�M�t[X�#T�*$t�K�Ɯe�1ib�����R�|"W��ğ��Iȟtk����$����C��qyUi������xy��>���?����	�'�<�6
ό!7td5O� ��	���d�O���;��~�ƈ��3~�tC���x�,-C�A^�k�H�JtC� T�����H�O~	�H>��bP @j�a���=!k��'L�!�?)��?����?aN~�(O�����d�Py"aO$!RJ, ��,8`���O����M�?a�X���	;��U�+L�p�R����P��ݟD)�ߦ)�u��ͨN�i4Jso\����U�-�*m��OM��x�'���'���'���'���6t`���ba2f�`��%�B�(�'�"�'�2��4�'�j7�h�tc��!B�Q��LҜXC
�6��O*�d9��"����]:�6������cW��^�:ŦM�mx��sc�Ope��D��~�|R����ПT�㍑�jv6a��$�$W�q���C����I� �ILy��>!.O��$T�b��6Md���<uJ�㟔�Ob���Ob�Ob��ᅿI��F�U��\�!��<�G�`{��2�4��O��,��y��@	�U12ʚ�5MJ�k&BB�?���?����?i���j�TP2:b��������}�d��O��'���'G061�	�?!���+U�&U�0m��+�H��fϟ<�Iퟤ����|m�w~Zw`�t��֟��RFbϢ+����k�1y�d�&&�Ĵ<����?���?Q��?��:(7tɴGD�}:bH*&IL���$�J}�'���'���y�EEG�,X�A��� ���7d�N��?1���Ş;�v��0U~$H�L^!d�ƭ"����Ms&Z�,�h�7��d5�d�<Q%%U�(�(L�J�<~�,)���ܠ�?���?y���?������r}"�'��Y`��$]i���1�$���'�d7-"�ɻ����OX��s���0!-(�Ui�NGPD�h�S��% T7�$?q��C=2d �Sy�Sڼ;�aN��Y
OB���,�~���O����O�d�O��$;�g�? �Ic6ˁ!0���5��5yc�'���'l듒�$o�"b����G܄m��aq�rhɖ'��O���O�+$�p���k"�iG�^-'�����>F�������	���	W�IEy�O�b�'T���"(/�dSE(R�=��LB#'	��'��	:���<������b� �eޖ5��cD�ӬX�I����O��$-��~*�c�u����U���4��=�.��"Yv��7�ŦI�'��4�_i?�M>!Bd�4�p@����{��1Q��#�?���?���?!O~�-O�Q�	:�:�SN�j�r1�R�#/�����<��i*�O`1�'���Q�vy6x�U댤!���p�.Ća^"�'�dX�!�i`�I��vY2C��
.y��5���%.��2��2*�_���	����I��	ğ��O-�p �O�?P���ANf�B�Z�W���'����禭�E��=QDV�hӮ��%�.X�L����H$��%?�Z�"P�����#a7��h�'��c�����'��6A�I?1L>�(O�I�O��x�J�"��0����d8b@�O��d�O���<QSZ���	ş,�	�B���Rr�ìb��)A׼-O��?�gU�h����8%��Bѭ'v6��T��d��Ȼ!C�iy�� Gظ÷i�i>�Q �OL�I0V<������2�����'>B�'g��']�>�͓i�L"T,N�g�vQz5�X�<�����-���O��d�����?���YP*�DQi��q�#��yv١���?����?A£I��Mk�O��~w�SD�$j�YihQC
V=�h�&�L�'���'&B�'���'.�2�S|�����ɉ�f
���6Z�X­O��?�������c�(@b��#h�V$���B�f��?�����Şp��,󁅜�N��x�g/�3K���XSgK+�M#�O*�[`�	��~|�T�t
�9`�8@��Ü�2�����Dß���ݟ���՟��	py���>a�bc�)���'wRy��))�nA���ě���Ar}�'2?O�2'�ҕUu��x�C�c��-Hq䒤i��V��`R�&�>�Q>AϻB]&e�U�ͭc�-�o��Zf��	Ɵ�	ƟD�Iߟ��	y�O	T@\!0a�`�Ça�81Z ����I����O
ʓI���D��g��+��dK~-1AOJ7��'+B�'��N��\^�v���SG�ٵv��+��ݤC�2���(ߠ��Y! �O$�O���|���?a��Zg� �4�]�X�rA:@��?ǒ����?�/OT\�'���'"�?Mb@R
f6�Ƞ&�'Q�b�D�<I�S�\����D&��O@���n��)���:r�ս/�t�$Ԙ|�r$��4YO�I�?�3��O��O�ev�­d&*D!����`�0�ժ�O��d�O,���OƓ��˓a��O�0� y�`�ĵdXjU�L��	Ny��c�V� ��O`�@�!�v �WEBac�؀Bz���O� z�$zӞ�Ӻ�u�T���Ԝ?=j0%�5z��N��`ς�B���ONʓ�?���?���?�����Q�)`���
ܛa��D���z������O���*�DX�QϓRv�b%jA�UeP,��X��؟p�N<�M~�7�^)�M3�'&��#7�	1W>�-��V�H!��H��s�*�Ń�O~��L>�-O���O�s�)աx=���_;rr�%;� �O,��O����<�u]��I�����'�2�S��!
�q�Ƅ�7sM��?��^� ��ɟP�N<7dt]�um��I�H�f� 
E=�ɵu�&��-'��|����OP�'���s$/-}�5���3���q��?���?���h��ɥ��9�_t�v�����Y���w}�[��ܴ��'�-�28��K�!��D�Ш�7}��'��l� |0Ɗn���ag�P�����ם����c�C�b�;h�2	�Od��?!��?1��?���^M*X�qC ��҄n-d<��+O<��'�R�'8"��D�'?^�C��\�L���'ɱC��e�6F�>q�i��6�8O1�4�+��W$���k���Vg��D-�һ��.O���9�?A��;���<�ƈH7�&��&pP��咖�?���?���?������H}��'jz�95j�0ij�C���(I�:O|6�&�	�����O���t�A���E��X��"��s�N��nV	#2x7-7?1e�Q:YE��|ҝw������я<U"�s�@��b����?����?i��?����R����ZpFlRB@a��m�S�'���'����d�˦�<	TK�3d���C�i��=ÐL�e�� �����8�+�ڦ�Γ�?�h��KĎmH&f� L�޽�n�#P@PT,��d&�<���$�'�2�'�ZqP��?)��ԩ�e�yBx��$�'�_��a�O0�$�O��d)���X(o0���'�z�.|�!ty��>���?M>��Ni s�S�'/*���
(��HА�2&U��iL���bQ袟�'���F�J^�����#��
��T"���������	���&?�'���S)�$t���;VJ<٠�1v��'��a����O��ܡ���R�*��4�`T㗩6��$�O�d�	i�.��i"�ʁ���T]��k"CȘ]��b�E�)�\�&ޟ��'r�'9��'���'|�3� ��H�$?@�<ݣ"��/P b��Ʊ>���?I��䧂?Y��iA�$J1��1W+O�Pt�*E!-5�'��'���'��$P�^m�F6Ob�Rv�(.\,Qu���R�h�Oj���ES�~�|�Y����Ɵ�2�OS ��	$���J��2dYӟ ��֟��IJyΨ>a���?	�bڜ�B��>|&y����!S�������>A��i�N6�r�	�e�FՋ��GmZX&���$j��'~�k ֓Y��i���Aҟ�i�3O�H@A�HH�f!G��~M���'�2�'��'��>]�/�fd�� �\h Qa�#S.V������ ?�ڴ��'���cɕ>hn)�6)�s���EDv���'��'��]�w�is�I�y�X!U?�
�f�XJt,2 CNs��� -��<I��?Y���?���?іI�KK���i�2	hVm�!�У��D�s}�'J��'9�OK��>s���3�1b�Y��ͺꓹ?����Ş��Hj���"+��;%J [�/�tC 6�,?!�>J���s�Gy��o ��s�"8T�-B���g�R�'G��'���'S�	���$�O��a��A+U�`,a�&Ύ��͸~��n�M����I̟��	�<�$�((�����I�ʔ���[�c�.uo�}~rl[n�<G�4>�*�J��Y#zMhi�`F�d�A��'?��'@B�'���'>�
�N�pz4���D��"�#�O��$�O���'�"�'6�7�:�I_W����	�*�� 7n�t�H�OL�d�O@�d�-��6- ?U��(��(OZ� H��	�$R�(D.�O��M>	,O���O����O�}�Th��wp|�j��L��d1��Oh��<Y�P���	ܟ���X��XYNN��gC	KS�rÀ��d�\}��'Yb�|J?u����z��s���c� i�lP1n*�H&��0B�I�?���'��%�j�L�!L��eAuΑK�}�E��X��şp��ßH'?-�'�z�
6����Е9�M8�oFD'��'r�p��㟰Z�O��� :]�Ɛ�)~<`V\Y�,�$�O~�R"�w���M���t�柌�HE�0�H82؆c��J���'��IΟx�	ҟ`��ǟ���}��Sθ%�t�.���5a��=��I䟀�	�D%?���/�Mۚ'NJ�ŋ-v]�=*��b�Ɛ���?AO>�M~"�-S��MS�'v�0��x�)S4@�3W����`9g��O�8{M>!/O���OL�"4-X�)���5윦?z�R�B�O �$�OL���<�U�������	�}sڑ���K*M���@����z�H�?�_��ڴD���B1���AX2�V(ON>I�'��%&�X�8�c,]�V�d�H~zC���S�x�Ы�<@�f��&JC�|�B������*v=1��2t�\�+ƭӥ;�Y�`���q��HF�h�Jr���5r�]pb�(@]�AS��V�K+��[�9+�8��?o�Xua��OU�@�3b�e��v�S�_~@���#F�Zl��V�Zah0��*F�T5zO�>����S �c�t���S�mݼX�A�O
1I8��&(C�C�U��J�(!�T���WTГ����X\+tƚ?X#�(��0c$��øXK�I�t���$|@p�qg�j��;5��5M7�h{B�2�h1��h 7Q��%G��4� 	<D�n�SP拑G\�	��L4�8��f���-5  ��i�N\z�웩nO�se)�f�Ȭ;0f��d��i`
ÓkȤ9k��5"�	Se�/Q��b�ɔ?)����玚;xM�����*�4	3,��h��	#��94���"qˑ5�j�)e��-L%`� � 0$���ʀ����SLQK�}s�jՆԸ@���H.�L�!�2�n�Y;K�Cq�&j�y�Kɳf|�������	�
�k�J�[�0�E
��_�t����Sw����I�#�|�p�����c������(e�<�a����͟��IL��#�:�ǉ�W�j�j�*]?E�2���ҟ\�'|R�|��'}�/{M�����1�bH5zѲ�i�H����pʞ'R�'����C�~��V���y�MØ<I\.k\d%���?H>����?��k_��?��O�lAÍ���\�8ť�-� u�'���'��"�'`�]>�����	?6�
dI%�w��iT@l@%���IԟX�UOIԟ�$��өtD�XƯ�����
�����1��O�]m�П`�	����	���˛I��8�J�%.����挚j����OV��͢&J��t�O� �i��?���>}�� �WC�(Lb�'��'Q��'6�]�P�Iӟ�2V�U����Be�^}�4��
ҟ<����P�S��B� �y��'�yЀ��¹t�ݢ*�eXexӚ���O��D�O�'
��ʟ�̓Sk��dBy���d�n��u�?� ��2�?1���<A��?��|ʸ��q�J*ƽ{Rش	{�����?���C&��gyB�'��'1�a��F^�
�6���C�7�"Z���u�̛S�w�|�I�P�IC���>ָ�lB�5�`� piЏ�?��S���'�"�|R�'�R�Vl����⌭7�!��1d��X��'�0%��'bb�'VҒ�� ៼��!c+_ �m�dDc� ���'7���x&�����t��Ș������ۭ�zͨE��b��Ί!F@����L���T'?ݖO�"+R��<��!Η5&�h�P�L�?���'��'���'N�8J��d�.��AA���@�9#Q	Ռs�2�'��O��y�'V��'�?���?-��A��f�:j*D� E�UzL>���?ᣌ����'��)�BY��9�^8&�J����r*�"�yr�'�x6�OL�$�O��d�Oy
� �"g2~�,PS���KA0}Y��'p�ɟ��	X�I�D�^�]q
\���Ƣl��py�.��{ARը��'ym����OZ�$�O�%���	�Qʔ �K�R�C�GT���O|���OV�O�ϒj���O8ݱ�EB�R)�)SI#^a�PB�ݦ�����(��ҟ��K<�O��$M�R� �d��<��ƶ���'I�'������D�|2'gEK�ؠ��EL�:a`D�Y��?���?�,O�˧��'�����G�d��K懡�J؊e�|�	Xa]�%q�Ob���O��z��b�O�|�c�$P�v�4�9�%�O�˓�?����'�=O�M��W%J�9�N�F���!��'��غ�M�!��d�OD�4��������3h���U��-S4��DA��?Q���?9�B�'��I�c�`(b��HO�\�1�Բ>gX�a��^	���?����+O��'�y��ڷ�:.n-<�0���VW��	W���?�*O�e��>w+M&.��ݐ�J��Q1+���(�I���7�~�T�I�����O���r�	�D�8������S����C:�Ĥ<���?�O~�Ȓy�D�=K��EP KO.1�f�[�>��$�,O����O��d�O��D�<��-x�1J���C� ���0y���O�ʓ(?�Fx�O|��:d��6a�tA+"5�
h��Q#p��؟���ڟ������$
�܉�S���+Ε��FL&R��˓�P�Gx�O���'�R�լFܱ�+Ԗ)+��6�J(@^7��Or�$�O��k�)Z�'��VDԅ�LB�f��z\���?qH>�����ϓ�?���?��x�0�Q�R�x� �K/�?���?ɰ�xʟ4�O���g�W��3�G>^�m+��<��OB��g��\��ןx�S�<ebO�a�0�SQ.q��k0����'"�'��O��Dw�Lȃ�KK�ҥ�+#�b�����O@�F+�S���OP���O���@��8��8K'�C >���R�bI�P��?1��䓏�4��D�Z�����O­bb�:�b�	��Z27O �D�OV��2�)Kl�T�'X�W�d_�U�U�Y'z��1V����P��U�`y�O�b�?]��_07�EH� �%u�x0��O����O���8O����Z���'ur2��X;��¡[(q3�ڹ^��5!��|�^���I���%?�Ɋ\6����.�3z���ĝ�WhD�Ɂ@��I����ش�?a���?	��K��$���x&͇����ff�O<���I͟���!����İ|�v���H dØ*s�����3ElI��
�4up���'n�'�"a�>1+Op}z�f@�l��)#���)w(��@��7�L�h��$�O����i�����O�؉�>�Ђ0Jd��Xӂ]ݦa�I՟�Iȟ@��O���?�'(4��"� }�0A3�L&^�<tz/OLʓl$���<�ϧ�?a��?�fӭi��A����Gy:iVϑ��?���?��W�ė'�RV���;f\���G4:i�25�і'�"�'6*q�S�'��'�s��P��A`�;��̋'���Jܟ�;�ONʓ�?�/OL�D�O ��}՘���&9v�a�b���9�8O�m���Od��O<����'Gs���X���D�@ 4�:�s�Լ�?�-O�d�<����?A�F����@֮���BC�����囙Z�0��u�0��ӟ��Iv�S���)�O�@���Irn �GJ
.O����O����<���?���$(������;>�8�sƘ9��xjg��\HR�'$�P�y"�'oꧠ?���?��L p,�1e��ܨH@������OX��O�-�v����'_�)U�J�(M9G��b�������6`aa+�y��'q
7m�O0���O2�$�a}�D�ej4J�jŨ?���[�%G�h7��'��(��yb�'i�I~��L�k�����T�F�{���%E!Zua��'�� t���$�O4�D�O��'!�ɠ,)hU���:A���ؔ�G�#+p)�I���IO�u���	�y2�'�>�A��M�M"=XV� D�<2�c�~�D�OH���O}�'"��ş`�3�8����V���Lh�M�Gydy���,�'��h��'G^C�O)��'��K�HӴY�ʌw�l8T�Mm"�'���>1+OR���<9�wd�,�"lP�L�,�C�3��I�*O���u=O29��>O����O8��,�tĉ�f��l+ B+>z�|���A֟8p�OH��?�(OJ���Or��͝s>ܼp$KD�9=*�3�(�$�b71O�	b$<OF���O��D�|2�}��D��CTTMKJJ�<7�� ��K���O0��2���O2�D��hI�D�)�p���18pP�H�
f��ay�'���'����n�~
�iu��)	�b�0����,oG�����?�N>����?1��-�?��O�${4嘭a�:�8QW�Ѐ1�B�'db�'ێ�q�'����~����?���!�h��m|��Q��iR�$�O����n���u����,�c ,��,ӻ�$�$�P?�d�OP�o����	ڟ��	���?��<
G���]�ƙ�u��q�'�R�'�$Ld�'��'���9�!���˼$�B<���*O����ʟ���6�M����?a��?1�x��'�n��!{�Xs�S�n`n����?qf(�'�?�N>�(�D|B�5O��D�#YV���f�� pY�1���	�;�4n����I���>��'N�>O� ��Sr�Ξ^[f͸4	�;e_ȩk��'��'G�E��'X�'��'����N������#e���C��E���'I҉/�$�OP��1�яk2�!T�_�_�����o�~�cz����<�B�͓�?���?1̟��s��¥
�e�F�ն#��kB�'�(O���O*˓�?i��?yfD��H���p��C	���8��ApJ�̓Z���ϓ�?���?YJ~R3�OM�Ȫe��i���K#PD+.O��$�O�O��|�D2a��Ona��؛�&� �K�)o���޹'~��O��O���t�O	R�dl�i�g�>Ƞ8���C3A���'i�'���'?챙�'��ɮM����〖-��ȠeJ!\#����O���W�%Y���OF��O�b�'��mC�AG��,�����Z.\��'���'�ԑ��'��'��)^�j��x%$D.q��d�$��.��!E1�y��'��7-�O4���O���wy�MG�e�`j�['Xs8�Q���?���?a���<9N>�-�~�(��2��й����A1������O�\m��D���T�	'��'tlp���� aˢ�9�����p���'�m��'��'��S�cu��Iڟ�3�E1eI:�U��!V��Ё
��M���?1���?�b�x�Oz�%� ����� !�Ì:���<i+O���Ս4��$�O��$�O�qW��!ЈP
W�0cv����O���O�x'��SZ�'6�<�v�اG�$;ӮԭȘ�K>��a7f���?���?�������T�|8�{��As9�x;�O��?�)O��D�O���$�d�O�找{۞�����
5%����A�+J���%ec$Q��=Od�D�O���-��T�?���̤0%aU:���0wA�O��D�OV�$�Ov⟠Q M�<A���~d�.lr4�$��i��Q�bce����̟����?E�O��'/"F^j�a���8B4�!āF�D���'��'��P��+�i/}����x��:��� ��E3&�?i��?�Ā;�?	����i�O��$�O�=���̒e*�i����N ���1�>���O�ʓL��"�3V�x$ f
��!��>$�D����8����?��i�b�'���'U�8JA+�ɐ7#�
q�r�W�3�ZXIN>������'S�d�'6j�yQ�J��3eŨW��1�A���'j��'f��'��W���O�L�����N!�%j`�R�XS� [�xS`G>��|J�ƄSy�ቀjN$���iFp�z�x��CI�%Q/�N4�g+� �<T���jJ"��iu�b���O|�$��O�ƭ"a�������dûCt�6_������?���JO~����y�ɜ)�T��,L1b@u�&LB.����"��8��(��A�3d�T��
�'�h��n��p(飧NG:��p���]3f�e�O����[]�1���Z-�	�wn�A��EP��i[���`�c�>��	^uT=�gF�t8����ËOL�EZ�M�s,�`��Sn"�ه�W�?��$XfC�\hV��ɟg嚂�J�o"\L ��3A�H�A��}��h�j�<��(P�B��	��:��|��C�	|(IPC��i�Fq�6i�2������
}b*M�#�]����	� i �@1�AԤ?�z���ɜZ��lZٟ��	�x�'t�&���29~���*R�i�|����5O*�K %J។���Mk���M|�>�0A�zv�rB:,.T�Ӡh��.v�����Obq�� �
8'>c����G?&��jp.�HL�0D ����$X��'=ў��
=bob ��/�-q�
a��\��!򄎗_�"(��e�+i��P���1:���p�����<�֋�%T��Jс6���� <@]sR�i'��'K�V���	ܟ��''�r�Q�Y�f�b��d�[7;�(9�U�F�V>�	k��t��[r��^��9o��R��P3�VXC@�Y ���'H�2�4�����DC>��т@��$}
��(n�,ll���'����O`�A�cm� Wƪ k�X���P��'
J�a�O>Be�]���.v`QN��@��O�ʓ,���X�Z?�I�����O��A�voĸ4�H�ǇD��d�O~���O�0�f͞�W�JE�JK�{�m�i�S�C΅�[��I9Nj5�6��9Ӯ�U���ò�������eq�x�fQ�h�4�)2)A���O> ���'�����DL�r�*5��g\bQ��[���JX�l�e���G���F���TD("��2�O����=ۜ�q�M+Z�$�v��3\�DJ�k�+�M��?O~z��M��;M,���.@�ΥQb�
�!�R��
�Va
fK0�|rN|*�-`t��Q���, ���sC�~}B��+X$�fj[ i}��������i�D�F哐Or:���lA��+�����۟ �4�?���	�<7W=�En9u���I�ŵh���?I����ō�~Jp�B�Ɛ@׮̓��I �M����O�x��G�>�=i�OĘ)I�$����ON���O^��D���IƟ���oy�'=��yKs�)5T$Ը�O�"V��O�P��k��q�&��?O_�\�CG@'�����/�dx�g��?1fdF(�DS���}�"�{uzX)!"ǲ#3"�Q(R/��mZΟ�P^g/b����<����M+�f�N���x���1���'�c��@�'UZ%�7�ԍO��bk@�"��T?��i�J7- ��|:+O�\1� \�ѳ(	8#I*�zAHT�8�m2�&��MS���?�������O\��z>i��'���f*�.=+���3F_$����
�[>:�9_���3-��>x�q�]?7a����M1��8f*� ����b(�c�P�������?���D\?�ۦ�T6�|��5�.	�m�0�$D�X��/�x�����N�/!�����=}2$�>a.O��'ĦU�����n#)�T8p�W!eKX �G�
"��1*O����OH�Dʼ"n��8�i�s�<�XP`�)p��e�%�p) pD�$J�
=ܸ)3)��X�0=��l#��OZ���'����!b���>������?�ԁe"O$���@�C&I�ǝ�J��t��'bx���6�N�rE*Z%1��˅���Si�C�I1u�X�2���d����7?�C�I�Y*8�PQ�؄
�X[͍qQ �',
�F�[��|�ƫ�%,�Rò{B� j�nW�I(4�.Y)�y��ЫNE�`!���F_�ѫ����y���%o�y��g%h���5f���yr Ȗ0~��1`�'h�B��U.��y�\��N�C��ƛf�H�!e+��y�'��Uڱ
�B�Ĉ�d	��yҠ����L�cX!3E4I�� ��y`ކ��	CD�/�tTa���2�y2�E��a��O]�/K��� d��y҈��:��n!'�^-�����4��
%�٭R����'��8B2D���]Kf���E�&���D���!�ȓb�ݲ쟞4�"Qj7K��e����ĬSX���H���c�5��bP�HR3Aľy-HMH���x�pɄȓ=p:]
�
�-����gX�O�E��E���5�U.O�����l��E�ȓ���R��&/\��e/��v�8���#�M�0�ϔC�
�pv���؅ȓF�L��F4��1K�{xJM��4L���5_�L�t��e��4U����ȓV2�A�3�I-f|�G&K�9�L��{PŚ��+�$�[�o@3㪼��A0ź��=aF|;�Mh��4�ȓ�}QGN̾F�f=�C�� m�؇ȓ$5�!�5Q��?z���2�D��fNA�Z�4 �K�+9ȓE�h�)��ܞ*Z y:��ͭ.���08KFςb>L�N�VL��ȓ% !���D��XI���?��Ň�)L0�Ѫ�'UuZ)��6G�8؇�o�ĥ���6�uHw
�D)��ȓs.���]Ҡ���ށ#����`�aL�
�M�v\�B�	��v�s���
=��lRe�)TB�	c���K���$�!�	y[B��
U��P��2Q����n�;i��C��!8�Z3쁗pڜb�O@�E�B�3#�R�c�#��X��/܊U�B�ɇ%�4��&P��3�.	O��C��$=�DW-
D4Q���~�vC�I �8Z ��7�@���m+6^C�2ЕhRdS�Ph>��#̞0C�	?3}d���=vp�� ��H��B䉕�$�����8Qb�!��ī�B�I�u]� P�Y�&��w*�3�C䉼{Px�Ĥ)�^Q(�%O$f�C�I:Wr�bvO� v:�ҷG^��C�]�1q�@#v�����	���C�<F��4�D���t��8��d@!50�B�)� �̱�΂N�ŧN�S�j-J�"ON� �S�n�"�[�)	L�Ij"O���MA�[���)hC�s�D�6"O�Q�q�EJ	���R�B�&X�P"O2��S'Q'#w1	t�K*M(Uh�"O8]�To©QL$ti�D�NHB�jb"O@<���%8Ih�m�	88H��"O:X�ԁ21Z�A�mE�@��zc"O��ґ�ڊx�,�� kD�f����6"O�E����r����4A��r�R"Oȵ��c��^�b�����r�8��"O>�!Ҭ�f��MۢO�x���{""O,% RK�P�\!-�c��"O�`�I1Z2��@�Oq�|Ău"O�mJ�/�2��ђW��K�F舄"Ov,I�J7�\i�c�b�||� "O�M	!b��1b�<("ǏM(�"O��:G@�72A��Ta�$��1�"O>!�o���CW�R[�$��"O�!��ЪI��ţ�O���zQ'"O�ha��U�sX)����;\Հh�"OR��Bkش;t��Y�Ο�M��}!v"O�}� Lu�H(q�\�2E�e�����@ ��3dqO>m���ȉ&D%��%:�(�YF(<D� ;�@߅x�D ���q��I�7�đs��]ⵌ7O�H	�>]� ���FJ+`��z�x���W��)�=�OJ~5����|*�	j�k^:f^�eA��5� �*��ܡg��s�eV8���p�H��;��f�	�����f�!�*��	bzQ���	�'��XB&a� �"睰b1Lu��3QUb=c��P2mwRB�ɰc4@���D#K�D9�
�$q�*��(�H4���3��� �R�i�<��D"J񟲙 2烼()�!ذ��f ���)�k�Li�@�h�x�#�>����!΄�B7�� e�Lk�៦|"84�a�*vk�% FN �`�}�O�X��?��%71����C�}S���7��F~"�Ɇ����ϊ[�T?1��/����Fk�	��(-t<T�Cg�;�l��DOx����'��=��gטnV\L�� �G>$T���;8r�'�vT�e�qp��b��L�
�s�(f�uI�f\��S�cC8)�#�RV����Ov؟��f�ս�UR��=��iYpÃ($9�Q6'ۦ����i[00�j�Cc�y*��M}��L �0�Adߧf����q������I�@�iZ�ᚌoV��O?���Έ!��E	E.I�t����F�(~瘠P¯X�T�l	'K�*hF$�'}��⟼�(�gX$q6a�(8��r�aօҦc�t��B�; I�H��I�S
�<��N��}R�%PPL�;��3�	�z%�:e�8�� `�9��{��K�ļ{b�^9�a�SÜ%M���ӦY� 83�M��i��I�̴sBbޔ=�]�c�\��yGdݡ;~z�KY3&�T;t��0?)Q)�#$���`�
�<�~� 5�82$qA��͘3���í�S��C��G[Ќ������OeQF�Z��5̍�Z���6e�2�� ��ɫX���I��Т��!,�x�JF��l���1LũW}6��QC�����';�X��W�9����ڰX��l�'�r����>g��'j$��⏯Dg�%?���*�{!,tX�j�)gbh��#D��:���U"�i�-��\Z�"�>!��h~�7JЋ���0��'r� �a}�u"���v�U��C]�/�U����	�&��m�f:~8�4m�6gpA IT�	��q�S��Q�E�'WA2�" �	�`)"��e�
�%��eƁK5�>����[�����On<��l�&^d�8�B�C�C����of2ų�f����?�0�ԓ2��QX��H��x�!Sb�}��B�D��OH5�h�&+��O�nO�[@�-���JD���ԑ�!��� ��&՗3p��9��Y�/H�	�U[��c�n�)�'��H2���
q�l�1C�(q���ȓ !�����ī�	����t�<��I�����$F�JB(�q�1b��\{S/_#8�!�$�n� [5��|��1p5GJ0M�!�d��T]�*�_c����!�D��ys��p_
����E�#�!�d�������aO����+k�f�����02�|���i����CN�rty�����Q��� �5 �kc\8@���q6v�p&�O�P;�bA#����	�{�:��%rE����<׶��I�\�(���EȀ>�t�y�ú"QHIJR��()j����\h<� ��2��b�\�ԉ��#�J�'�p���<5	}������I�D<HԳ�AI�V,!�$�4�<T��N݊=P��Hw��4�x#IB6\�̅�S��<E��'�:f�9&�"�h+;Pa!�'ʄ r��`T����]Fur<i�'ٔ�P�EN*H���Ht�'�����,ݿJ+F S���)����O�QR!"آ����I��*X�eQ�L۝p[��j�(��be�,fH�a�.4�Dr/�2r��ڲ��1�|���O1?��%їb��2�G��M$�M@N���D���.81�>��@�7e4��S����>��熹f�ܕ g�]?Aj���7�B�kM�ih�eлh��+Ԇ
�t ̓��<i�К���y��K�\Z̼8��T�*���fhL�(O�|�^_ƨ�i�(���D�c0>���g��	�
����O��Ť�Y�Dx Fh�$6c���=�OIʱ�^�#^��[vDX[�JepPP��]	��\�fA������Oq�X��uj��&��rIô ٸ�Rצ� |޼�m^:,�>X#�͛i�	z��~���l�c��\D�9F�0']�����L0D)R̀�$��gSvS�ψOX	��IB-Me�$*`K��`�p�i�0]��I�G�hE{�ŉ�Lk�h�a
	�HRjM!�N �%��x0M�7�vLc�EV���F�cA10�� �Q֟D�D�n�,A���"T��`�R�2��U@E���Ձ�tq��Ʌ�F���O��MI��А-l�[���,u���}�#rL�)�G��Z�OW�=j�D�Y��� �C5k�JPk@��UC�8�%��t�W��G!�5D��0O�l�gݑ.z��E�{�@�eaM${I�5��/}Bk"�g}rD�u��a�JM�q#p��CF
B�!PG�[���Hz���".2p������O�YB7��.&��� �ݛ?*��2r�iꬌ������Gzb��=-��j��Z&rZƨ�O.}��%�u�
\�*��u�d����W���)Q`Ț�Ʉ�yj��(X�QB�0'*�4�fBA9��'�J8 w���]��c�	%dI^�q$�?A�R����҇�ǆ^�x� v�:��?=���v��B#�>���/>��%����]Zhk��6ݪӯ\�	�*��%���T#��}z�'>A�N�5-�4!΄}�rq`S�"�,T�J>y���O��b���J2Hi� ��
x����b�	-�|��Dc�4
���蟜-����Ƀ}ɠ����)C����*��.P�I�\�"T��-.�pҒ T�xò!K6���p�R���F�)��0g4֡��AW*D��'5ҩ����i� �F�J/&:(��_8'j�����d�:z\9v�ӗ
VBl0?��S"0D�j7�
#Y,٫p��]��	�PSݚ0i^�:�az#�8eb���/�M�ha �	31P���F*=�� �)Pn2�����VQj>�c�E�9�)�`�����C^�{�~���OM�Vn��:�ؔQ��Ce��@Gj�����M�G�0Px�,��v�e��.ԃ8��ʓy֝λP�\���,�O�T�r�,�.�i��	�5^ ��TJ�*w�е�Bʋ=2F,i�� ^� ���
-����#d�剸u/`���)F}�F�=f�}�`�ƀs���E|2�H NԮpz��{ܧi�4��u��:˒rsϗ�S�$�ZrԄ3@��#1�r=(ϓj�j(;4(՚��<:�/<�b��'����Ǒq�S�T̟!},�������g�j4�#�_�0�ԁ�CF���2O$���ѽw6�8�D�t�B� B�ɨBx`����d�����F\�fɒ�C۟'s4{��XD�<�u��U���S��q����b!9Ye��h� �,?P�/O?牧%2J<� b�+e��ڰ-�6YlHB�I	�X�e7G4�@[7`,y���2/��-���ڻ �az�	?|)b�"�>M����Wڱ��>I1b�X;�'C8t�\���ȩ
p��ߑu�!�W���%��Υ	�d�U�T�K�!�d�&E�����Q�v��1ʊ.g!�A'=tv�veZ�|�zH;�j�([!�d˔K~�I
��/��pr���%]!�$2����N��Y1%�*SK!�D�.T�����]�w�|��b�ȵ/N!�d�!C���u��$�*�c�	K.!�䑞n*N�P���#;�8��G
5!�d�Fa�d�ʓ�$�:-�f��9�!��I*�����>����d�ެ$�!�d#_�D��,��^�R��$�H�!�Ė�#I�L�!ʁ���
[_(lq��S�? �ԓA͒5z>)��jήG^u��"O�}�#V}�M(�g�9�,�t"ORLZC�;��z�96�2�	�"O(��Ԭ
62�`���I<M����0"O�A3��7Dߤ\1E�@�d��驧"O0��GϻJ�p#pK�>L��y{2"O>�:�N�*�b���Pa�D�Ab"On���2F"�4ʂl{�j�"O�RS'�W�ұǣN�b�.�H�"O.�7 ^y���t@�H�4��4"O������ V|r�e�(c�ģ�"O6\�E�D�s5�=21.���Ȫ'"OY�L�2x�Ɓ����%���Qq"O"	�c֊w�pH��R*x����"O�(*���[~�#�l�5y�Q�R"Oi��JҹG�Y�rjԢ[c�5�b"O�4I��6s4F�xG6lx��&"O�	�Č�tF�je�]g$���>	%*C8'�t����&��m�p.�C�G4�1Ǝ�"�P�p`
E�i� ��ȓl�88���ϊ]��Y`�U�p� Ą�D>�vn���L8��-�tgP��k��tC����g�1��*�A�ȓ�bp���A�Z}&�ǈ�;zS(q��^��(�R��"�i�)�V�4\��NDH�ӮNwHfG<L�&X��_��-9E�˸N���� ֻ2X�����:�	�Tnf��ISD�::N����r\��a��fĨ��F:V��a��>��c&�Ĵf��h�s�U�>�>4��h(p�[� R.H0�p��\�)��ȓ9�>1a	
�tdwB6���� ��QwD��T+���uh°^��t��7T���B��Q`�ks�5�j؅ȓM����K�<8�s�(O�U`E�ȓ[�X�Ƕ��l@��~Ȟ\��'\��wm�<��ۖHI����'%���/_�r��DSV��xI^]Y�'��	S&�Ͳx�B}��.�wK�	J�'�f�Q�N�O�Z�0Յ ��=��'@Ԕ�!,Ɨ<M��Jg����	�'wZ���i� /+��A��)rj���'#2�L\ �1���
	5���'p��d��,~�*�鈈t\ֱS�'`���U,�4����3��(p���P�'�~QSQ�dX:$ϙk�@�`K�a�<�Q�B�/�JhÃ@�{����CBc�<�Pd�-�PL�s�l�"�b�IU�<Y��ޗ��a��G�+��\z''T�<��̈́�"B�q�@��wp�!��Q�<�b�
H��� �������%g�<ɴ'H(!�p���N�;W�,H�a`�<1e�ٿR���P���Tp�@S a�`�<���k.�8['B	#@�F���`�c�<Qr/ĳyT^�s�J���<3�cGc�<9�O:��3woJ�f�����{�<a򡂒��ɔ�ıH���_�<1���T�$�� հj1���B�<Y�W�c�R]*�M�+b�^�4ƑA�<� F��#8JTi6�^�9�T� P^@�<a��Oar��ꐌ^-zrkUW�<�B V�Js)�f��v�vu�E��Q�<0�ˣ@��iD��^=�F�H�<��厀E����5��)Ɉ��H�D�<��H�WlF%�U�Մ"��%�pO�w�<� d���)�L�Q	G�Ns,�c%"OXA��'D����5�8+Vp���"O�%����?���j�T.^N���"O�A˰@��8�Na�AiԩJ���g"O��c�)o�R�wAE�Cz��U"OZ�oIJ�Ɇ;-�I:3aS��y����<٘��D�N�:a,!����yR�>9��F��.�X�sO=�yB�"%x����Ѽ$�j�8Cc�$�����}A���>E��Ì�W���%@P� 8�3�䁽�yR]fXD��I�G&�cI¼��'.-��I�~8�h���+@��,�p�%�����#�H���EjH�рG�9~єHI˥
L4�
O|mr��L你��T��#��'�p� ���*BX�!^�<��-ꇪ�	��]�ȓW����@��Z��\#fπI^ʱ�O�5��̟C�S��z;�0 恭)���S�r��1�ȓ-0���9B�p�
ɉ_}T��ȓS�F��安! ̪�c#�Ӂ`��a�ȓQw�1����T����El׃U2��ȓ^<��A�ً2fRI��46����ȓe0��S#e۲A���)�M�1f�̈́� ���"X�pԹ�$m�(b�,Їȓi{P�RS�͜��`D-J� Zɇ�^2���J��HS�ۜ�ȇ�= ���G�sn�y�2D�E,<Dzb�>PfQ?	��.}���&C'x�|ȩ��2D��1&� X+~���KS.Tղ��#� ����	T�(��Op�AIB��E���V*VB剔",�&JY,k���"T�'4L��J"a[��O��p��)��|*��L�S�≑���.*tl���Fx�����n�tm��ަ��E`eg��!놃�f^P����'FX�2��	�.�(k��X�}` m�|��{r��$S���r6k
X� �G,���&T��A
L�2�q�`�Nf�ԟ��	�^PB���.$�ic��@�`��T�PW -�F��v�H��d��B<@c�� ՠhx1�V'S ����&�#tv�	 U�Ont0j8扄~U�O��9�k��y	fe�:
�$��'
蝃s�M�BD�Yڂ���R0GF:x��)�ʟ���핡TƐ�6��q���H.LVUi�aZ��X����'90PZQ���)n�a��Z� ��H��71-v�`�Ȓ!=s�)뤫�\�}��(頣ɼt�p�j�+
,�<A��W?��E�!�[3h���E��x�D��&P������1(�������O��97�����0��	6c�]0�&��3s�9a)SZ�a1��'(
P����Nn�j�Ɉ2b�bxz��
�����f�{�`�0Eo��2��:6���`	�Px2H���R@�*�y��XÇE�o2`���	�|GR��Ǫ�Y0P�B�
�;IJ��a�C�+9m�% ��� �"���/9/�ӓ�+,��F��d[��r��HU� �"o�Xr~��{�ly?������:�2�7��C���A&mB�v���X�a�ħO��w��`C6��c`��zH�Lj�D�^�6�kU�G�8�~� k�1}�@e�!b�e|5��׀M2azB�EAQ2M���#�p��4�^�-�4ql��:F�'��x��M�F�8���I� &� s
O<@��G6e��M��J�%X��m��jC���<�fᅒ0�ق�ŦX��iâ�R�H+H���]*Q#�}[֫�5��x�C�*7)D���eI�~Vd1��)ª|2��9�a"{vB��G��S]���O�Bw�)R'�Yc�GV~6MA`��צ2nT�0@�P�`!@�j��!�(�F �fU"��PΝ�W� ��?R�G�S�X��Qnɴcg�<�X=V�W�)X��Uf9�OV=�%Β�F�8�s���~t��`ųb,i���3yg���d
��p%��S!��u#`��N15�B�ɵTK���bDN�B/��iu"�?!k�����<]،ɫQ�p-N��#l]�b׾�	*�,,����^�h�I���r���xԡ.�+,��ȁK�.�c4o��(�h�k�������O̙g%�mZ�2A�:�LU�4��=9Ȑ}��E\�	�P��Ȗ0&&�'���" �q�LM�#	�/Q���L>��7:屆GނCC��8��*@Pb̹t�C>+����daX���Ď:��	���րB�E�5�N튤K)��D�1�^�D�`�Lr�7�j�g�]4V���26B³L�ℚO�� �K`�q$��SD�͟'� k����v�Z9Al��	�&��ėRX�( ���34��H]D�" �>i^�0�1gI#\2r��$�)��1�5oY�r���mP�=����3`��|�t���Y[|~tۧ�����ׯ. GJ��Ǔ^�(�(�荕yby��
��%%�x	��*V>�$�!�©r�Y��(�W��O2����Z(.�>�����{�P��#34���HҤ��=#�Ad��$L�T��B�d!C�龟�?���b�]���8��R���p&T��n D���&���PY@��~�c���>��*�"Z�h]�go3u�NY�Ћ\l�'�"p��b$^�ș@רΙHE�;ӓ2dL�iP�\�bԌ��tl�{�!�9Q9"59@��E��ՓE�����+Rs��"EU6�PħU�P0��Z�`'�I����X�hW	r�Tdc@5 �Zҧb��%����+EUR�w�e~�ۿS����ӓ�������F,*`§&�J)��i�a˩Ol�j��<�B��H��:���� �i/���#��?n<L����ћ>x��"O�-�Ou�`��f�52����@��O�i`HK���-�.��Ԁ��>!��Z:�m3c	S&�楳v��9�B���ɜ4V�y9
L�p�
i��3rU!!��#q�(�G+'�(�2��@7V�j�z�@m�D��j����u�$Oj��TI �A�v!��p'���9�O�b��j.L/7h)z�+_;*�b�����5nҀ����/s\QAF���AW� �[<����>� A�תĚF�����F��I�uMR�0G��6�M+�GP��O��B��x�~�S�$F���vHL�4u��A�'%=eL�=
��9@ �)": q�U��O�ء��#$ฑ!��?�< aT?!�<�tN�4m���3��.wPƱI�^x��7��7�ưK�..'4H�������p���	$*`�T�Z���I
�A��&\O��ȐnɿvƤ�aPoH�!J��D�|RgX�Z�J��@j��L)�ha@R+f5U��S�DB͗�	F�֢DO���/���y�MB?27@%��*�:�� P&�ٖY$�!wDzo2p��EBm��t�'@J5�6;�R�[�G� M�����-H9��O��C�H�j�����#jJ��r��D̄�m34��cBA�+:. �چ�� VU"=!��ם���J�k�\ ���	vX��5���MVj�&�3,����gT,P,yX�,X���P�@��g���#͂�M�txp�'�ʸ#B��@����ʑ7Z�(K<w��/���;UnH)��	���0P7�8��=O�1��H.`u�y�d�_�xw0=���G��B�Ox�L�?>�])��6E��T͐�>	ty��ť"�naP�FD�x�D�7;6�}i43��U	5��p b��=E@����2:�T)�"OA饡��u�Pi����,���R�i	�>��X���r`:�$�G%Z�����N��M%Y���3�0���I�.��uYU��_�����I�5u���A9S!61gǚG.�#a&Q�[�*�HT^��,�r��
R�T�A���@����ɍ^�4bSG1I*� �Ɔ%dT➌Y_7���W̓�&�j�! E$#����[��xQ��YkxI#�$���j��de�/q��C�	�gb��Z��A~����FR)��y *��u_���拒)+��"��'���|"��k�Źd�mL	�Aə?���*D�H5�@�Kԉyjľ� �y�*СTS
u�L��`F�H���7l�H��$�3t�V�B��
1eB1!��F]0a{"�\f�>ً�V�'(�TФI�^�)��AL#���CħH5-�u��	�6l�`LQ=E�� ����\m�㟴Җ�]J�=F��a�)�py��91��!xqOP����R�(gة�t�I�� s�·�7H ��	͸Q�H���ih|�kt��I�\�(MBf
�
���3c�F�e��U����rm����'��c��>/�� ����L���dC?F���pf����O^�ab�_4i1�-[֫�z�1��'����wM�Ϛl uWjŴ�0޴\�I��X�	��ҧ����L
)@`DqB��Nb�M(���y�9�T��@�nlp���-����wn��1��Hx�@3##���MѲD�6���a:D��!�aP�nE88�W��<K
LB�#D�Pc0oR�N��؊⊋�5M��g�,D�x�(��$�\ ���<�ءZ��0D���WH��Lh�$#ä �9��I)D�# �͝u�`��A
A)b���鴉)D� �rg��x�,�PI��z���+D���+:r�t�ۍL4l�%�*D�����B�{8���O٣^�uA'(D���%� Fע�`F��1�1IcN0D�� ��h>TL"4y�f�5(i6���"O��cu�[�x�����K�XtP�d"O�<�FN)�9�� B$PhI!�"O�1Q��ҐaU
��`��N��P�"Oj�k��[42��m1��+o'�$[�"O氢�d�3���BvA��!2x0c"OƥS2�!]�f��s!�J���B1"O��x&4K4p<�q�� �89pf"O,IJ`�G�>���A@�e�j`��"ODZv�	�9�*�%�4n��
�"O�<i�Q0:49w���Uc"O�ʂH�!���6F�� �"O�|� J�f�,��̆�,�`�S#"Oֹ��N���P��A�KzL8(@"OQX��ӭ7p}���Lxw���&"O��z1C�jD([C��]@Tk"O���6m�hd�D����01"OܸȦ69d�!�ď�q82�"OD���
a�T����:>�e"O<����-%��@��):�c�"O(�P�m@�B�0;�#$�Vpӑ"O����S0T��hHn��/2r���"O�����˨I���ìN+D!`�zT"O|�jĉ�1��8�kY�r
���"O.�S�%��e?2A �ҟ(��A"OP ���$l�glثej���"O�|A�ǀ�Ts�	cɘ*)i�ٳR"O�T�fH��^�h�@�h�tְ "OP)�(�����J��Z$B`�c"O�5fƺ�4�٣(ޜ"K�PF"O���先K�НhAB�hj�1�"ON�
g�
�G�Α�V@�)xC.\�v"OTY������,%��5Y�6`�"O�<�G�˒$���iRU��"O��#AI���%�q�1i�4؁"O���a���o�s�5���"O�abM�32Y��ژr�p)�4"O���A��<��#'Ë9a<���"OH�FEۯo�$���Oڞf.�y
�"O�	R�*��5cAѐX�=9"O��	A�=��#��7��d�7"O�P�)χ���ҐϜ�FԐ�R"O���3
�gw�8B�B	#��R"Odq8Q" 4uq� �J `�x�xC"OX�ـm)�@�q�8e2���"O����)��V��!��B��Di�"O�l��K߃o4��d�S��P�"O�,p��Z�@9�'�DF�@I�"O&,�w�ޣ_P�]�C�W?��a"O�%�榟�gC���W��B�ܼ��"O�SU�1/d��G�?=t��A`"Od�Hċ��IC%h��9�n��"O*��P&��Q���>q�Ւ�"O�,��ʿ@�Υ�UN�'�8͡�"O dq�f��z͖��tn�4}����#"O����(��]�b�a�-��m0�U0!"O��v�K_WeȀ�d~���"O�|{E ';�$J� w>Dj�"Oda���9L/���� Ʀ6�d�R"O�0�V�3K�*������k�"OR��g�
��t�֮��.�ȭb�"O&|�%�pќ�3d���Z"O*a��F�3���{��Ύ}�X���"O�q�,U{�J�J����"O� �t�$���$�f�7 jIi"O��f�=[2^�+�)^�v�����"OP��gY���ر4�ʊc��qp�"OE#�F�(��#�u��U�"O.y��,�o��@�7q��r"O<Ԩq� }e��1#)W�aR�"O��a�/T,`���[�Fd�#R"OF��,ٞDIm��GY1,FP��"O�@��H=$�2Aňg@\��"O�؃�n��f���# E�w�D5i�"OP�CC玩i�bT��<%b�q�A"Oؕ{5k�D�p�NΌ�P���"Ot��$`A�5u�q���ȪfM�TB"O���*_�:2��㑥Q:��؋�"O���Ҭ�6z�Z�C��|�t)�"OkB�&vaU�D��
]a����"O���&�T��:ڦ��FO� S6"OLH���B��ݐ&@;��g"O�,:e��֐�T�ԍd���� "O���B��Ws:,0	ΓG�����"O��Õ�24`��w,Kƶ��4"O�x)��Ŵ(L�Ա���6����y2��\���D0�� ���$�yҸd8{!`ƯujL��v�F�v��l��&��Q�E �6A��QcW��5x�ԅȓ_s�`zgl�xu�3ݳE�`�ȓ5��Y�7#b0T�B���$p�ȓpDİ
 �KZ�:��_�?��ȓ00Z���Nϕ}�t�a�N�8עA�ȓC������#K����gaB>"��8�ʓS���:�h2�\SG�^2��B�	�@�t��7��R�,���\o�B�	>R&>H�0�σ 6 Y֭PX�B��M�$\�Fŗ>C�aSw�P`��C�$:8�a�T�l�̣��ói�B�ɇq`�� �J�4h�n�  C�I�h�����1-�A�G�=c%^C�� �)���Ա��9��:m C�f�,�Ņǡg��a"�
	��B�9/l��G�'TW���ՑfH�B䉗m��	��G1�p�Xw,\��B�	P��ū�n�GI��� �.�\B�	!B7L�q��3+)N�Rd�NZRHB䉖N��&Gq�;�C
�&7�C�I�!K�X�-�m�|��$D��!�ʥm�: Õ&�w�h��XGh!�D֊6��a!*DKުe ���3T�!�DH>f��k�.���W �Yp!�d^h�Ny��n���K���nw!�Ȩ�aj@2��N\;<Y!�$�4/C~�Cg�X�+VA�-��GV!�
�s�R�Yw���K�(5Ӄ�lM!򤍃B��ͺ�OW����(�f̽"C!�d�:����
��lDa֜B!��7Az��*�~p�́���65!����U��N�Fa�0{��<!!�u�\�N��O� �(@朌^�!�d�N4�1aQ�	%Q��L�� %�!�M�r�<A" 
l�>
SN��p�!�DY�|U>�xVEԹv���CK^�m�!��_>m��q�֌З��t8�	!H9!��7�)��a�	V$��bUO҅@�!�� h� �V�\�D$d\�3a�3!򄖤X�x�'�
����ñ>���S�? z�P$�^0�]��n�uT5�"OR�K�/�%�jyr��Z�wȴ"O�E��I+������<j}���"O:��f(I�4�IA��~o-�f"Oz�(!F�v��0P >SaH�A"O&""O�?�����T�H\�@�"O��1�%ӏS����#�ϱB͊Ui`"O�X��*äP8�q1�4}�����"Oh� �J&b�~xAЫ)�H�I�"Oĕ���s&�ȑȒ���p4"O4�+`���a�gȁ
o��*0"Odi���+~�feh��˝]��I��"Oҵ{e�^�7��T�s�	{}�Y��"O��J��M�l%*q��kY}��k"O����8�Nh�
P	.��
�''>��u/]BD`'���ɖ�y-�#ER�Ձ`gTn�fmg���y�:s��� fBFE��.
 �y��݉KF�)�l�7`p����)U6�y�.��
5� *qh�'R�rQ�4O��y��Qb�bQC����<]8�t/��y2M
�p'85�Ԯ�.�������yRʛ�S�N����'b��1�!��yB��6]��!�1
qb_��ybSU����(T��m�#c��y�Dʳ	�\`�e��~I���[��y��.]LpY�R˗��`�AR�@��y�&��"�r���e/=��sQ$��yrEX�]�x���U�)j
��Ս��y� D�]�0đ ̀U�ে��y�M�=P�x�E��M/�a�g,T��y��B ��	�M�,C�~%�ׂ���y�K��i�� B��t@�MP�y�(K�&}[�C��=v�
f+)�Px��i�ɛe�Ċ*m�R��ʭo���'����`��}G2X�*�!l0�Z�'��B,B�\�H�0N_&mL��'�(A����-fn���A��^�h<��'�Pb���i�콓�	ʛ_�DhY�''��KFC�rxX��B��W86��	�'S�ċ�
�\��Q�W*V�~4a�'�Z���""r�|8a��Y���'�t̓���?W
��	T!M�X|�P	�'���K�֛op QӬ�6\.\�a�'�0yxd�NL�X���G$Gݮ��'^�\�&.I+�� ُ<{0=!�'P�l+0��%���;#K��D�TY�'h�+GBRg��b+Kقh��' �a��E!�z���n�:=�d���'�|l����|ɦ��!^5�*p�
�'�^�u�Ǎ{��*W��-���
�'#|P`�R2��iҥ�U���'D$�S��5<�Ȑ��ƹKA�I3�'r����K�oCh�$n�qq�Q
�'#\�AH�wp��⑸b��T 
�'�p�a��Q!~�0I���ڣis�	�'�l�{)�:�`@�r� �82>�P�'k��)u��7�:T`NO30�`�i�'2�X�#%�D�h�A"[���'K
 ���J�EX�� ��#Y��'1F2��� v��� �-��l*��
�'��|�%�Zk��S��h���'��T��o�9Ǭӥ^P���'�t��Aݰ>`TA��B�`���
��� �Ģ�B�x��u�PE�	8+�"O"h�dP*�2%ܫ����p"OZ� �)�A7x�@׉�R���b"O�{U(<-P��F�6�L��"OF�)U�J�v��}�c��Mɒm�s"O�m(ң\�3Ғ ���2��"ONEH7!�	D�f���B��M���S"OF�ɦF�}.��xr�ݮ�F�"O���4c[&��4��?Qy�"Ox}`e �1�.�����+N�Q�p"O�)!���)
@�A�Ȳn���1�"O�XRҠ)H��E�"�������"O�<�M�|�8(�VJ�sɀ�i�"O$��Aҷ0�� ���=N����"O�����z#�M8��=)^�2"O
 ��d�h�v`C����+�n�<a`��&g�ۥŏ"uP��H%K�q�<a�3^�(�sTX�L���h�<��^&HW6� �BQ�qW���|�<��ߞD�$��#�8��2nI|�<�a�۟y;�5�֧�3"lͳ��N�<	ulE=��x!èqhb�bCb�<!���4��qF$CX��	��]�<)�,�Wg�z�����"d�s�V�<�ǘO20yb�'
:��\��nR�<��/ٱ3�`9��e�(|,Q8��BO�<Y��;�ri� ����8]���[M�<�%�Qb��6j�*���P�[M�<ab��2[<� `@�-$x��E�O�<��m7�R,�*�0}C����B�<��P�%��k��֯Db�a�!�w�<A͟3�}���F�d#x�Q�%v�<�.f�`��̖��:���Lt�<�&Kn����y5�,A �Ls�<9E��<�J��gH_
��H!%Kn�<�7dX.�R`b�
�!�r]rW�D�<��NH53?���/̸1��T���S}�<�3B�Rڈ���7{�.lzD�OU�<ir`�%�������
�.�C�B䉵@o
��ƃ��H���c�0�B�5X��pc��5�{4�FVk�B�ɗ5��7�C�`�Ҥ ���PB�	%Ͳ$��̔�`y�#%��B�B�ɪt�� j���4���@�@K�H5�C�	f#�}HBG�#��c�`��pB��S��E�iݜ/�f�B���E0�C�I"kJ�剑�ޙw�@ �vNK.�C�I0j�L���� [_p�s����B�I z0i���YZ�X�ԏE�p�B�I)UH�@��_��(1�>W�C䉜L\0b�էr���5�EK{�B�5CvN}��
�fa�M�e��<S�B䉂V$t�QG�^�p^^����1K~B�5%y�|�/�2@J��;|�j"O�#&"��k���*G���<�"OX�gZ,i>A[Ј��"���"O�$B�c���Y�IB7O��H�"On-�	J�n򌙨��Ԑ|����"O�m��*B%O����aGIa�DP:u"O,(R�H�	A�ytE'u�"�hg"OAe� ]�V�.(郗(5!�$L(������h
���炎G�!��Ϫ?윅pt��1�`���M�'e!��J��D�`�߯t�]B���@�!�� �9 U"!<�i���x��D�r"Ol�@A���y���!m�)?���S"O��S���#�Dk3�؀���`�"O������Y��;��ɩb�.���'�r�� ��!˄"e/� B�N�2�'r~u�S��v�@�%��$Ko��'�2̈ק��A��,���_�z H��'w��4@�'�~�j+=s�4ya	�'��1
PǟHM<q ˽�~��	�'7h�&�� �f!2C�\�AӤ�*	�'��\�#FN�zt;��C�@fF��'`��($��\ :a���'���':���h�2fX:���m�: $nE��'7���ɐ�Var���+�7fb�"�'��9GcL��`y0��H"`%��'2��jdN�l��
7c�7�'��#�L�(A�s%e �h��-ҏyb�)�S
#��Ap���x�()��O��	�C�	?Zhp���?R� 9�	G�"rB�ɣ;�Z�3S'�C���%K{,:B䉩.κ}{�T�p��g��z`B�I=���Y�!�#A�A0)�(B�ɱ6��N�&=6��S�_�B�Iv���Ӄ��m�ri��J�0SB�ɛ#r��+P{�03��G)l *B�	m:J,;V�\�D�(a�g�6$B�ɬmKD�I�E�[+a0�d�>\�B�	%,�x�@��nZ��1G�ANB�]��T�vk�or*��=V��B䉊j�<K�
Y�)�*�jW����B䉗P84�!$��+y{���C���B��#	2j4o��b ��l�2?�`B�I1!���S��
u��Q��=�C�ɋepd�BR��[�4A��
�.8tC�	�HV���Me�\M� V�(�RC�6�	�A�<{�4�q���8"�PC�I�FLNI�d�ԵW'}�Sc:Fx8C�I�0�j`�4)�#�0�a�C�B�	01UpQ�6n�A-�xط�+^J�B�I%c�`��	=Bl�Q���\�=#�B䉟4��xs�J�?�Țt��A�JB��K����G p�k�ȇ$L4B䉄/�FyH$e��A{�l��ᆋVGB䉤E/v�:g�B���0uj>��C��%s� 1����	6�:���­T��C�I&�n�z�i˩[�mZ�'�45�C�Inm2�Q9)9�D�Q�>��C�Ʌz9��J2Ɉ:�q����Z��B䉦J���зrj�V�"r��B�I!�>|�*�v6-���aq�B�	�o�n1J璠�8a��J[�L��B��-,
�W�5R�&��a���9�lC�I�&��� u-�d:��;���-{@C�IW�=�1hw%�u��C��FB�	�X}3 L�e���V��(�C�I�~�6�PRL�97�a��Q�h�fB�I�x��\��P�{�Ac�P�MAHB�	>cy�Ơ��DGh�9T�N%YC8B�I��rH	0DM8%��%��C�ɋ!^�t��N�Z�0}�r���C�C�1B�Q��I4;�U�Wϓ;��B�x�����Ve��=P0��RMآ>ш�)J�[L
hI3�@D���A֦G,N!�I�)Ӑ@Ig���L{Wo�7IR�)�� ά��O�0���b"��=��"O��*�'�
*m��%a��l��@"Ox�P`�E+3?d��o��=�0,�"O��j��PXLC!HT�}HA��"O|91%�W�\ z��ҧ��$�\�A%"O���q���R� �Ɋ"�~�r"O�M�G.�:(��v��9��(��"O8�y�m��A�i{d�H.��X�"O��
��Ѧ����#�� ��=��"O�|±Nǩd`��P��"Ԡ܊4"O�%	�KHL�y�!��44x�b�"O|S �Y�(�ܬ$L�k���"OV���$y68���:���	�"O���Sg =~J7��{�8�ɂ"O���F.>'�0�Vb�<%���t"Oy0��J:&9lhk�gˆ� "O>9����E��W ְP�sS"OPe��]%i���;�Y�p��3"OĒ���TLT&Nޔ���� "Oh�;$��;E�b&mB���K1"O��CSZ�-0]�7�[iy2��`"O�qr�a��4'4����A�_X@�9�"OV��GO��y���s�ܕ$!�Lxc"O,"�&��T4,��iS�P=e�"OЀ��K�E�0�{t5$-l�A�"O.�j��B�_?�z�.c��Ŋ�"OJš�ɂ?3<�Ѱ�=J�P"O8`�G���Z�√�`Ww;~e�u"O�蠡�Ė_ p�p�	b� s�"Oȥ�@�U,��!��n�:@"Op�ç/�&A��i�Pn$]p�Ԃ5"O�8[�H^(y��틘0�ڙ�5"O���T叼=��)�I߮@���p"O�IA"	I���1qg]�C�dT[�"ON�#���T�0!(U�m�4R�"O�]�#V�Y��q'Ǆ�_���;�"O���%�*[���KJ<8ל��"O2�w�D�1�>���͚�a�h���"Oµ�k�<0�"f�K�]{X��D{��i��)����2 E]��1F��)!�A�RtH	�anܵ ۾I���Y=w��F�)��18��E�)ܘP(�*�l�2�!��q�8G{�O�O:�����(�l,qCk�I y��"O� �J*&88���ވ~ܲUc�"O�m1H��Z���!��nD�"Od�rL
�7C�LC�D&5c^�9e"O2Ax2`��D�u ӳ]�|:�"Ot�I �F;`�zf@�`DZ�a!"O��Q��J6Ħ	��̛'4��"Od�����XK1�EEفs�Ie"O|���V�����	�}u�y�"Of��aiژ���`�/$X�"O6�+7�֨<0�\��I�U)|�"O�yQq��V$#E�РVfq�#"OP��b��=W�tq�r�Ћ'P��"O�ɵˊ�[�fyrS��#4�ы "O��(��S�����W�B�r"O\��h��ӊ�%F	z���"O��#=E�d(�㖬?�D�"O��S�ɀ�p�x$bW"Y�T�R�2"O��F^>/^@����%YS��:�"O�@�T�U5ƌ@T��*F�4�7"O�HZ��w%�"BL $	�P@�"Oވ)�ělV�����ß\��q��"O� �a J�!1����M�9��Ċs"O�@	2���_R�5�2JS����"O��aF�۸{Y2좠H��l�9Kr"O&�I�S�;��J	|�*0"Oވ�#�Ԟn�����24U�Y�"O��ʥKL͚��� ?N�ٕ"O�T��
�a�mY�,5��i�"O����_1@ �2'�A)��bB"OV�څ��'(4[w,D�y �$��"OF�����;ZАk!��#rn��"O8�$`R	F�aqW��6� ��R"ONeٲiN�Q ����rf���"O5R%#^�lH�y�@�3
��	�"Or�k3� ��1a�R�Y�ʔ�u"O � �2������C�<
�u�"O����M�/��Pv挢�q�5"O��1�A��:����.I�P���"OH!B�D-Z�����-��G�~y�V"O���wkS0]?T 0 #����"O��`�F=f�r��[3BWp�"�"O����:5���֮E�}��"O��j�M1Uz3�d�U6�pw"OX�ʀKD�3����A���t��u8"O$� U��B� ���ʙ=tKF�s�"O�)k`��2tBfjL#B�6	��"O<�V+ټ@������C�j	�'�D�U�Z��EȒl[�h|�
�'��� S�W�(���
X�! \<s�'�<�AwK�$D���4`�h�hy�
�'��m�"NV ��d� �h�����'�\�A7n '�tX�hW�f��I�'$�H5F�//h\=H�bԶ1����	�'���'!�s�$@eBĔ����	�'�Y��� )b�x��]f`B	�'�(�{�� ���6���`y�0[�'�ɋf��"R�9ń�*٤  �'J�݈ף �4L0�&R��`�'�lp��͖�L���r7F���>�"�'����v�LU3��8(���<y1
�'	�Ij�i+ �(X�M��B5	�'��Nt�<Ir�;6��Gk؎�y���6w��­�(�rQ(D�]<�y�A����1�ƾpnI�sϞ�yRhQ�>�v�Ss�A܆l�S�\��y��y���gmMR6��dEH#�y��Ќ/%�5Z7��<j�it�֭�y��
Qk��� �v��c��/�y���Y�j$9�`Pv+b��/é�y�h�5�`IA�.+{q 18î�yBDХBn�	$�M�A���sc���y"c-a����v�);&�ȱn��y�[^8@b�����Q�QbM�yR��oR`�{r˸DR���@��yb��i�Հ��BN�zA�G6�y�DɊVc@dk���),Q1�-���yR�۽r���X���6� �� C�0�y�D�6n�Zp pf��ඣU�y�B� \6x��������а�yr��J��i�mDv��E���yb�'_Bx���^���t�t�%�y�v�:����{+�Bt��"�y"&�Y
2��G���}�n�kӥ���y�� 4��!��D�G��x�����y���S=BY(�%ۘ*�2aɱ�ˇ�y
� <m�B�B9L�*3*�7t'V�!`"O�1�KI�6������C9;���E"O��$1��i����
$�y��"Od��[�E�>HP�R+��� "O�]Z6�S�d1М� �\�V,��"O� [��ϖ	h��OM�A�Ji�"O3��B�F��խP�D{��H*O���7@%$�)"f$�*5G�lC�'�9p��1��逥E���HP�'8 1Cŋ�+4���hՀ�ha@�'�����t�:����ݥ	���q�'���Bh˝G�����<l�a�	�'�MZt��")�`����k�] 
�'L�\+���a?*����Ǚs%��0
�'#�=�D)�$k��p��	��f�Q�	�'s���,ºM�>�a��;XC,M��'�\��7-�6��B*c=r�+�'L������r�z�hI(`��(��'Ȗ��0��)�H3j߭QF��'�*(�-��[�T�A�Hƀt��'���q���&Z�KrjR�v�*@`�')�8��.ީDO�H���>z�ɋ	�'4��9�ڗ	eT�AR�f����'��������/�����V$0��@�'8:�'cշJ�3���w�8��'s�$��]�MZ���u���!�'������U8	 �ˏ<-&�H�'��aU/���	�T�O-3ꨵ�'<\�ZC��� �ǈ�<1>���'�x= ��� GL.��U3#��
�'���ysAO�?���!!$��	�'�x4�S�T�K�ޥ!SK����	�'�L5x��֢oIfT�+W��]��'�`M0%���d�.P�.�(O��i��M��c���.͡,H��f� D�<
dj�5�JT#�h�_���(D�x��́��pM�ƈ�h���ۡh&D��K/�DDv��gK�#u��T#D��9�
A�o.YS���+i�����?D���R%�d_�Q�ǌ�r;"IA�<D��HM�J���yQ�	�x���.D�|�'.E�[F|ɢ�G�uy�P�$/D�\���HH^�ѐ��
�C��-D��+g�F�l|�K2��;w-��zG)*D�� r��6��#�X*����&+D�@jՁ��)P@H�Dۧ���N*D���Ѓ�Vd:E����iLʽ@(D����皅n�(=��n١de�u2�$'D��8��ii&�ZӍ��k��D@�%D�42P�(GN��[�"D'o���1�#D��C%�f����7�\� �&`k�!D�D���#/x�R��`��2Fi2D��ٱOT-p�>�f)݊R��0��-D���� S�L�$�N����I�a�5D���ǇS�"F����@�r��@�(4D���"�T���,KR�	B������7D��3RF�E����F�
o���g�5D�� dn0t~�T���.|�Q��c8D�l�
��Z��X����p��EBӆ2D�0�s�
>`WD�5C��@c�1D�8c��+U�\)�]R|�q�e;>�!��X||��� I�!V��x�Jп�!�D���8%�9Qz�"a�291!�$l�ha�"��.��<�4l+}!�� �:�#�>gG��!+�(*'"O�0ـbS fXl�!�M��xK"O�T���^� ��s7�E� j4�rw"O����Է@�<
�Oد`��"O��DK�r��И��'0q��D"O��U@��A�,e��5e�vA	�"O�`h`h�2a֖�p��S�s^@I��"O�<����{�hyC���+�f��"O�L3�䁲��M %��t�δC�"O8H ԅ�\�8�����(���c5"O<�cA�:�@4{'`���Р �"O,9��D:C`��2v��d�<ї"O*�	4L�
0�0qPp&M r�:m��"O�ҡF̢�fH��ҹ,Qi5"O,QE�G*\�@�sЃ@�5̰9�2"O�Ic6���yx����UД�D"Oh���Ҟi�>�ःћ59�̪R"O�02��/M�`��d�W�cL����"O$���O�͜	񡪘���6"O�郍H6!�`���Ѯl}=�"O��3�E:>��1�w��}��m��"O:��r���͠C@�'+��RP"O� �qx,{#�|5	J%"O��Вh�5p:��`�ؔ9 �f7O�&�)�'P�8q���Ϊ$o�i�8@x�ȓ<6��E燉	�mb����:�!��`|T��$�I'D۰�3���Js�5��i�:���KۂZ}T�e�cWX�ȓn".�+�+źH�콲ҡć{X�ȓ�b�q$�\*��Y����5h����i�T��2C37��)"T���h�Ņ�X����V�	T��!W�T�S,�9�'}ў"|j0��;3	�4�]�e16|����d�<�t��&`�t\c��M�5���(�*Nb�<���,?e���ab͟J��E`�V[�<	�^�H�0e'▙}ؤU�S�Z�<�S	�?zЕs� �<X2rC�^�<Y�U�c�0��L-�y�dHb�<��f.)^]��hV)^���p�G~r�)�(O�,�%��J�͑Ta�]�a؂>O��=E�4��"z��ّsj߲�J!녦��yR ��b��t��D�^N��d���y�&��vB@��,)�p�j���y���BBq:�ɔI�~ B�2�y�
�5K�����+�z����]��y�	W�YHy��)��+Q ):`�+�y��'��O1�6ʓC%�u&�?G�0 � ��?m���M>-O1�1OR�n�.%�)�ր؎�S"OtS��])^��U�B��4���b�"O�hх"��m��NQ��.}# "O	HA	͢j.�@0�LK�8ܜ)҇"O84���V�0%�9�KƝ-�$<��"O�9B�b��ZQj9�������d4�Şs���@���V�#�З ޤGx��'5d�;�H�8�Z�{�͆55��a�'���)�O� 1�	CH=P�T�
�'� ���E1��K����;xH��']� ѩ��3��0(�F?/_:�K�O���hO�V��@e@��(G���nʴ7�B�	�g����q��u3�����j�2B䉓U�s�yi,�h�fֲ�\C�1s��mkآb��  �'c<C䉵mxlڀU��\�&Oͬu
�B�	�'x)Z��T@�1�K�~f�B�)� �Y����H��X���5W��`""O�ʰ��'.��$1���6炰��"O�P"5$��H -�RC�&��a"O�m�FH�P��$�T�J�5�.U���'�ўDPdDB�z�  +��ڼ^�b��5�>D��fL�4p@�zw�Y�(�~�9�*7D����v_�uH!XN�B!�5D��y��(]�VJ$eN�c��g��E{��	Tv�uy�Ɏ _*�s+،+!�N%)h@���Q�HCp(���h�TE���Gu�T`��*G���QlE5�0<�����'T�p9Ӎ�+P���A������'n���IM,k#����F��lT+�'����5w��!���R ��r�'�LU)Pf�� �S��]�p�q�'�b0�4�W�8��cW�P���R�'m�U�Q��(|ך,k�E7H���Ȋ��8�S��3vA�=��.�,����df���0=)���F�].����"+��-P��y���.~a�!� �Od�ԩd�C�y�F�|r���c��K�Bu�3����y��Ӳrh6"åAa����^��yB�V�U��	q���7!�\�E��+�y�$?t����+���P���?ʘ'�"�󉒬6����DA -a20C"*Ш�!���h<e�%@V;cf���Ǌ?j�!�����͛��\,7�����i�3�!��:
	B�"BN@�ҙ��ވ*�!��X�̬k���I�Q�Ս�!��	
�0�` ��"B��h�P�]8e�!��ܺ`�H���v>D�w��R!��#"̨ @(�p���͓Sb!��bx��➁3�4-��AJC�B㉏k4�Q�O�D|2�%�*A
C�I1&��LI�'3@ �G&S�c �B��'$���'ż{�Ђ�	SS��">ɍ�	�%��Ջ��H�z�q�H˞3��D��D��D��7�X�+�d����y�H �K���r�+O�2�6�11"��y� �!j���r �Y<(K��/V>�y�*X���z�`�&Uj��Eć��yb�� Q$���I�>?>�0���y"FA�	�8qs�ɘ+���4���O�ʓ�h�Z��ӬK�Ks0e����<U���� �'H�����@�S(?�N��F�۵>�!��RX�d���Z��?N�!�d>`�1�B��cV����5Z�!�d��=�n`ɶ�f$�QQ.N-4g!�$�$-ၰ!�'_��8����mN!��#J�,)��KâP����*S6!�E53�����X�ȁ
v�Ʉ�!��I�Nv����,o�MI�Í�\��=E��'��h����U�B��'���)�'>)�ƺxD�ء�F*~�'�V�8b&C�Q-�i� (�Tu��0�'Oؼ��5|�`��KI�}0�'��d�d�N0O���ՂH��pr�'i>�9FdJ��20Q�I�@�`��'
�	Y���uLdEP�`	�>�fy�'}�h�х��]y�t9�E�5j��ɏyB�'��:tC�0&\!谅W�����'��ݘ�c�Q"�Cк g$,��'��}`��IT="@S"5��
�'t���D<|S|�p�]���	�
��� B�S���~���d�K.@����5�Ş	b� �t�ʯ�R��je��Dx2�'������U!=�	�`�����'j�3�D^%I������i�D��'hRE)���'��+��ZG���'�N��c��9�h��� ˳Z�y��'.BU��!j `Ђ��S� ��
�'�h�fg�1>�E��N�� G����O�=E����,��eAF��\��pQhҳ�y���1h�
@G��WT�(�gؑ�y2��?t&	��GL�ڈ�T)ˏ�y�mȱZ�"���K\�@a����cߧ�y��')���r�#4� ��eeד�y�0&�4b�bΠ,����dN�yҫW3bs�\0��C�#�̅{ե�ybDJ�E�\@K&��bJتC.�y��X�(}^�����TF�뚄�y��4�١�
i栀��������<I�0T�1xס� j�R��A'�
�d���I�V0Z�O�*(%F`x��J/Zx�ȓ{����4g��K � FY'tVDt��f#��e�V���TG�q��t�ȓCf=�@F7�=�-"���P!�D@�<ƴI������}�o�1T!�d̉+V̊��A��*|P4.D�KS�d�<	�)8|X) +��+�>�PW透'6��ȓrx�Y"#�� A�\!�h��rJ���h��D�#�� Di�m ���IB�����I��Q
K�D3n�q��(�ȓk:��Y�:�{5g0*��ȓ3�n��nµA}��D�ܖR@�����l�2uJ�A0���
�%i8��yh��)�T����]�&���*b��H�E�[�|Qqc�m��ćȓh���x�&��1�P�bAJ*��a���?����2�P�"���u	������X�<�7�T�d��I�*��8P�X�<YvJ
 zt�F��B!(�,W�<��	x|zXC%�AY���#]Z�<��
Ԗ��Du�,���+��a�<��]�&����w�&qb$R5EY�<�p&��d9(���&�i�h��<Y���?ɉ��I�.�>��`B�O�Z�S�%?�!�ߛ4?�p�q&�9���DJ6R�!�H
40�T15�I�-�,�*��h�II���������\ ��h)a�(�9�"Ohe3V�\=���g&ƻVtTi�"On���@�r~<$x�e� s���O���ϾV|�}��X�7��)`����1O�=�|"�'ss� ����4 �`�2��j�<1UMp�tS�4#� i�*�e�<)!bʮ&�v�8W�Є��P�Q�U��hO?�ɿ1���焏���ub�,��q��B�I�o�����7��!ԩ-;��B�	�4V�Ⱥ�*"
�T�qD�^1-�HC䉭�~�6	ʉydZ�qG@?{�B��+�*=a��<��hSٜ6JB䉫6�}�/Ʊf��`��8p��B�	�#�`���'�iX��
ת�������<��*�?uܲl�K[�}�x�"O��bB�ݸ7q��i`DY�(��y1�"O�4��`A��Zp�QI�3]ؐ�#"O�y��F�@�p7H]!>Y&`��"O����t�\ dGP�x�h���"O� ���V��+]�ٙ�e]:6�ޠ�u"O�a%��de�����2y��"O�h��m�eh�IB�Jh~�q;�"Oh���x��UY���0�ő�"O�a��������"��|ȸ��"O@����6hܚE�����_���H&"O�h�� 9��Xw���k]���a"ON�kU��0�ʤ����uv� �"Oj��]D�L:5-�g����"O:� ��d�V��p�]�M��5K�"O����\>U#
-cfjIm�����"O^�9��K�9P��q�Kx��5��"Oh��g����l C��h%�qQq"OnJ���f^�]	��
��(�"OH1��唆f��Ɇ�ʬ'.pp�"O0�m&o��x ���"��0��"O"�YV�ǫJ_b$��Ν	s�v���"O���K��d��60z.��"O���
��V� !,�1qP�{�"Oνr�G�2���QL�quHk "O�q���N���Ią�XD�"O-���\=(��rvN�85�	�b"O����I�Zl������ )NE�"O�@��ޜ/��a%O7�)�"O����e�ך5y�c�9$�""O&��QcK��P�C�K
"��f"O��j��XO�pI'��d�T9�f"O���tf�(X:h�@�-c؊Xp�"O ���ܲH@ %Z�y����"O��@�A�Oy۶��T8�YYf�H�O"��
]!�����%�r���'�:�eH����+7���Ĵ	�'*�dc�Xz�b�e*���'׊��ҧ���m��m�̀�'	��
��j��=�"@�.��5�']����%)�!ʱE�/�H��'�pE�`]:~����
$x&�mY���-�S���٠5�@,+�L�E��xgaU��ygC�9��Pfɢ@��D�-#�y�6x�����I�}��]��yc¬|����1KE/<#��J��κ�yr���G<|�#�Y!2��Y�G��y��P[J�a��;#���U��#�y2oʀ�LcF�+��$�5�Ov���+�����X1 W�I�$ �X�<�VjX�7$h��2J�;&�tY��(�z�<�áG35���˧Kƴs��I+Sk�<�/�u��dQ��JB��TB�l�<D'��2f؅ �	j��@�i�S�<��$@0�A�*�d*���
R�<ӆ�L�z�K3��~F��q��P���=��N
A�h zwA;6N��Zf�<�,ޏH���1D�{�:dن,�v�<�  �2)�l��#�
;XT�a��v�<�cA��H����E�!v[*�k��j�<��V$T���_��W���;#*C�	�!��	9wG�)�E��+rC�IV�V�©ǧ1p�����>
�B�I 螅Qq�UK���#v�����C�I�8`�i��,�s��˰��!��C䉮FDD��4��;2
��@�`�fB�I�rO���gc^�oA�zFCF#.��B�I�-�q6�X�?܆(j��E�*�B�Iɲ%8���F5�u�Θ�K�B�)� �����B�IJ�H��C
FU�w"Oְ�A;f�䡈 �?'�ִ��"O<�d�8y�����lA2�"O´�� 4]qn��w��D44y�B"O�c��
r���I�ǌ�M�u�"O�Y�R'�6z�FY	sĒ�7�i�C"O$쨁�������cV\�Vq34"O��tn�e��!T�&���"O4�Y��Q�0ոd���_�S���!w"O.}� �Y
�pe�@�S\:��"O\�	m�>P��	���]xN��!"O�h�"!��|TxY���TB����"O�e��9X�FA0�W)`<��"O��!W�{�>���@�+w,��"OFݡ��8j������H4n��"O"��C��q�z�;�'�}y�"O��%	�K2��f�$a�
���"O�y��JPb|���EȌgѪX�q"O
�C���_�D�EoJ|��1j "O�L[A)�d�j1I��K�C�� 
�"O��I�z�:\��PW@Ƶ�v"O�ܲ1#G�B,A�-O;I\"q(u"O�ms�F��=�P1�c�N!THlP��"O����L
LQv8h�*S�)�f"O�%�ox�Rc�S����h�"O%����+��]ㄦ�K����3"Oژ���ĘY�$�'%Z7Ic$��"O,���Nb��	xઘ� �T�@p"O: `���[��Ĺ�ˌ;Y� �"��'D�'���ʆ�Nx\�EK�C?8ٹ�'vnѹ%B�c��Ĕ�?�ʍ��'��	���˭܂��b��A֘��'�8<�q˜�_��Lj;��Ԩ�'��Xv ��.>,����5ݪܚ�'���%�W�}/Lչ���#Ċ��'�l����	��	��A�f�����'�,��!K	r��Ҥ�`;><��'�xL١!�Q��y;b�a�P �'���F���Ҩ�ZF���'�fȑ,������b��KE\��'�\���锌:�T�
�,%z)s�'��t�Q̂�?J��G�\�"�^�	�'ռ��dZ:E��16&M9!�����'�x��эE5x|He��E��Z�J�'h^詒�AU���U!��̌��'˾���,�����#�	8䄱�'qV�3E��4o��]��@�1W���C	�'�<y�Ą���*Ј�&�"�)�'Xn����0,@NP�@�6�	��'�����Dp��G�����'Dp�������mքr�Az�'Lx9��ER�j��	���?r�:) �'�0���MW�uEn��D ߜr 	��'�d�Yu��4��;e�,@��)��'~�b4a�+6�!��f	h�b(��'��@�sK8P�ħ\��\z�'�(�k�+VmR��%GI�A����'-����#=���[���N���
�'���Q�AiF�#&�Fi�U��'-���ծف]8�Ⴃ�<<Xj���'�~��dɓS�#�cT�-P"�:�'���Ʌ6���U�(~>���'_*��'
U#++�I��	ÐOf�A�
�'ڸ1�s�A�)Ď�H���|����� �U��	(�ʴɧ��&5�೧"O��0�BеLLb�I���$[|�s6"O �H��K�B0��O߰�Ii�"O�~��#w��a"�� �yR��|����kq�v�������y�a���"\x"�Q�X�:亅���y�Cy^�@w#G5VrAX&��y�g��~�txt�W��J�`U��yrC�;�@ܓC.�x�с�ŝ�yr	�#Sz,��i��,����#.H	�y�޽F R|����bh@R���yB�ʯ �\��#l
�B ��!���yҥ��`��M�&:8�A!���y2!Ф4j
@����-~|R�d��y�D�$?��騦G�QA�M�7 +�y�oU��.!�ʓ�u�@��7���y���o���F�	d�\H�E�y�d�+�¡�%�[�i@Di�c��y2h��;8�`� ӢbӔ����=�yB�Yy�0�2e)υ�>�;��!�y�K� ��:AKR1Ttж	�y�$T �~��7L�7+{j�c��;�yB��"Y��	�!�V�"�]�C\�y��>po"}3���h������	�y���y��h	bNG<(�
�:sdڂ�yR��0\��l���̈́mJ�RBk�y�
R�kN��b�7~Aa˕��yҍޟr�\J�'Y{K �x��E��y�c��HM>��i�4c�h��Lڤ�y���i)�P1�G��n�4�0�����y�k�x���y�����%aծ)�PybI��>��Ur׈��C^U:�*�e�<I 	� ���!��.C�i9� C\�<�@���J�d�p�̌�U.�T�<��l�
J���
�a7��(�OS|�<13 ��t�^�Z`a�5c�B��c��M�<��(.	d-��H�5/ܤ���H�<�� ����F�4#A�-RaSY�<i���Az����A�E��)fOp�<��9WڌpA'Bi��%[E�Ik�<�ǬՁ�<���~0��F�\�<�!�U��h�Ñ3V�T}�JOq�<���]�3*�HUG-v��Rr�/��9�O�,i�K�HF
%�C)Y��lհ "O�##b�d�t��H��?),Q�u"O� �g�"5���� /$���2"O�F�%m�V,Q�d^�f^��"O��)v�Lr��I4Y�6[Є�!"O*�P2��/w�����[E*�	�"Ol�Q��0u
�CR��4!@��3@"O�@i��T�a�d���T�d-Au"O6ЁT�QP�03ς�nn`���"O�� d��_����@��<`��Z�"Oh�÷�l��A���>u֥��"O��z�d_���8GE�	e�Y�"ON��--ּݹ�-V�O^�X��"O�iGh�k�u1�QKh~�I"O�LA�B.L
���#�S�?c6�#"O�H(��C�9�H w���:ad�R�"O���0	rxzܳ�NT*P mz�"O��z�&��u��LB*5 �AY�"O���b�H�B4��.� �"O��1��ڶFW�8	�JoD�sG"O��{Cʄc�y�Ѧg�I�"O� �Q@&C(q��h�r+T�)\rh0A"O�-�׌K�!�>m�p�߷��b�"O8}���;���K��9�@i�"O��Po�\��diF���ᔠc5"Or��a�1\����Bж@��"O��C�����f[c��A�$"O~��$i
�TbJ�#b@�2�9Z�"O@T�&� J$�D ���]��"O���g�g��p�ѫ^�"���"O�)r�͏7&� ��dL�y�Z%�"O��J�޺T}R91u�ƌ[�����"O�"���w���$���4z���G{���!;�T�QD�\�U�D @��z�!�d��E8�� �K\���#Z��!�D��n��q��S��P�����B��D�� �1�A =�\ȒP�,&>C�$T.��6��6<r���N�fL�B�	:	�ܠ ���`-t�s1���c��#>����h��i�"�ڦW���T��Q�\$BE�<|O��#����;���p�RW��+g��ox�h�i\1e��T���	Y�*}0Fa2D���PX.��@�S�U���3�&+D�hP���7���4��18�t��Q (D��Y����|�&�X�f� ��%D����O�||$a�"ӣ�|1���"OX�=�,�:4b0$��M�X�H��hO?-��9F�<\XTM;s��(�J�JO�B�	�AFX@ɌcHZm1��F�B��(�Y�#`�cubx{���]�B�
Y`���R0��0â�ȟ+�tB�(.U�������6����+8�*C�Ʉ^,F)�O�� �/P��B䉝acl�a���~�B�s樅$}��b��G{�|"L���!�3H��㯐!y�b�'IZ|��`��(�N�<�� K�'�>prc-�K����Á3���'4��"S��\Cά���'#�h��'F�̫PA�RQ��pB�Tuv�`:�'S�p���6L�p��˟g����'���5��i��̖�jV���'�,SQņo8�Bd"iO��p�';�Bg�4�X�wLW��A3&k��y�CӲu朜J�f3���kH��y2�۠G4,Ҡ`��V���GH�yb��w�M�FK�&#����怦�y��W��h��1���S	���yb4h����L8K��e·��0?9-O@��i\\x�\$_�|Hz��Dy��S3�h��+N�jG\ɋ�,R[�JC�	+"��Q��%Hg �A7��҄C䉡/�~s�;I>4e��0ufC�Ir�<�G�ޏw�0s�hX!Z��B��2#��R,�>�α�6l�$�B�-�έ˱@۰t����ܝ}���l���O7�I�bw���dI��~�!V#ۜZ�pB��5.����A�c�r�3��[wC䉧 �n�pJ�b^��U ӟ��B䉯+����m�y�j�CŘK�B�	B�@BO�1(�2	��%Cjh�C䉎	�i��K&qa	�@" :��8�ɡC+�0����S�e %%�4#����hO>}:uM�j	T�7m�A���l;�����A7Эc����h���Qc>4��C��Xz\����-eP��G�$Bn�C�)� �=� ���-�����H �o\�+F"O8Z�Ax*�d�g�""b��"O^���
�U~��	���0��u3W"O��
dEe�� ��|�e"O���i�" }2��(foH@@s��l��	�V�D]Y�H*H���{�J��D"C�	?K��9e!B140�1 �ȕ?��B�	�M�� S�"�rr�`[�eU-c �B�I�,o"$�UlЁB�����b�̾B�	"M��d"�(W�H��w��N��C�>~�r����'�Ј��-L	�C�V�Hz���b�{H�����?������|��PCT>U�H���A�,�!�D�/0�X��+*|&)��y�!�.��!r7"K%fFh���C@218!��1���A"�;^I��Sj#!���u����[�b��Pfº!�d�s�1�4-�s����k�	lm!��50������!��8x�k+e�$"�ī<�|�'&MB�E��!��K!}�
�'b�:�HQ�b�K"�K	�'y�1"�'��|�6����*��eJ
�'�,Y�Ci�+W�4UB�$G�(pb��	�'�rM�pÀ�I���ӄk^��'�d�	�)�"Yk�x��)R!^���'�v,i�C�bcP#�ϊR�T�'/�A�)�<Yg���l�� �,6R���/[d�<I�� ��XHtj�?�.��Sn�i�<�QʌLq��ǯǄe���#�h�<�2��-vشd����H�k��Ra�<i�-Ե� (2�4jBȩ�\�<�׉T�`0x�y�`��58Ze)�WT�<�K�d�$i����m�*�چ ��<I�3��h4��y�����-rV�]��^v�`��hܶhx`)�"C����:�	�n�
QB�]�B�L@H���`�R��I������F�8�Q�ȓ#��`B�U=#�<	K� � �x������I`�	j	 ������h����&NB�	5z�A5c��.adA6	mB�	�MY6A���W��:`��c_�F��C�	%(���`-�+Bq��V ]���C��/�:dx�M�)���R9MfC䉧7���Vi�!&
�!��Ϩ)�PC�	1r%��x�13T��i.I��fC�ɭDdA��H�m��#I�1�F5�'(�Ir�)".OЩ׈��	^��B��ƉF7^m�d"O\�� �`�>�;e-� J�]�e"O���ǘ�{w:py�<`D��V"O��2�*�}m�l��-c>���"OP�!���j@9�X	
���"Ox�+F�E�%���h@��)cf諰"O<]z1jP7�&�t.�'�b-�2�$'�S�'/���!�BZzĄ�\1�"7�#D�XQ1fлE2P��4�����X�#D��0�� �H�Ι�͔$f
�#D�0�� ��u�<�i�H�U�ޭ	�=D�p��H8A�Q�&�ĬM���q�J-D���a��$� ˂���{���t 6D��0��sj������@<̰�4D�<kBK�'�`����j�r�L7D�$h��<��E��8n�*�cU;D��8��
���tH�5-��s@;D����!�G.TT�W
�/=@1I�6D�� ��qBK�9\ظu)�E
u�B��"OI��9�>1��C��w���"Oj	�4�"r�:�A��Tlb���"O�aM�=\wX�JrF�FL�ɗ"O������
�| �1��v>�eK#"O����.3J��A�sm"w6����"Ob����S�!��lG8c!�"#"O� ��B�K�I�4C�sl<��"Ov��!	N]���oF�("O"�;�*P��l�c��#y	T�a"O�!1A�	��`��R?z�ġ��"O��h%*��ZXI"��׽��MKc"O�e@�IX�PdԒ���Z�
H��"OF9[�]Y@]�Sc(|(��"O����*8�8���O�
Oܑ!�"O����:�8�r���0��"Ol�Kb�s�r�*����z�H��"O�D��e���rI&,�Όhr"O6�1�j�q��p0&H�@�pݸ�"O���b�F�%�pb7O�W�M; "O�a��X:����7�|`P"Oxs�	@Y���Bv�[�t$���"O���h� {���i#LM4T]H`�r"O�ʂoN�[���8ހl�w��O��D �Ļ<�|Γa����f�!*'�p��gP3#�Ɇ�;n$DQ��ۯG:�qs��7�,�ȓ1��ɐ��1�a3r�ߍZ��݅�5(�l	ׂ�rqz��/�Z�ȓGA4%���ͯt? �����/|�����������e&P�0��)v4ȇȓGt���%H��^�����,w,��<�������O�����)K����@IO�r�"q`�'��
�%�@����Giٕ;<(x��'�@#&
�:~�sP��9"�NV�<!�j�>!|:}Y�N�*�d	�`GO�<���  �n��kZ�����eI�<Y�M�S&�E"�8,�Mx@��I�<�U�_Ā�����v0�����D�<�a��@�;F�аAT���4��}�<�&ǈ�^�0�`��4��6Eʂ�yb��
�ixw�$,�b��D�Q3�y�_�c���RC��(�hh�F��y��D�A��Q���,��E�R,�yB�RFbXT�◬a����Ǒ�y���n_h<���9w+��,P�ȓWP5���(S��!!fU�0������1Yqõ5��¤n)�����&���e+7d��b��a��хȓo$�Q��#F��,�3��a��y�ȓ��m�Eu��d��AB;P�4=��x�l� �K_!SC,�'Ÿ!Z��ȓ�N�a��	4*�`s�j���Sm�s�KJ�:<RwaD���ȓ����s
6�)`��2tp I�ȓXo���[=>��Y��G�&!�2���[��p)��?-X&�l��X��%������^=�r����0�&$��f�}�󅃫JSht�CI:�e���X�+#ڑ`#�Esq�@y�ąȓg+戁5�l �(�G�tY��}edD���1Y&�tJ.ћ]1�E��lXW�@�]ul���Q(Ҹ�ȓ<*\pҠ�,y*�4�ٖ+��ȓr-�#��p�D�󶀑���)��S�? .-�$��&+�hA1��p��"O����DZ�CX�J�g���|�C"Ok�Hte�����@�&��rMTj�<��ێ�R�����pʘ=S�b��<9��I	H�;�:��m����}�<��DA�e�� �Q�G$.������S�<�C��I��$z�EWu��OQ�<9��o�� �S��z��J"��A�<y"˺���2��^%�Eb�+Rr�<���]([Y�ċ6�P�Մ��$�m�<!�� ���0#���c��Qa�d�<�V��=��I�3�����h�G�<�U@L%F"0s�D�2���u��D�<I�Q$CY�1��DL�^���i�<I���<�������z:�4���\�<�PZ�0�@���\W��2�CDr�<���f�
8���4���P��Vq�<9PF$^��R�F��R���"�m�<�fۆ/��8�aT�7�<p�S�Ja�<�DJ*�bPJ��Cr��ǋ�`�<��ٸG\�9�eN� 7~�1�c�<qЈ�aB@Ha6�7r��&gU[�<��iҾp�Lm����9f4Pr��ZM�<ك�PCv<+GE@p�s1OH�<17�Ҝn�d}r�PƬ��%��A�<I���2�)�V�I�X�yrgP�<��E
{ �8����4"/���1#�z�<�`��!+�&��T�8.B�ȨRdB�<�t D�d��%��3
V�o�V�<y ǂ�:jȋad��C�f�Jլ�N�<��]�?�4���	�cD�����U�<I'��iBDѺW��'^���Bk�k�<�� ��V��i��B�K�԰�C�Fk�<Q��;q���Qe܍J���Z�,Sh�<Y�L��JӴ���"v�EX�+L�<�	G35��Q苘0R�@���p�<��`�2\i�	��
��c��KF�<�fe޾ �ܴSaB�*,���3��B�<iU@�
xr��D
��L�pt�B�J�<9Wʔ3��l[��O;YA}��M�B�<��,�l�F|N�;F�8g��f�<�ômY��[��O� �Cg�`�<��bW�T�<�2U��'�h���Dx�<�����w�@$���R�*pd�gj�<tm�4&��+�����
m���f�<�C��}��\�MW	^|�lyS�	J�<I��){=���4K^�i���
skI�<��h�uO�Xɒ)V�P�d�E�F�<	����$Y����%K4m�6D@�<	�N���m20�׆�}����e�<��	��(�hA�ր\,ٹWdc�<	�N��`/L�W	��ك�\�<���	�t�1��~��E�@o�U�<�t(H�q�8]�E�����`SE�TH�<I��)���dGQ8R�d��_�<��J\2/�<q�-�7xE:��i]�<qGS��ޥY��O*<2#��\�<)⇞C�+�8�넎B�HqC�	$/��Q���ya6����6!�B�I)&�X�a��O�h��Mը
-�B�M=��H6-Dv�P�%���3ԠB�	�;�����/�4$~�:�핧5�>C�	&R��E#��D���Q$��oFC�	�<�������1[?���f�ÂYt&C�)� ��ʗ �n��� q�Ʊg�HQ�"O�1D*�s��hÑM��$���"O*���ٜv�&�W�V\(؛b"O!kS+�pJT%95��&mm0�X�"OL�Z�$�|����#��'b ,�
!"OD�8�IY,�p�tE�	����"Op9ȑ�E�\Z�h`�ʼᬼ�5"O��"���3��xQ
V�h�8I`�"Ol [Tg]>��%I�.�&rӊy�"O<e�u"_g�l1u�"i`Ic'"O��'l-��� 3�:��Q r"O�l2�0&�h��,����a�"O��1��U<���g왨w����'"O�yp �&���`�Ū
��!XB"O��O0f�"�� k^j_��R"O�)
�Y�s�&�1�LJ*{�`yV"ON��kM��b�y�n����]"O\�k�'ޫw��{$,�W�,! a"O��ha��=?���R��ܽ%�`�"O�%�R� ������(�d-R�"O>!Y�@�kO��K�F}�IY�"O�p�6L.F*h;`_�tx�ءg"O$taf��?0�3䫍�4?<�W"O^l#���1�����a�.,��B"O���hX&j�Ψ0U&�<�"O����  �.܁S��3��u�"OH\�3��L`d9�5�L ~�fd34"O�����A�Jx(�s��'-<x�"Oxm����H�R]����Q#^�Q4"OJx�*
3L�s�͝�e4��s�"On$�A�RE�:���,�L0���v"O(M)@�,C�������f�°�U"O��3 �|��e��z��h�F��z�<ɡ+�.z������ 2��xRNLO�<	�l��u�]�f�|�M@�JL�<!���<[]�����xl�KI�|�<���E#x,ب;��#�" ��N�<�퇢N|�S%Y�H�B2]����t���2C����Rx;���v�<	�ȓ�\�3�+2z��K���D�� �ȓu�:$n�d��`S��2H�ր��
�j�=x�����-i�`��
Z����K�($�0��R(�@���twLi�G����:���@�Z���d��p �L��@H�|J3�� hB�ȓU�:�(��>՜��f��E�ȓm���J�9_�=�A�8#�|��;ՠ��G����Xe�Ʒ!�:����J5a�*B�ؘ��*@�)XH�ȓѦ�Ac� �"�26�J�>
�]��>�zQb��?A�\H���ΩS���ȓ9�������B�8���CP�dY��)���^�V���W�x�ȓZ�|lCB�4/BiJ��V8)�ȓH��mIA�Q,Լ@�/\`48�"O�8���EOt���i��M`*��e"O�4�`���K�(�r`	�JZ-��"O��2�څ6F��'�N�=$�W"O�<�@�U�/=�E��g�QX�"R"O�`'k�
y��2��/k����"O^�KG����Lr�%�2h�,c�"O�a��H*���EL+@{$�1�"Ok�&p�V��F��/y^y�"O*\ F������,Z'Ķ�JV"O� ��Dg�
A�,	Yrk��>���@"O�E�S�φw�Z���CA�\�jȩg"O2| 7�S+�>!��)`��H"O��"�O4C|�16��zL\Hr"O*dXBL�2	�:�!��B�9r,�"Ol�sV��1v���s�J�h_����"O���AL
E�Ĵ�r��YDlZ�"OΔ &gN��l��Q��9�"O��3wL��h�z)�CН5@��@"O�0�w��5%�něr�@�&8YK"O,ycVH˴&��Aqq$R�_�lQx�"O(�:QF�s� @#�[��v$��"OH��T<-���Y����"O�8h�-�"u()����p;�"O\�Z�b�t�6e��"��CF"Oh����5�z�(+��L�7"O>x���>3;��ȇ$I�)�2��"O�(�֪.Dʌ��ש;���rv"O�@s�Ǜ�;�1�$!3#���؂"OT�"q$��j|�I!� �E�x��"O�PQ��L 08Vm�|�"�"O���'l�(ת��F+�jJ�T"O<5A(l��k��ڽ�W"O:�(n�-?�,����XDJ0"O�5��E~ҔA჋E�qb���%"OF�2� �{��$��4Z�% p"O�Y��@�%�P5{!���di��"O�m!�/��x� v�`YH9K�"O�1)t�[1
���ңNA ���D"ORP�N�J=>�z�h��H(���"O���¥S�Doܵ!a���>�J�;S"O��ʋ*o�	Z���vє0ˀ"O|(x�"���!��nI�c�¸�R"O�H��O+~O�E�|�>@�v"O�lc�4�;A���
�2�sc�C��y�%M�+�&�0�K�uz�@�P<�yr	@��+�^�s�tyXЁ �y�a:czyR6�%e��00���y��T�k�N�H�ֽci�	�$���y�G�.B�T��]�2�����y���|���hs�W�U���e�	�y  I��0�*|�" ������y��ӰOi�Q�g��zߘL�t���y�N��7M�e�Ƈ�F@(H�V���y�̙�O�d]�4*_<:7uZ���yRI[�mil�`e	���H7�yB �N��-Y�K ��(4�˲�y�(�a��к�G��~��d�6�
�y�+�'_,��g	��pL�ĒƣQ��y"�Ú̔�2��$tN*�&a�#�y�~��@���@u��2�&���yƝn8��B��1'�A#֤V��y�lS&��ӏ�0�*� ��Y��y�퉻r��"D"�
��D�.Jp��'�ti�F��\�X���	�'*6t��%6����,?w�$I��'`XX��C�.����W�C�v ���'����Ξ)�)g#�=�.p�'�F9ks)+�EC&-դE�����'$zɁ���O�訑U̜6���'��L�CW"J, \�4��\���+� b㞜R�JH�Y���X��]�N�}[t�6D��c'�;!�|�T��Hl��Z/2D�x�s>hP�S5���.���V�5D�� ����9r����a̺,2�A���	~X��P�Wo>V��W�C�B��g-D����+�T²�k��#Xtr]�GNx�$C��D�L�S` �2�P@I��{��{"���X�kӅF��Ĭ��Ϙ:�!򄜏.P~���)Q�6t@�HH-�!�$�~VU@��S1����&T<m�!�d#(�8�5�F����D@�;C!�d�w��Хa�I&�IT��'&a|B�iX�b�'�4@ɣM�-�^�����+ccx	�'x����P�MT����ϩc�BL���T7E�Q?��qH��7�X�*�.Qa5�Ƀ��<D�d�Q�R�~$ u�-��U0��w� (E�)�=ź�(���0�XQ��H�-�y�ȓ�
u�g��	�݀��n�t�$��E{����Y�l�"��g��HP�ʘ��y��\�vj�Y�F��6~��c����y���3	Z��3''�?JT8eC`�3�HO���-��.%*#���2��ِ	?%������+քڎ��#A�>ښM��F����a�0�b�
���=C�f(���tSd脚F�49�a�Ѝw�>��l��`��c����lFX�<ćȓ`]�q*�/W�]iv�V5�.X��k�� ��+�#t�0�s0+��*��ȓ6�*tBi��X�> ��A�3����N���S��s��ؒP��!m�H0���LM��.c���"�z	�ȓH����TL<���₲.L�ȓ(��P"���H��xT��E��m�ȓ~	HWcH H/���l�8�ȓ)�f�Rsa(U.\�c�*�&:�E}b�2��iB+_cȵp4o�@V�B䉴/�xx�ő�W��m�RHC�:��hO�>%!*3;W�4�J\�Bֵ	E�0D�0x7�"oҡ�	�"��Yp��,��<�O��qd�1eM����5�JH+�"O�ab!NO x"�����Z=4�$(��"Ob��`
*�VРbׇ4�h��c�'��<� ^w��Lj�낆F�̅`W��I�<���#D�	��D*8��K�jWG�<�aEL;d���)��� \^��	��SY�<�&m�<
v ��"�34�1�HW�<$F�'.�� �$�	e�BMa`LTH�<�$D΁�4��0�W�6_|�M�D�<!�AP9	,RL���8�� ��*�C�<�Ո��:pТ�E3v�������[�<Y��!Ċp� 脩,�${��U�<av�N�	&ʵ��Ƥ1H,ūH�<)G�X��>Tҥ�Y}��T�ßB�<�� �c:��y���&��0��C�<����^H�kS�u�`��-�V�<�VT�\�q
�iǱ��(Pi�<���טc���҂�-M�Gg�<��MR�i:~�����uZ�+���a�'Uў�')�ɨ&h�T�(�P�=8Qzхȓ#�$�
2�D�	ݸ�b�F�n@.!z�4�O?�I�I������D�$�Q�eK�B�I�+u��`)ðinj����3�Ԕ�"'D���7�ȱr\�ĺ�� �ʣ8">�ڴ��1�ħGU(���qє�e�U�*��U�ȓ�&A##덲Z�,���#V�^S�iE{"�O[���G`U53JI"UJC�I"�y	�'�MH�c`�*��9`����� ��D��3zYQ F&ؽ6��4u"O�,:�X%@a\�Pu'�2ܤ�{�"Oz���
�	f]��F�+Nn���D"OЕÆ`A�Vo 81�EM�5e�d��"O<<�dB*�R�:��><MqQ"O�dJ"�	:e6H#�R>PU�Ua"OL@�w�WQ��0W����-�"O�\�7*	6	���Wl`� E�D"O�u�Q�G��j��Cv��m��"Oh\�SP�x欝jS��d�,���"O�`�%�
y���"��lF��7"O����Y,V�H������C�dm�e"O,����1i3"�x�Ā#��A�"O��pd��/]d9�b���Z��"O`Y�H��=�)��`A�;D���"O�]��A*g�@�)�=~�lLZd"O$1p��ʈ 
�(�t�Ii�I�v"O�����_θQ��� JI��%"O6H)r�ݹy�&��7��.AHP�"ON�5� �N���ꄀ	���0&"O����'R�o�
���
u$�C0"O��	�i�"p���C$~P�"O0�a�k�~j�XueZ:VH͋�"O��)�b�/"U���D�'�ju��"O2��ޚC����΁�
�B]c"O~�[EF,���V�V�~�qg"O*����K%�v�Y����P��1K�"O�I��B+j�TL��&�H�ص"O�)���(EŊsƐ8Y�f�Z�"O��`�,�+����c�Hw&|�t"O\IapM3�BU)�l� 3d���"O~E�Ѡ�"�R��,`M����"O\H�b`_�8Zt+���7 >�bA"O�p�S��vSd�[���n�~"f"O��٥Q���ؚ��?��qc"O 1��Y� �$��A�8m��"O*�衢ΒW����n; ����"OL��u��i�M��J��4ZU"O���Lmb�h7�"9�6h�"O��[��u��CRF�/���"ON��FA��a�)_-��	�"Oz��m�AC��'ݶf�ne�0"O�Yɢl��� (�Ad�80����"ON���Z�P
fl#��N�;
 Kt"O�th& ;{t�@���'@�E�t"O�q���*�P�w��u�^�""Ot������_2@��*�V���"OnH�'�r��� II5�HY�0"O|}yp�Y2E�����H�%�z��T"O:=ʱ��rT�K��z��5(e"O$���&�b!�B�# Pk"O�L��H-k�.���@Z�j`�"On�P�VF �PR�]`�4�k�"O�4��)nL �*�ք��"Od��w	>Z��iS��ӗOpRqB"O�qSSJ_-��y*3ӻ��@��"O���צ��h
F �� �U�.�V"Or![�:ۼ�aQ�D:<�؉�"O�UBm��1r��)�V�u�H�@"O���#鉺]+�S���>���"ON�o�0Mj*�e�S`��"O��@gZ&Y��a�ƥR?�*��"O�T"'.�����`V�4-�-ؓ"O�hʀNO�L��E
���b��"O� 08aBJ�@��0&��+�h� ""O")��mG�MZ�X��� Uw���"O�+(���b����\)Y���"O�Ń1� -z�\�#�,�(j"l �"OL���C�X��7)��J{��kG"O,E�`�_�N�˱ݻl�hI6"O��a��L=�91/d[d�c�"O6E�r��,{\��r΁Hq>!13"O,�yEٰ[\f�8&z�x�"O.M�tNN� ����`�)d�Xh"O��+�v 4uys双.P��{�"O¬��ݥR�a��*�)���"OF�0G��sT�d Bɇ?����"O~��	tlH��S�d!z���"O�-�W��&���zrIڀf�@�"OT�vh�.n8�p�gΚb���"O<�@ [:Z�&I���9����%"O�(��j(D�[Ӡ�
�Ri���'����mHֈ��h]>����dZ$i�C�	
q/ e�$��|7��A��ִ8:�C�	${Hr��l���;G��s�|78� ���d�M��+ly&]�(lO`㞘���Ζo-�-�U��x�h��9D�(Pl�T����L�q�8`��#D�����?4 �X'Igs`#D�� �_�x�q��c�W+�!Y#�>D�@
��0hr"qy�,Q.o���#n)D�h��! �X�jݰ���� g&D����-��m�H�R�>Oj����($lO��L>��Q�Cj���
F�BTBF�<)���R�����Ui��:W��D��hO�'2�Hp�"�x��q�0 W�9j�]��I�<Y���fk�4
��[W�]�f�K_�<qC��(WJ�Ђ��H��`%cD_�C���O�v��q�ۊǪ9)��ɜ'[D�:ش�Px"�Y'
���M���Ҧ���y�ǙnV�yhP+��hyI�Q��=I�yr�_�>&H��RNV�5�̐A��6�y�<Doj�p��-�t`��m��<	���"�^�sG�P�>v�}�4A	�T;!� :n&!�4G֚W>j�YR�K#+!���6�>EH�K�>=�)�S��5m!�dr���[)_;���"D��w�!�D٢ke4|��9b��s���O�!���	:X�q�Tz��ؕ����!�$�j���)`%[ ����&dX�2�!�d�$A$H;�.��.�U�6(M3"��'|a|
��Z�Z�c�ĉ93/�l�#�$�y�"X�\���,1i|�B���y���-y��)�s͗u�@	ۣ��p<A��$��T�Vl����0y��9j� �</OQ��E{*�������*��<@��:DӚ��S�>�����q��X5�(�q���B80��E{���'<���N>2|h�UB�U����'� YÀ�&��s�FO�^��q3�'U�I�%i�*dc����!8|X�'bh+�k��g@<�9��֮��ܘ�'
�!�7o߸O��5�SE��hA�'�d��D#�z��P`���u�t,�
�'T��� !��(�.�j@�T�nl�8
�'CR-��
!=9G�}P����'m�z�$ԗq���F�"�>d[����y��ϣ<!~�Z1��XV���yr�A_RͰ�A�$x�Q)ӏ
��y
� ��0�A۱ �����(~c���"O�d�L��^H�tE��wLR��w"OFkQ D?\������-I��:t"Obd��j��`�����\�0K��+��D'LO�]�RC���qh�8.~���"O��+������G�,��I�"OZ���P�h�1DEo�����/��M��S�	sy"��/�(���>72ؑ�h0�!�D��"X՚�*�9,`�sӡ��(�!��A�J��H�瑌(!�4�7��=���j�EF�3�H�A�N xF@�h<Gx��'�*��7�0U���X�A
�CTN[gH<�pd�(]�i!���4vev%0��y؞\�=�Bʞ;N7$e3��W�K��])ǆ>��x��ܱ����E��+9b8!cw�U5�0=q�2�G�0o���O�CBR��V�L'A�p�=E��� ��an	� �t#�@��Xx	��I�%O���4͆�5EԈ��B-^yI����\��Ib v�!G�G(� �������Oڣ=�}2R��9,���i��!�0E�R#�wx�P�'2bD�bƓt��L)T+�*H�&��N�����)��$]ڽ�5AȐ<ꘈ�
 �L�'3��0|J&B<��\q �@$ur�CIv�'��x���Uϒ�@X�0.ǚxp!�D�#'�X���@���t�Cw�϶#r!�$��*9�V�
6%�x�p��U�!�D�z��!�DSU��h3s�Ô{�!�$�#����x�t ��H�X<!�DQX-�m���)嬍���
!��B
&��T��I�u���AEO9!��0Q��uS�/Ib�(�3!��'C!��<M�}Qwe���4���,L�~̡�Dw�*�rFD�&uJU'@�Xl�Ek2ʓ��<Q�u"����$B�x�j&a�c�<Rf\�H�5�U(��G����P�F���'U��k��ט>T̑q�؂@��a��'����s.EX���"A�P��
�'�p)���X��2<e�YxB䉪�@��D=|�\1b��S�C�0iٶd1��VYPc��QqbC�I�/K>9��9��̩�B��C�I�5���KG�ġ���,WHC�	�����g��
e��Z1�֤`�2C䉨|V̙�VFՕ1ֵ�S�%"��'+����<L��PjÔz��U䊋
��B�I����cԎN�mp���4J���O�����2$ js��6��M��� VaB�O>���EM�G���W���y���"Ob9G�^��ձr��weH�%"OXy�s�\��L� 6Lt�x0�'s�ɅE �q��F)>�4�*�Ȉ|��㟼��ɽ��U�0c��T%( B��@18ݴB䉶g�-ZU�	��H�
b��6m&�S��MSp�π2�v�9s��$���#�AZ�<ѳ�Ӆ&�6�"����{Gj�V�<��+@)H��5�$��ҲXKv��[�<)Պ��r�ِ��۾K@R<�b�IZ�t$�\�&,�6���@�ƽ3}`I����V�<A�e�
P>ݻ$\�`F�ᶣYw�'�r�'��gy�Z�N���(]7|���Y�υ<�?�2�<��A����*]�h�ґX��Iώ㞰F{J?��e�{LPs ׂ%#4a�s�2D�`۶�ǃ<�r�yr�Q��8�����$���g~���)��B#�4M�`}T�
�y
� �5ɰ�G�2���B�Ǐ�_wN����<D{���$��a-KR�X�k��Q�'�ўb?�+�JW�^�p�O�%7�����i(��1�O�%�ʀJ`��J&	ZWӀ1&��5OR���$��K�	iy{��7�!�$M���f��*�:P�$��;q!�$ܲr&��$�0.�U�3�ѢPi!�L�*�RXa4�L"ɄL� ��4h!��n0���QѢ	����&M�=E��'T�{�,���(V��`R�'��Jd I�Ҳm��Y֖<�	�'i�EP��*�Ľ�g�>���2�'���x�-A=l>�b��AU��'�ў"~
��G�`���D�ф7��	�E�E�<��j�&L�&o�E�i��l�}��֟�0>$(��=	x�*�˟�rS��U-z�<Rg�&~Qj�R��ܢ����Ĝl�<����>ąBTiD/�1(�'�k�<	q��.�t�ɶ�z����+Tk�<+I3�&\�3�Ѝ%wN͉p'�c�<��ƈ ^�Q���ǲ2à�CaG^�<����!?|z(Y�Q�}z,9F��T�<YW�A�uVq�D�Y�d�!�)�S�<�èГD�ļ�ġ^�-��Z	�M�<��@jM�� ��l�<���UE�<�2�$XP���b�L@��� BE�<�t��!����H�~�0A� �H�<I���?[$��ঘ)^�Ly��z�<ٓ��k\�(�g�>jM�a�R@�<id�S"�6�K�ٗ-
$A �)�T�<�%�^�Vt©�E�LhR��KE�<Y��T����!]�P	�Ղ��C�<i��
zZ	��-����@)�XH�<���"t���`��vx�!�)G�<y��O���`��
o-����_B�<Q��^�Lsnt���J1��@�gH}�<ɢ ةqE��S`U6H�R�SK�{�<���#t�nU�@DW&@dj�ç�Cv�<q��>���괇��<t����Y�<qF��>J45㒂�\�2$���Q�<� E1G���z��-�TAZѬ�<���^�oz�1�AEK��\�4(�q�<��@����c˝$��i�6�@j�<Y@+V+,��!A�ęj�Dc�f�<)@ɍ,4��H�5��!p�~i�E�h�<�"�����c�W�&�8��Cg�<��������h�e�Tt�N	`�<qb�;J�r�U熆*f�r��[�<a��D9\����+R�\yʰkX�<Y�gȗ�R�ݲ/_�0�W��S�<�T��6	�؈P�\@Dx0�Cu�<�R�^��fT�c�ȝ"T�1�0/�s�<�-&_8�3`��Vg�T2��[�<��AL�Y�@s���G�P����b�d�3:��٤�B� �1�둀o!�O��/�$����RgS?`���!"O&9�ĭ?ȌZ�'H�8m�ɒ�"O�%&�'bО��T�+ODM5D� �ѩ!P�F5�R�~g���<D�X8�ğ%9�HH:�P�t4��K�*OBxˀf �R���˳Z3�+�"O��0����,��@1B�9J��"O�:�bR�w�I1PoT�^��3�"OP00�V�����6n�R�"O�{��@cN�s�NO$sܢ���"O� ��ie��	")�iS7ђe�*�9C"O��٦�B�}�vxz�aP:��:�"O��X���vb1*ä́/!�r���"O�aӆe�R^`q��=��s�"O؍3T�ZD�%Is�^�'k����y�	��k�*����(Lp�Hr&։�y"�P% �\P�ӥق5�v�ۑ-W��y%/i"����.�"I�0�
�yBbT���# ��Ⴒgڗ�yB���$ �	/��B��1�yB�s����%Ѵ-�X��X2�ybF�72���у��$`"&���y��vT��;��E�o{��n�y��$��Y8�@]�\x�Dc����y"��Yi~�b���W }�dB���y�ϓ�{摁�G-��d����y2���zڬ!�F� gA��"L)�y2MH/:R�}Z���"��!n2�y��3 ͸PL��*q@!�_"�y�g֊X����$x�s�C8�yiýJG`8C�F�jA���5���y�b��\C���ɝ�5d��l���yBbѝn��(A%n���n�y�	�yr�1�0���Ϣ�:(C�O�y2��x׎��7b����L۫�y2��[E@՛��ʝcI>@R䁊�yr�3������^kP=�!Ċ��yBG���dX�`X�~ᐵ�� 8�yr�._vD#am䒰�ЇjZb��ȓ]�pɸ��=��K���zt� ��K��Հ���/G]�$Q!g��6d����M�~�ˤ���ʴmU�y��x�ȓ?0$l�/wF�u���h��\��=#B��+N$,�Jܠk>&9�ȓY �ACqC�qu�l��q�ȓ6���2 L eΊ ����.kB�ȓH
�� �L��v�����"�8��q��}`7X%����B@����x��Ei�bE%;d-��҂I�����&ŰM��\������m�����ȓ6sv	�Ҧ�L8�-�q#��=�t��*4�� ��]:��ݠ�y�b9�ȓ/
:�b�%4���{6$����ȓ;�n4��d�6nP426a�
�.a�ȓ9۪Js)�>PMyI���k�6݅ȓ|M�8#�)��X�� �&�e���ȓ~Z� ���cA$���ۻY�ʐ��n+�e��/���`h&��FOԨ��K1�U���ßly<�C��Q�w�݅ȓk�u�0�^/.��h�@8b�҅�ȓ��Ā�� 7fl����ޯM�D���q���S�G`b";↵�ȓM�N�*��vC�I��wwj)�ȓ"ѦU�4����h�̟J|H��z�jѐ��>�����I-�Y��:���iPI׏rdv$)ui��k�Na��4����5"[�<J�d��]82��g�0�b!�7`���ǥ[�i(�ȓKl�4A7�G�r7.D#0��
x�H�ȓ3�<F�PUb��&f��H6D�|���(Z�H���/<���c�:D�Tk�ȏq8��l�4\Ҧ�(��=D��闌��&#���2�`�(�.?1f�]�d,�"|0��0Kpʨ��P&m�I����]�<� ��Z��'5���HS�t)��|�S  ~9��'R*Aز�,��|�0b�0��N<�!D8kc���'yC\e�2��G.���3Z%c)�L0%�>�P�A��ˎ?Q�]"��)�O�i� D�2�X������j��f��\�ɣ�`��6ŐLD{C�D(^�^,���F>oS���z�f���\�^)��a4)�&2O!�$$x��I+��Q�&�Z�j1.W'�Cb\�1�eZBM��8�J%�_�7'�M;�o�'��Ob�)�2_ Q:����)
�q��K&OȸR�'xgBA0N�|r�I�	�dH2��̞.m1@�I&3�p�ؠL�%w���� ����'f6(�+�)�	| � �aKs���g(%?Q�C�4���1ҏ0}����1"OQ	d�.U2���36�Dj�!�t)T�1� 5�([Ӿ���`'�z����E-�/�8�R�i-G��Ty��@*X��[�4!� �T���T%��^b4���ґ*
�!`�;9ynY8"���q�@�����	sp���P�+�f��C*{F*�;q��`�P�ʠ�ן9��̈d�8�ZqiVJԩ�l���	+B֤#�#ρ$�I�s�e�Q�d�b�;A2�42����S,V�l��&T�W�N�P�aBIP�"��n�@�;U�
!,�T��~G�>�	��hͨ&H>R��8����6|牌{d���O�i(4ApS�����?��0�A�\_����	e�.��"5�x��o�d��@�*Ү8X5Bc�'��D"��%!�b��e,
l
�����mZ�Yɾph�� j��P
Ӂ
�!�j����ˆo��wǸ��.U M��9R�H��4b�q��0̶I[W�0��4h����oʩ���C�(h;�(˃����צ�}G2�h�62��<`�O��$Р����	\ �!�� ���S@��9T��\�C�
�?�h�#T��:5aN+��"�ΰg���S$����C���)@-���\�&��	�k�<�Vy P�C�yr��U�.1���Gy���|oZՊt��w��9�~����x&����!�y��B�I"�N�Z$'ч.ܒ��A �[�8�4L��d�	��*O�CmA�i��@�<A�&\5�8���g�4}�$�J���CB��4���q�`�>qༀ���|I��1^&�	-��A���zsџ\��� Qs�X)�O҉�\[�f?��8e��$Ϳ74p�g�c(D� Ab��rG�o���"	q��S#(�6�r�*��1�J\����>Q���)-u��'��HP���Q]ɧu��
hta�Ti�C"�`�T�yB��4�r��"�x����%K����"��k���OQ>͈��?)��8d䝆o*�8��!D�\���%~f勂���o��]�צ=�ɤn��U���'f�Q� ���!�Ņv5b��']Xa0���.�A��i �d��'(`�z�h w�\��q�Tn���'v��!D�#'��Y1l�;䐅8�'����:�H9A��;X��HAٴ�R��	��S��M�e/Җ
d�����m�#�[h�<)bC�.he����ݭ1:�1ZB-�a?!ӥ�~�d��Ѭ1LO\�b�c9��@"�I+����C0�O�-p�GM��R�J��M4���
-R|�S��'t��B�=T�h q�n�	`e�M�s��]��#<!�+�0~���Pbdݛ��O��"5��(P��K&^m,A��'�@����K��E��!V��\�D��{��q�p�hѰ*O?�	0@Bl�� :"ZI�dN)p�B�ɡl4@��E��qQ*B	+��K_��H�,Q�(���	GE"��%J�X��I�N^h=��Q�dĚ�H-�~J�F�
�b�cBH%g�J嚷�QL��k�ۅd�`�'N8���(<��5�����ɣ�Oz����B v����Bb�#��<Ʌn�?Q�E\�-9�)򁅐9<�����$�O^��L�H������T�InV� ���X���}}Bi�����4ĥ)O��!�A2�s���`nA9�RɒUL�)2�B�k�)$��D��0���Xݲe,	���'?@8	C�-y
l�4��<W3Ƞ��$`� �C�;N佊aF!�qO�S�,�2)C���(��� Ș� ��"���6=F�
	�~��a�Sܧ C¼%a�`����&r�xuC��
�HCLe9V�-o�t�;G�|B����)Y
V4"u! Bѹ:rr`�,���pu�rk'��'�tx�3�EӘ8��b!&T!��H�� �5a�eׅ3̐�3�Ig�B<�Ҡ�lG���a�2���+�#MU@ 8 �@=�p9����6kD)�@ K��
:Pn!B!�#Px��u����'�ʴ�#��:~��$C:@���ӛ?�@bG�gu2:�L�}3L}�Ц6�I�Q,��CH�}�>ḁ�͊v�*p����U��Q��&Ԏ-Ԍ '��K2j)�_�lmB�}�'a�a��T3��C/���g�f�Q�'ɕ�)o���>�S�? 4 �C�������F$r�$�*5��.;�H����ht|J�.S�V����X�(�����m�`��W�c�7MK�f��D�T��HOh����f��3A%��Ly)f�[�W��	tII��X����`U�#?Y��H�N@6�����O앛�߀?��(Ɂ��G[���1�D30�{�GV�r���CI��� 6:t@�hՏ1�1���)u~By�>aS��Le1Ç�h��W'_�VcT��a�B�В#Аs�8�Ƅ:"5i���1�>��R����5G��'�rU@��M(}�,2%*�=_w�'�F��'�.���#ם%1�X�G�O�R߀��#�Ҏ<<t�ibCʷy���{eI;��D�&N��kQ@�7&�ؼF�$h��@tk����3ulH
D$KҮ sʒ�9=�y�m_Bi�5Q��˱2� m��c���2�$e���ܴ
?�6�N\��"�,�g�H$Ex�Չ&r4��m��:/���u�r����y5�!b�	�P�{�/8I��$�iejY���_��0=)ӧ�8B�b%�'Լ���K�2|̘�֣O�9AM˸qJ~zbmK�s�H�8o��u��^H���o�6%�����'��=�W��>�0<�"L�l����N�O��;A��",Ǿ���	[�����ʿ��I.b |�]+�� �w�<`�p ڷ��%���D3QH�=� %..J�a��2+�i�qB�(e�����  d�����l����9O�	@%)Oo<���pb��|iZ��I; �"���G>7q���at�>Lnɰ�'	Q��)�5OJ��cdW-t��)�o <O��&o�� @�u�)5Z�x�u'A�6qO���'�`���?q�Ҥ��`��-V��3�5zw������Jh<)�aP�Y�䐂��E
F=�Rx�'Q�IJ�&B�W�$�%��Μ*��(ˀ�38]��X�C��!�$�|���&A�(n�H1������)��ڝc������<E��'6��0d�X�Y
�{�X7n[�!�'�zE�c��y�z$��ٰ3���'���넃��uȂ��鉡�z}aTgӀ{�XqC�#�T��$�4,� ��V�^ؾ�1�J�QR�$B��e����ȓ<�I�	_�2@��@A�,d�ȓ��젆�]94ld)�^b�i��
X�92��+72���N�NI~(�ȓyS|i#V�+�@a��V</bD��c T �C��<�D�X�]�$c��ȓ/������c������?����#hm؆c�-��\��Ɨx�2��ȓc]n�8�_�=�"��Vɔ�P�tņ�0:����E�Ize���F|踤�ȓo�l��ׯ��9�)r���a�N-�ȓd+���7Mă8׮��'�>L����ȓ���(H�uX�
M�x��C��*D��C��X�A^tqp�Ȉ@_pL0�%:D�T���/a6);!�F|o�P��%D���%$ 3��E���P%L
�K�m#D��AC[�D��5�Ίd ����>D�������G@����!�(�9�"!D���c��e8��ee� ��kd3D����HGAv��k�҈���{`g/D�t��Ҿ*l�\xBʒ����E�.D����D�P��)7 3n�jc��0D�0Ps�H�D�8u�3:�&�p�k2D����� �b�3}�k��?D�D7A�N����Ǡ��9���d�:D�dЇE��O+B<)��Y�3c��J� *D�H�"��#ߢYRe��!IȜ�d�*D��Rc��^T��N/h���%�+D�xB_�GU�;DN]�_b�0�%'D���DC�h�.% ¡Δ8Z���%D�(��Cn�:`��T5@��� T�@��!c��Pq��k`���"O(����E�St���6pXb"O���1ナ��챕�J� ��M��'�8���0!¹土q�|P)�'����o�6l���ٴh�%1�'Q"՛ec�M��)d�F��=��B�)� V\)AA�1i:��f�ú�Z�A"O�!��B��&�جm� ���"O�t�@��8�rF�0c���qc"O@I���-u ���Q�Z�~�y�"O�`�ʀ�>��P%ҝ+� �&"O@TxD��*I���Ź=��!�#"O�M��W�7�t�C��H~�A�"O l���R=L�Z�q��G��X@Yv"Opy���E%(�p�'��)ؒ<Ж"Ofy2�G�	&�J�e�d�:�j�"Ob���܇�ʭ�-�s��e3v"O���(=XxĒ"Zs�U"O>ip�ҁr��!z�4D���J�"O`]�YhT�1� E�~A "O���#���4aҳ�� ebؑ�"O4���Oq�BqB���td@�:�"OJh�E�G.
��z":A� Y�"O*8{U�ތ7��,Q IƱKFd=q5"O�=q�G0g#H�y���"Oi��G�;$��#S!P#")�s"O`y�@"mrd�����3>��A"O��b�Nw�82�'BC;@E	P"O&�z ��FL��C�t� �"Op%x�n�	:y ,hb��?�b`"O���@ņl���^�s�,���"O4�q��qֲ!ႭX�e蒝Q"O�J�O[�}Kf}�@-�17��X��"O٪�)��U�8����2�ZX�"ObaXV�ϑjc$ ��EH`"�!�q"OȅP�Д&^|���d,.|	�"O��P�]�|�2�3""�K	�eZ'"O��c2�4i&<[��_H*5"OhX[�+�$�*�:F�BF|�+�"O�	Ţ��8=T�K�MY�l� ��3"O� `mʡQ�JbBʃ7,��Ku"OT�I��ŹJ!* j�J
�-�f"Ot�sb�D�q��P�)+;�f|��"O [%eT����ɞ0G�|�
�"O�m+ƈ�"T,q'хB�@q34"OԔ[Pƛ�]�%�&�&�q"O|��	3撥8�R�]��Ѩ�"Ot�j��ٻp�@�&,P�Nk�)�d"O8�)'ę�hy��єNyB���a"O"y������1�� 
0$Q��"O��6�K0s+D0�ӆ�8:�qJ&"O0e�Ao� ��Ju�W9b��|`�"O�l�І@�i	~��4�:"���3$"Oے��
A��Y�� �F〰��"O��T�\��`!��.W�$���"O�hi�+)%�Z�95L�� ��3"O���44ƞ��bk�1KTU�"O`����+R�2uYpG�%8����"OMJ����RZĸ�e��(] �"O��3q
$P�D̫s��]=�!��"O�QA!�:0�eB�ڷ5
,aҖ"OH���w����ʎ,-�Lq�"O�հ�@X9&֥Yw�D	�mI�"O�)��� Et��9to�,u$���"Ob���ǐ�W�������"O�1kS(D�5+l��=)E�䪇"O�5��D�c�����$й|6J��""OX����@k��@������m�"O��ە e`��32��):�'��a��K���0uM˘F2Jy���� ��4"��6��iP�O�v� ��"OZ��оn��I&(
	GL���"O���L�	e���d%+Y��������`H.KWqO>yC j9j8�����H^)v"/D���$A�C���C��E2*��я0�$��G7 ���0O�vA2��'�@.N���8�x��]�DA�=�OPf��@1����pC�p�%�T���@��B��
v4���b8�2fŎ;25(e�Qe��=����'����=������!aS�c��ӴS�P�88y��]I�r\ UG�8�l�1Fԗw-�B�	H�~L�ԉFtA6Xt���/�����	5I�`�aw�C�D�bX�N_1h��L��	Fu@�4��P��&[�ބs��� Z�`�M��:�&1X�l��З>�0��'�!p�.`ߚ��'�=K>q b���yPV-X;z���O� �?��脏Yv�x�od�f���DV~Ҧ�Ū�ڧ�TI�T?Ţ�oՊ*����kcSJ�[rR��̱&�� ��F养#�4)�@�'RX`�%�V�=h�;a�I�\c
h�U%�v��HE��(�r��	j����2��"�1�k�(���A�F�4�u	Ê:���7#�2R�aR
�j�4L����/�	���W��l�C�ۗ^��P���Um��J���8��M�5N$-��թL\$K�F1�WNB�3�H�UFn�'��U���!|�0Dp�.�d�]�0Z޼��[�5���
FBQ�@�}[�̚~��M
��*b!�[���仌���l�j5��d�+5tP�e�[��y���*OH�b���YC���'��(	��OUl�fN߻e���Ц�"�L�SC�%EM�T�gA�(	l�e�+T>6�NT��I5]j�a!��0}�^�+��GK\�\��'&�&KD�j̘�%�5_o�u�̄0�L�[` ��K[���3Ɇ��4JД
��5G4����dArg~�)�LЎ%h���R+(���"dKG$K�HҀV@.*��ro�A�xy��$j�ST?�q�I����ǁ1YxZ�*#J}��DI�'�$`��N(Q�h�'(@L�C��>p_6�jG��(N��I��'�0�&�C���l��t��l�9&`Qؾv�8uZ%+���B#ݔ�C7[� 3·����b��O�8��r¦N��ͳeeY�,�H��'�N�r�ȗt�����u�^�X�O����%��.@N�s���<��	U�����8��A4���D/G�9��� fΏ�Iia~���7
�-дυ�AѪ���䕂M)*hX2M[�(�X�'<��`��7hƨ�G�,Ѳ���(��jN�1�(��O�ɢA��{���P��ӥ�R�j�l���)��_�p(����4:e���&�O"m�6�F��ձ�Cn!���U_�4bV�-�i!��X�ޜ��ӺFlڹ.�PX�!�V̺�x���x�<��N�&b�p7&��#�Ux�$_Qy�a�V#|�`F�|��͒S�����93����!R 2�!�ߏ0�I�کq���a��$1O��q6�I��p<�u�ǂ�9�΍=����J�<�f/�`4���%H){ޠ)D�J�<�"_����)�;=�K')HE�<)tB�φ��D+O�sI���.�F�<��
X&Y��Q;pC���x�VO���8kjL'�"~n�hb�@���Fw��+d�Y �C�	0\�B'�8W���0�W�;���	;�έr��0y�az��ͩ �歒��[+C�E�׮���0>"�R=uR��q�F� 9�@P�;Z`19&��?x�>9��'=$����l�d@�Diہk��Ɂ��R1:Xn`����!�Z�?�8�G4ts�}J�"�{̠b��/D� �N^>W�l`4��c���S葒���u��C$�������D̟d�a{�cݻGS�U#D�H!��<a����hL$hC6=� AV0�L�3��x���R�`��$��Pjy�צ��/ NxZbP�Ba|Rb��$��*mN�9 gL�G�XyVI˭t�M	�O�TA��
%e���"!�/t�m�g�	��|P�"⊤L�h�R2m5{��H�cCH���ś`)_m�<��h�?�|L�%O�x෡)>��1��-��g�Jy��9O s㛾E�
Q�A�̖I�(�҅"O�c��/6.u{&'2B���ѕ�Obt�!	��;��z��-�Ƶ�=�O��(����CM��ם0J(x��;c�X��GV�n����/jѤx+�g�(P0���?��|��4���K}�Aj&�͍�l��0D�`4���pX��4<D`r c��i��cӔ��p��s����	]E���p�..�lX��ɐέc%i�
� 0$Z�!Y�\�8<Ie�MMT@��A"O��`��_�n�h��c�4uJų��ݓB�t�JGcA�h���6*��b�N�S	��rd"O>�����B!��
�L�q	�8/�pX��	�H��I)"�H%b�*�9c"��&�,��B�I-��Y "l7\+ł�,]�6�ݾH
X4� Ƃ��=�&�=����-~f0��F
�؞�ύ�\�X����'8 yL�;}����U��XJHb�'�l����8:.����Co�
x)�}����Y��5Dc�O��3�n]�֎��#�Ԝf�����'U���q`J�$�0�"�X����w�ڸ�\@J>����Òh�M��qDt	�$��m�L�ʥ"Oh���@[��Y���0q����7O:h���p>�¤ �� �A��>\𚙁�ߦ����%6l%�"~n!O��1	�I�+A������F2�C䉾n�n}*s`�[?���у7k��	�G���1/!I�az���f�t�&�]�v8n�qX��0>�Q��c�,�څF��1%�jҠ���$,���F2��5�'%DP�6w!�B�$�?`�{��Du�^����>o�F�?aC�Ñ�>�� ��� B�@2D��r҇��	gh �w	� �|e6KB�%z����y�������I�dW����Ը\�R쀃��=(!�$�:YP�혤+Ҳ\�5��F@��D�J�:���Ёr�h���w~�kA��+�pT��H	�6�a|�B�CF �i�C�=*�P��lR��|��d�<��=څOHp@,z|&hɴ��������7�B�����(2��D�j%d�c`�b�dۭ:[�X q�f�<�f�شw�!��ڜ]�>U����i��UC���Aʦ��-O?�9O���id-�f�����/ȡ0MFC䉕t?�4�
�(�,�{$c��nwh��V4�T�5��":az�G�sjE��̖B�,�9q�\8߰>YS�R�q��un�V�r)�An��X}b�ؚb�!�?b���8��=[�vt��a�!�$�NTPc��ڗQn��k����[!�DK�D��L*���yZ�� g,�>p�!�	-I��bs�H8�����`�!��^F���6 �W�1c�m�~�!�D	,F)Q���<�Tʥ�F�8�!���qi� ό�%�P8�*Ͽ�!�Ĉ0�[�"G�*թ���EV!�D�}P���K��X�	{��D�gH!��4(���Roh����@��!��0��% �n�v��\�B��}�!��O
{���[fJ�;A�I����2{�!�U��, Z�OA��A�'ߗx!�dș
t���a�(]rF<(��
�:y!�DD�f�E��=Ug��y"�X�!�X�I|e*��U�\H B�Ť�!�R8U��y��?oM���v�ǚAt!�0��ls�!Ҧ$�Ċ���Bn!�Ҏw�� A�3>L����mX8nC!���nڮY��JV+�A3�M@�J!򄎫y��8���&Ѓ�^�i!���#��0��٣5��Zq䘮MQ!�Z=cZu�bf�/@c�Y[����$U!��ϫER:A��膴W�I�%U!��U�^�Ș1@{@(�
B$�uW!�$d�vADD�fMb����/TY!�dǒ.Z�$�B���ZF�H�!a�X{!��Z�r��MA�M��~�j�óN�Rl!򤂊��q�6��!��;EY�LA!�$�)w�hpI�H��5r�!��J�l�d�xS�"Y(ƘI�َ)f��?y�-*j��� \��� E�M|�<�%ϓkR´[��G�e�",W�WL�<� �C0"�#\�ƈ�vB1a���"O~�*i�C�.�8&G�{i@�:�"O���E�� B�y��u�	R"O*$q���FK�49���<^J@�k"O�R��ȱ46��r����-:%"OxH�taJ�e���i� �FU���T��%L�O��ӕ�~	#�A�	����Ӻ���>���aH�5^�B-qEǛ` ʓH�0��IíO���)��2���`�\�Bh4)�a�7pQ:x
�`�B��ô��
çn�X��.�.$֑��A�/T�&<�F����L��t��va)�.�	'��8H��ф���FA�De�>aB��$�� u��&���.ʧ.o<x�$]~Q`q!��'���F�3Kڕ�W��6D�Z��H��d�S:�����]�J�n�"����h�3O�<��U��h�/R�Ԡ*A&���)sb�E*`��C\�]Tra[�]�0#��$�X8̅���,�SD�'9 �e�ʅ+2��� F�e����U*T�e�b4�<�8�'�?� �5N�N��l�����Ƥß@��o��[ŎQ!��nH��ӑR��j�k�J_�:C�Ð5� 	����Y��E@��?y�� �b�C G�#���C�[�5��閤�8�xd2,L�<y#aK�lMq����cSc��S�f��n�)����ΐ941����u7�X�Ę����퓵�ԅJOV=��!pE�)#¨I��'�l��C� S�b�~���I
�m�v�iV�����̓�b��d! ��p���c�4x�S�O����	���sg�;��]� �HU�=�)�ԟ�O����80��5�p��J��y�L/w�ȒE�\�10�E� ��y���HND�D����젡��W�y���-,�D=h3L4wx��%���yL�_�Dt��P "��c�@��y�N: 
��k�*�fhS�aF�y��(�����̿Z�F�r�@�y�NK`M�nI�f슱����ynW���=pe�0c�xĐ1�ô�y)� �A�!+�
[���P��2�y�+-��iK_�$���J��y­?6	������;+��%X�jԡ�y�% �DNh�"��H�v&�} ��yB
�1OB�iX�mW�T��$�K��y���iw�����7�r���&��y�F{�)�BH�zY:�l���y�Ã\\������C��)�P-���y�I'qD��h�,U�nfn��KE��y2ȏ�"�p�j��f,�k���yR��11P���d'�'ǻ�yb"ٙ�������\��q#%M��yB�n��%����XМt�t�^�y"H�T�C֏��V��a1����y�ǟexx�ꗧ�@���kȼ�y@�:d�0��B��0���o���y2��\e���N�<]6�pB����yr��y@! �2uw�*�y��7����l�{B̌X�ޚ�y��J:#	�t�T��c_I�+� �y�5-nJ�����.X}�8��D��y2S���@��}VD�M
�yrD�MQv!`c��N.�/ʾ�y��fd�D�$�1N��!�gǲ�yr-,E���Kp��Z�"����y�K��rk��� nE^�z]t
��y���^	�J�� d���ɢ�y升$Έ]R�F:jCb ��X��y�Aͥudv�"��b���p�D��y₌�-h4�r�ˏ�����7�y� t���� �!2渜��.	?J�!�_+iْ�y��ɑ=��S��6�!��ȅB��%����[���J���3B�!�D����Q�:�2Y���o�!�� ����0g��h�-?b9L��"Orؐu�\�|u��7Y�ƽ1�"OT�5�6���Rw�F>T�"O� o��z>\���6:�.���"Ol1��@�� ���h�O�p��u"O�;1 ����J���-8s��"O��P4�L+���Ф�[�U��"OV�1���c^x�b��ѽIn�g"O�8Ӡ��/NډI"�E�P��	�"Ov��"Ρ53pP�ca���� i"OH}�@bG�p���t*B�G���"O�YY�猸E�x�Ѕ�
;x��h�"O� ������Q��/8��5H�"O~���T�p�.���L_�>v`r�"O�$���^�s�̠%��,FR"�P"OV����eˈ�X�h^�K���u"O(�7��s}��m)r���S"O@��@��������|)��"OĠ�F�Ac����&b�J
���R"O�@�`h��?=d��X_5ds���U�<Q6) �5Hw$��4�E3a��F�<��q���V�εxPT��g��D�<Yr��;dRz���5l3�#ԏ�i�<���Y&"��Q�M��BՒ�G��b�<i6�
r�;�fG_���"��%q!�ʝ1�,T�5b��h�k�gl�!�$��lu�����3������!�O�lհ̢PM�~^&P:�#E'|!�$���2��2J���@�ʅHy!��ج��	cUb�N>́s����q	!���6��9F��6��"-˻u�!��:_=�Z��܇`v�����Q�!���*ny�h�%�׊|R(�t�Ty`!�W� �D�u�o=M���G�q!�d@0Ȥ �E�(h��4��bl!��#AT�)+�Ȋ2 �>m[׍2$>!򤙨#ZN]"q��X�D�3I:&!�ăewZ�0ѭ\!*����l��5B!�D�gzU�ϑ�fjH�bu��3!����{�(�b���zd��f�� !����m���c0I��J�F!�d �;"�a��Xs*I�v �$�!��M�"N�p��e��%�3!S�}!��Q^p�A��ѧ՘���`ԑ]f!���>8��Zbi�;�Y��(*R!�D�4���*`�X@�P	�vG�=l�!�d�b��x��
��b�%{!�DA�5.��`�o�,<��@b!#�
Dv!�dНgxd)��)@�2�r0!ջP !�8uwu�&�n���J��g�!�Dٶq�45ӄ�F̖�Q�H��|!��x5S��R" ���Ն�6|p!�D��Th�y�Hī�~�A0R�Y!�Zzg��	����m�6�8���O?!�$�!�
����GAC�W>!���I��Fϑ�k����G�E !�6Z��r���' ��H��A!�=oR�y��*��mA8!�$I2 V�E��o	�>����%C��!��%z]x���腴������W�1�!�$��ho�P2�! .U�!�ro\;C!�DI-t�u��H�$~+ �Qo�	�!�D�sB�	�cA�v�M2o�>:�!��^�h�5`�4qc�n��7�!�� �	J�L�a�%�����9�:�"O���Vϲ��-��Z��L�"OPA��_\�=S�.ۧ���+D"O���OċCv9�f����"O ���N� ��:$�ȧ}(B�h�"OڱrE��707�!���\�l;D��"O���X�cY��*W��	%lQ�"O<IkFD�5c�00�(F��-�1"OTL��� �x4aΎ>�b"OF�q���
�n(�b���Z,R"O\��
�J��`���P���0A"O0����ρ]���iV�G�C����"OT�8A�1=,���eH��svfq��"O0���D�a�4mb����Q\�X�P"O��!ʹV�>!Z�NͿ-{޵�f"O�9�3��}3��rG��r�ԛ�"O�#"�GÄ!-�({e����"O�<cE^?E���Q���-��j�"Oح�u!΀b��@��	b�R���"O�Y��m�4ȁ狏�yp��S1"O����Ov1b,�"K�(B̊$�"O��@E\=1ض�(5ȁ�/��`�C"O� xg��<�: g��[� ��"O�h`� 92�b� &�#��,��"Op�j$$�4=�>�+p�F�w��w"O�4����x���k��to�t�"O���uC�k�%�p�W /�n���"O,X1�1A�a�u��8!�J`��"O�ܛ�i��M@t��ǫKc�b��"O��9��S�U
: ���$����s"O� ��eB�co̍��MP:I��c"O֔��\�XaX<�]��RƩ�	�y�o�:�d`��.4`��-qecư�y��2K��� �dA����(���y�D�ut��@o�c�fTk��3�y2������R��\՘�2խ���y��A�=�`�v��A���	��y��2-:���@��Xb���9�y�1i�*)�����
�P�$Z��y2�K�-�8u�1�2{��u���R�y��Wڢ��`�<:�`��.�y� �=)u1N���)ӓ�yR�E9个s���&9��r��H��yR�\#|݌��lѢ�E�I_��y�/�9=�4���]
 �]����y���?lx�cđ��6 ��δ�y2j� <���ّ��$|\Э����y�ʻ`в�D�]&�#�`���yF�/q�t�S�$�S!<��1�U&�y")�ymQ�%�x�bh�KԿ�yb����pZ�Vts�d��'*�y"��lB�ղ2k�sb�!�Cړ�y��x�4`���A{���`d��y��L2r�\��o�?H4��#M �yb�U
ʞ�MYI
����3�y�@"6��e�0o�@i��֊�yB�87��Yp3͋�"��=�6�D��y�U5JC�.�
L\��v�N�ycP07wv$���G/H=p@���
��yR��<YҰ���:�y����yb���d�ɟ1l��#�b�yR���=(���- 2	���yrB�>+����ݢ�~8i�(�y��[/?�@}0�$��TJB�� %	=�y
� \9�mR�8�6��R��a����W"O�uB ��^O>���΀���)8�"O��T@,o��)Q��Y�)�@�"OT`2�̈.ˠH;���y�����"OveK�k[�{�ș���u�܃�"O��bb(G-yfm����+i:M3p"O��8��lo�ى  �O>�B�"O�]�@':T��C�OQ #�h��"O�٢D�'y�b��,,��"O����%��q�$�<W��l�u"OvE�ȸ]��	
 :��A+t"O�9WcF6Kܽ���y��l�4"O.0 ��3�~Т� � |׶I��"Ob\�E(/~ژ�-E�9΢݉�"O2�@�lH�`sힺPl��D"O���u������$�0=��"Oָ�U�	�(�4T���8@Cbmð"O��EC���d�	?�H:�"O@��@�ϖt���ScļQ�>
U"Oh�j��U�G�Rq����;?X@��"O$b��=�!(�=x8�a �"O�)�S��I}��@p �7E2n�jB"O�xA� �D�4����۳C}��"O ��$&�&	j�1��Ȣ|Ӝ���"O�#�w�؀c4��N�I�R"O%���H.�~ru@U,���7"O�9�E��H�ȑY��W�_:
@�a��Od;0���M[��I�S�̡UA�*qډ�G#$P��D�O��d�*���M�,��|ⓧFߚ���NG�FM蝫��RdVc�43'��g���R���'Nֵ!�N�{TL��'Sұ�YBZ�1���f���H&�(�I�,9��D�O�Hn��$'>E�W@�:����F@�f��4���R4��<9�S���d̹{�Zqb�? �!ZF�6Q��xr8O�6���a��z�r���� `K���@�۾a��ݸ�"Ǌ6qh	@޴�?�,O˧�?����?�ܴx�Tt�� F?J^�(�G��lg��	d�|�'fN}�}&�訴�� E� %���۞lLI��hx�,�ӧ�|�L �g}�!f9����a�rU�L9�"wN���O��E�>�F������ ofʘ����Hd=X��!�?�N>��! �J���$q���-֜V|0��=��i(B���O@6mE&M2��"�!֑O��+b[���̱eӌ\n�����I���%��榝��_e��J2�8Š�B�+�9�>9h5g5�Ox�i"nS�q6����af�=b1�
�>�:��7党]H�݁e$Q:���$z2�<!�� ��"E@_l�����H�&�� ��'8���$�<A����dq�<H���5e����a{)�h
"O20��#�?D���F�))Pm�s"����2�M�'G���'��<�iy�4�Mˆ�V�qZ�)٢!
�qP�	�SbP�l���'
ɧ���'$4�T�x�/��Y~�Q�4r6��p��*��=�T�H!p~=1V��<	v�z��@^BJ���̛a��5�'�y����?��4t߆]�r��5bs�����8m)�\�O����OJ��J}���j�du3�7*�����Y��yR��t��灇.��Ls O�=Alm�� �'S d��`j�h��'��9S2n���D�7%�8'�>=;��I̟�����}$����}�SY��-���AH��B-��;Vc�\B$I�b{$Istb��U��9�@@��'[ c����`�4���D�7M(B�'��z��*�t|ҴꞨ�FqI$�5}�F����$�O>�*��᦮�z����M�Ϝ��	��M[бi���2g��b��R+$�j0J��E�(s�kܨq���'��)J��?Q��M�v\Qϲ��e&�b����R��'���U�g�%h��H-0+���wH��`{xp!��
!BHK�T����Y�P�7rtiCeK�y4u)�c5�?q�N��I�,��#|���A����6 �q���Ԫ~t�<i��LG{r� i���!��ƃ	r�siG�.q�D)ܴ>r�����7��'8uTTi�F��DҐ9�������>aq�- 
  �