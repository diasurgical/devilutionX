MPQ    F    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h�]G���|I,N>%�
ֹ�I�<_.11AQ���F��IР��^ʵ�
����:�)��31U�]ΌM$��z�zv-׼���\g)����<~SX�
�N_k��*������%��n$���\�wO��=+z��z���8�W{������`ۆa�jYp)�k��6n��noH��ֻ������C&$�dx|�Z��5d$1��M��;�p��%�z�4��@'�,*N�fR՗(>���Z��b�[�m9�H:S��f^Z�� `�|�K�����y�����+�TU�7ֹ��	�M�%z,x���b�� E�0uǇ�l�U�)�*,D�J�O�L~�u^5�J� S�3�P06	�k��ckC��:�+�Z؉�F�N,��Z�E�.����[�"���\���y������5�l�d��T��k|��5D���DMiج�?�s'v��3�L��{�)Cݨ0���<n�侬(%?���u��9��E��d��bMQ�z��X�'��d������՘�7p>�zr�}E%|?��R	М�N���~1�����
w�XF(=\�ʍmܿ�Y^ud��ȭ7��<���:ZXRa���Enև�?yc�^��`E�p�;HØ�J�\���7��x�͓�&���E6����0�
O�s�y�\�Xa�H��6i'f�1N5)��m�*,�9lk��_�k/;����yHb3A P��"�Zչ��q�����o+���Xa�s6�'
(��2�4n ��ه �.�AN�]3=�e�K�$S��D���7��S��bV\� �����C��=l�����I���XGX����n��0��`������Θ�L}�dr��x:�}�i5=�Ī��y��C��j������K:�+��S�Ё��u�4�d�!%
0�Wͮ/�F��z�9S{U|��!*v�#w �1�<G�4���O>���;���&���<�	K�3��ɞl�\Ї��&�`����]R�������4���|/�iY��K SR�ޯ���~�3j�V:�s����'��~��h��tL��rt������R�������(���KL��V_�ӏ���5�5��k�X���9�&^;�����Xv�+WJ��Y��VQ̻���l��n���9?��cL��*Jl>b�eR�����asL��¡��s�(X�r|ZMo��a���ʸ��6�ȎΖ3��*Rbd��_Ь.��+l�0�%_F���y��W��L$�"l{:��|�oo�Y&Kx��H
�X���0E7	2�˩�2I��������7���ihw�x`>7����D����Mt�8Qߍ$m�l��z@�s���TTtG�h#�#`r��I0�
v3
���LmYbht6�暰�~�T@�|Q��"Vi��Q�)'$�t�H�W�)>��E ����/�҃�N�cd,��j���磇J�)a���K�lM>���1 �t@�Q�.;BV��������~1�(yX��L�<4kL��Cq���bW�lo���µu�(�z���+��"m9����ܢ�m[&	��nۅ����.��c���Zc����̙��s��Z�P$Y��7���E#��
���hɂ�2�����ܝ	W�@F�w1��3i8�L;ϐ���T{�E������j�nnu=�|&Ȼ�o;e=��+�f��뤀���9��~3S�����+�\~��Z��-r�E&��h�y�S��n��Q���)hm�j�n�IR&����ȇ��FU��RF��>�Y�o�-�>m�|����"r�V7bΉ	�o�W]4��2�J4���ca��b['��و^h�O�@Z�B\K��ɂ�g&Ӡ ��+F�6�ExǑ��FGxjH�
T���.C;�a��q}�a���O
K��"QF�d/�:WKg3��G���&@bk�O1m���V�iM�Wx�-4���C�m�P�Um���`z��*�[,"`_���W+�9�qU#���Ts⊉n��z<�Q6/T��� Z�HH$��Kfv�ۼ��T-A;�PjŖ�M�f�AW(�"��?���O����>hV�\}��r�K�!�-�{ռ�i�҂2��6�c���Qj�j��2� ��O�PՁ�#+6}���1��([�j�>�� �s����Gs��ܵ1`4 ���2�T�]z���"��E����*��e
�h�ȿ$��] �ˍ�U'P�.xd Ԇ�~�sB�>8iKIe�G�v����'%��u3��6wݐ9Ulst�jz���l�	Ķp��v�a�j�Ƞ��Txr�)z{��-�$�4��ؔ�8Vɞ����p� #n��O�[N뻌i���?>\f��]����R�D8��B�,Zǅ�l�r��@�k��D����x{exP�n�R3�&�{١B �] �.��P������\����W_�4&�d�>�`�:>2�qa����[���Bƿ2*��t*��g`��C�����!Peo�(��I*���?yX*M�.~���P�^<�`�sJ�_�m/wi$�#��<=q����v��I �GeF�;�ٿ��f 
��GL��?�&[zj�Ȫ(W�� �.y����Qv��`�Fތޮv�	�86�߫�޲���>����l��7�� �!�A�=��̶���)���)M$��kj���ɦ�BψG QN��rFڊ`���z/)��8�󹶈�ND ��z�q�߾���a�~�0_�D�G�)���T/������Ȟ��7����r��N��uQ���2�RS�R�b��e�bY��|����A*&�̬���[6���u��`�Ķ34.ўq�pь�Y�Ċ|�]fz1���Zm�qF�Ǔ��)��$a�\1D����B5={���ؤ��%f��N�I�e�C�3��/�&"^�I�D���|v���k���rKT}۞R��j�(��W�۟4�-{�#��[�E�n��`��Nb*��^�,�=����=�>��������IH�Ugfa�6���t�!m�ͶKNA<<�R͘����,z��*Y�B#;(�EK�wݼ�S�{����J`��389C�:V��H"ˉ��&��g��
�o��pA��9?��P=dJLx� �&�m&���YA��u��7U����)}\;�O���+u�Az��X8����`4:�;
Sa�t�p����k��H��I���R�t���$z�|�l�0�h18CTM[��܋�2ڠ^�`��49ĝ'GT+I �R0��������m�6��9'�GH��'�L�^�(� �p�fWc�Ugž�ZW��a�T���ִ>k	7�%5����P�����?����$]p*�
a��gA��)u9f!�PE �iԞKS�6d����k+lsǵؖ5��ԁ�?,aw�@���=� �$���\�S|��A�Lq��У?�A+�jx�?s��48�)|�MD
���u5�<�v�iz��6#�C��ӟ=n��Ĭ?��������L�� ��d���b��;zy\�b�T������CE�L�Ҙ��pYJ�rAA�%Wrl�X���7�N�&���Y���@_�cw� �F��'��Za1^p8בcO���^�<Fe:���R<Ȕ�R�zkic������2p��H��Ja��q6ޙ�'��h*&#U���3�r)�v.Oo�vXg\�ܴ�Ƙ6O+i�:j�쭨Dt�`��*Kl�z&_[��;��2�H� k;"�T�Ք�qL䝀�v?�j���o�Xw�ˎc2'��u��4���t����RA�e�]�=����7@�ڠ=D�gk7Dk���Qb��u w���FY������2KIҭ�X�p���8�nF�<0οK�{�5��sߓ�y�d�s1��hX5��\�Ŏ��2ڴϮ
r5�%��e�:8-F���М�����K!`�0+�^�*��F%!���f{p+ל�V��X�l$<�G�/-��ܼ
�O��$���C��2��G1�-c����u��B�N�A|d�0�m]-�����|�冖j)��I�-Sm6��4'�~��Z��Wy8��O��MW��#d�tg��r�����a�̍=�.���#!��]N����d���7�x?�5p7	ѓH'��c�^
�+��$׸p5+r{����V,���Pa���n�1���r��E�bL���J���bu�ä�.��7sG����N�.ڜX�yrZ�Y;��{�96�5�6�x\���%���[��_|x.Ͻ]lN#����F�j�y��V�o�&$)\�"�u:p�a|1�oHLTKs�Ԛ�YX��0`��2 �������(^��N
Λ���Oh���ۓr7,��z�DTrJ���o��Q:�vm�3K������n�s��T� MGa;�#�ʄrR(0:��%�g
���h��Y���h���"~��o@�Y㳰�#䏍�,�$b�@tJ��RA)�tPE�*V�
� ����}�Y,�P�x1��WJ	12����|���w��@H1[}G@�1�),V-��yg�ճ+�Q��玨�wDL`�>�  ^#�����,�zc�4�����&4�"��x�e���̩�W]m6E�	!T	����(�.�c�|�Pc;�k����\�̕�]$��K�2�:�n#b�f���J9�67욫w������<n�r�,��r��pi���ђ�ʄE�-���P��5ni
y<���v��;7J�;Ƅfu�����ԁ�~.h��vg͸vM\�V�Z^Օr�ڊ�V�_��0�ƙF�]�����ch��jO�*$�S�����";AFK��bv�x��t��o��>H�|�bԽ�V2#�d����4.M�2��bJ����ܴ�UY�["���4��hc��@u��B�&���
쑢�d����ɂ���5�x�����G���#�(TȬ�;.>]Ga�}t� ��
�*",�dj.;W�v3��-�5�@��j@%g�F�1/�i�8Xx\RD��IX��ӛP����d۷���y,]�:��M�R��9z� U��'�oX�|�f�8< ��/�n�Z�U���)�f6������ėAv��P+�H7<fz�(�f&�ZE��������+\�M��m�)�4-PJ���*�M�ҩ�?�p�H���eY�2鎏��kf�ʞ�.}_��l��(�	��>N�I �u�s�8?��r��Ӱ���T4��.����鯰��郔�+撝Q5����Ci�ߨ�����
�w#�z�xhڢF#�U���iX� onT~��k�>#���K�q��l�v���Fu��w���i�V�a�KJ�l���j��ׂGr��f5�N��e3��ި��Tp�x��
z��-�Y��o�X�/	TV��^��t�+�#��Oʙ?N��������wf���7��+DS�pBUZ�!���G��?�k�R{���x6��P�BZR�C`�y�}1���i�.�T��RCp�eY����Wڑ[&�ղd
?���y�>-ebq���g�� ����22��teѭg�=C�	Ւ�B[P MM(�J1*nP��g3y�m���(j��8����`��)�zz:/������<x��$�q�lI{��e����*�,5�
p4{L+n[?|<�!�\j��(	e ��@6�ʵ���Q��,`�ݱއ=wv(H�8��;���C�����xlU��J�!B�=�6���ʤ9U���6$�o�x��ěB*K n8�0���[���K)�|�8� ��ܝN�ƓCF���$�9,��<�H�k��D�6b��"�?NMD��֚�$Y�]פ��n��Q��p�=Q���U�m�1�݈�e{����l�Q��b&��\�[!�N�i@%�gV���Ά���l�u��"����w|�Qz�+�����Ԭ��.a*�$�m�������O݊�� =V2��:�q�\��f�gj������ӡ3�\����^�<�SH��v�k�����Ÿ�aT�J�R<I�jkʺ��Í��>{�;zʶ���)�`�ASb�-59믱xu��U->����3RҘhD�c�3g�I�6ՎTtp�h�N<�ȁ�:��z�,�+5*�IdB��'��I�wx�S�����`C|"8T^�:�Ա�#p�����V���N��ʀ�p�E	�
?)o�]�L�����{�&�� Y��	uD�4�F�tž���\v,�O)��+pl�z<�8e��<I�~��Ya��p_�
��`�i��HTp��ă�y�bT$Y�`|"���+$I1��BM(�ܦ3z�TJ�;1�4t/'��D;oR��;��:�u��Ú�>�9b#�Hp���R-^� �[ɓ���������U���T��֯"	�9%�R���w�ˍ���~zi����.���*�%���l���8;�u�b��� �]��F��6�\t�_�ykF���0�Ж��Լ],�n�;���J������Ċ�
뢙������km��>�A�������S���~�M\��%@��p%v�1]v�=���nC���b�ns���z8�u����{˹��ջ�d���bCb�zTּ�:�<���vڧ�/�<��pt*�r�$%2�~���N��iN�O<�4� �����.6w/�F�>�@����A!^k,Ñ�����=�<*�9:-R(���ց���c㼿�b�p�P�H��6J�Ň�L�U�	����&�g�����-t���O�~�QW�\�J�~��6��i�.Å�- _�
��*�ll�_}_�d�;�&��H�(� ��"�c�oC�q�Է�<n��e���g%X�L˩��' �����4����-��z�Aۚ]�^��<~�{��K�Dn�7�8��w�b}q 2�*�j��3Y����I�-X}������n�v0����А����N��Md��:�nH	3_5�h����/7ڏ{WE���ʨ��G�:�N����:з���k{����!�NY0�*h�%/�F�mC�~{��,�oæ�Z�ak<I��*���iS���4�-e��z��r���y�ȲW�/E"����\�\!0����]B�0|�䆑x�g�(��S��w���g~lD���P򞩖�(WɨO��g2t�ldrj�{�]+�Ȧ�Ɉ��Ÿ�q��oT�	<��h�5K�V�μ�o_�^��Us��Ήs+�̹�O��V������K�n�k���� ��L�5�Jb��bP�%��S���sB���W���	X���ZCd~���t���B�6�H��L�ɐ��y���_�Z�.�¿l��A�[��F��y>���*�D$DY�"b-<:K3�|lH�o�^ZKn^���4.Xk�~0{�2������"�w�9�X���K9�hz�ۮ�7��aU݂D�3h���j�BQ�dim\���n�i�LNW%T��IG��\#���r��|0�O�@��
�[�C�3Y؏�h��~搴�~R�k@\VY��*Y_�u���Ȍt�5`�M��)�p�E����%��y~u�X�_,0>�k����JdX#��{T�b�]����1�uN@#1�$�VaLFV����J��T��qL����9�![}0�K7�����oI�k����b�Eq��!��"#j�� Z˸��p�ҟ	m�	\(^�<��|�.xn�7��c��_���e����$�U1�-����!a�!~|�'K�[���+j�H)�vS'�m���
���琾��J:�E��'�)@�,N�nd�0���1d];R�ޗ���fP�)��U��on~)��@�e�s�\�}Z�کr����0���Kƃ��Ҹ�H�l��h�Ozj��=��й�T�Ƚ��Fa�޽��3 ;�/to�D�>#��|$od�X�,V-<�������4I�2	��J���&:��S[Sɪ���h]z@�Z BRX���k�����V����4��x=�Y��eeGnC	��TZ�w�I��.9��aF�~}/�G�	 
A�"�Cd��/W9��3�ȏ�n�m@غ��oe����i��lx����!	�#�gPO��� .�V�����,��J�B��MQ09ՃU�!��]�›U�AdG<;��/��5���ZU������&��y�h���QA�q�P��{�Cp{fb�#(i��u ��ER��ˣ���N\C>b�h�#lo-9G�7c��u	҄�r�D=���`(2D=��c��Ȇ��s}:@��j�(Q�P�~�>��� �z�s����=������+�=4L5��ZO�
��y��첑��Q�Ϙ��~^��C7���B�
;�|�5:����<���QU��a�X� 
v�~�� ��wشc�K7�E�=m�v����]ꃎ��z��!��{'l���jp%�"-��,} ��+�`ġ�9Y��,4x��zq��-���ɪӧ��Q�V�6��Nh����#���E{ON��#��/+�u��f�ߵ�`�F���Dn�ZB�I6Z}�9��8�^�k�D�@�x���P�6]R)�};)
��sF����.��ƭ�>� A��n�WUT&��dE���n�>(�Wq�*�"!u;N�8�Q2�A�t�)�g�f`C�\d�O��P�J�(���*�z��Τy��5�d�������`bemӕ�/m���٦�<�-��=�l� I���e�����# 
K�>Lf�?�H�[jf�(ͧ� �/�	���H�Q�`=�Tނ�{v��-8�"\�����\����)��l����!�4_=^�<��_��	5⽆$4
��Y���B��N ǭ��K�Bڀu��.x)"u8m��~�UN��G����9Mߴ���B즟&D)�4�_L�kI��M���墟	,�8���	*T�0t��kt������ ���Y�X�eV�@F������&ymy�W� [<����Bl��,�nj�|�g���B�>�|��cz'�h������ދ���ܣ�l�ڭ�������8�8=1�'�u���~Hf�	����]����3� ��?�^u+��E���V�v��5�!���s�|T���R���jF�Ȭ��S�j�{�s���'�䥰`��b �pXc��}���<Z>��+֎�֘#�&~?�g\R6��(tP(����N7�1��=�5��,�{�*O�)B٠���gwh�S��k�PJ�`�?�8o�w:s����G���:���w����%dp��u�*0�?�X��u�L�ߢ�\79&���Y���u�n��W���t��\�kBO��d+kf�z�<8 {��8����ǻaG�+p����%ۆ�;zH`;��j|�� �=1$��|����&��1�AQMѢp��jږi4���4�d�'}V?�R�f�J���02��$����9���Hk��x�^k�� �셓���K� ��p�A.�T&P1֪ �	�J%�����F�[��f��L�=J����*=a{�{4q����}�u�'T�H� $q��AA6��Ҫka�ǫ��˛����,��6L/������}���7����Ţt{����WM��Z��ÿ���A�����DM�ͭ�`�^�D�v}�Ѣ�Ь�GC.���AnN�`���a���.D���vTxd�gb��z/�����������&���p�*�r7(G%8��\�m��N��y�
�FBXw�}RF�6��{��ܐB)^f@ˑV�h<
<E�6:�ƚR��-���e��"�cޛ-�q �pA�H|�JW�r�'���D�3����&W־V�ۀ���߮�O��:,vu\I筴*�6
�i8C�b͛z��V}�*���le�_��;�f��JUH�S� ��"���J�q���ׅ��`�!�%ҙX��M���'{�5��1�4����&�PvA_p]d��추��-���%DJ�A7z&I�ebg=� ��5�+����u�OIH�FX
ּ��n�a�0DM���������)��ѵdCk��iq�uv5nJ<�����l��jG���Rk����I�:�(�N9��Ҽ������hl!֠�0a�� ��F��e���{���גA���|)���<��t�%=����	�f>�H?��Ӂ�M�����E�c"�����}��иծ�w�ê&a�]���k�D�d������� ࿵�S�v �*n&~G<ټ�p�����!��h�噋&t��r��8�6�0��d9�����[�*\�$��n�h5&	T�	Q��
{;^ �4�������u+�=��bV�׉��N�=�Xn���J�Z��Q�L���J�|�b+rw�Qcߗm֠s=ǲ²����Y�X���Z��Mqoԩ��Y�k�n6|8�Χ���[���� _r�.��Qlă��UcF��Gy����P�$_vv"���:&�|�Ao~�8Ki�A�YzcX&q\0��$2�<��Y��]���i� PX����h5������7"6$0�D����e��Q���m!s��L����)(�T��G�+#�x�r��0��[q�
vHQ�`OY�2hErh�f ~��G@s���������������t���H*)O�BEQZ��@���� ��3yu,kK���<���J��4BCR�'���U�1э�@�P��4V���Ո�~x�b���P��=�LQUt�4�x�c�����/U�ӄ�F�Y���fz�f�"~2p��- ��B@�MN�m� �	�a�?�m���.�aC��G)c8O'�aY�`����$*!O�(��$@ ��g�Bl�,���a���N�P��8�h�@�D�C�}9J���˒�ɽE_L�d�����<n_�d�y1��c�;m���1[pf+�`�1��
{�~$�ޱ����.l\���ZT jr�d�̠�J���O��PҐ'��h��jE`�q��:�c�X��F��������)��6o	 >�	P|_�����sV(m��⥈904ds2��4J�U �R�����[���
�h��@��-Bͩd�\�Α��������Gx������`G��s���T�L���8�.4 a�0�}�grn�
�ٻ"�jqd�rW���3|�m�ɭ@����-]>_��i���x��,�zV�~�SP
�A�;hJђ���E,�X���̓H�90�>UT�
䥂A�����<�<vk�/%��j�Z��oU���6���� �z}A�O�P;V��>ɶf�J�($N�������Ʀ�A�\�N��c�9ǫI-�Gv�RI$�C7�_aU9{~d��[�2���+�ȡ��ʔ�}�n�i>(��
8�>�� F�}s�ϸ�Ϟ���f�4�V���ߗ�e�h@){�ZŒ�F���r}�s����(�ג>
�����t>��lG�<��U�~Y��x� ��t~���S�o)KR`⧸�%v�M������|����h��V���&l�L�j���e�g��G)K�[u��){��jx�Z�z�^
-cE+����e��V����cd���j#�!��|�N���|m�YWf�&����K��D���BK��ZX����k����k�V���<�x�{�P�J�R�RK�����װ.��.��4���H*�3mHW�6M&��d����1�>#��qrB�ݳV8��2��tۡg1�;C{ϯ��ǎP�h�(�X*d!���Vfy	T(����I��oԀ`Ӱڋ/�S���٭<��Z��g��I1 {ew)��*a��"2
&ВL��f?��wvj�b*(�f  2�G,c�����Q''�`�0�}[�v�$�8gl@�5#lz����d[�l�!����!�ݍ=�@��=ʚ���e�$oĠ;[���PB�R �1�f������^��)M�B8�ل�y��NU���	��{�/��m��o�D�ſ�*2��sL�Ҥ���ڤ�wz�DC�˶x�f��)B؃����i�ӟ#e1�l{,����}�&���T[W�ַ_����g��w�b��ѝY!�t�C|�Ǟz�n���i�"��dHǣx��5�{���u���f��ʼ=*+ٰ���m^f�˵�Z���tV3��쏗�|^Pb��W��M�v�e=�|'��.:�TΈ�R2Nbj!n��-���{�ˊ�lOɈ��|`5VTb��X��F����lT>��k��6�޿���Hg�zX6��Lt�[r̞&�N2�v�cu ��D&,���*��B��w����w�m�S�FP��">`�#�8��J:�1#��k^�4
#��Yi�6��gpP��Ev?b�ή�L)4r���&��YRۇu�hzЈ�jN�Ou�\���O_1"+f�_z�48��P�T������VXa�SZp�̉��
M��(H�o���q�oԂ�k�$�y�|X�!d�1I�M�=u���������X4���'�:hRAAO��KꂤY��=c9��H�]����^��� L����OO��i0�k�"�|�T��t֥�	HO�%f[<��Ь����ʜL��a��h��a*��x�6�����ބuʸ�6�� ���<�6uI}��#�k|�y�&����B�2�,2�ܮ1���N���GZ=��͊y��Ob���W�ס`���������pJ�-�D���\M�_��}���9�vx!�,��g�DCI���]Fn)����c�@��y�]Cn�1�-d3!�b9��z
���ჯrՋ�m�]�
����p�J�r�Ku%����	Kd���N����M��y%�w��F�t`�����+cI^at�t	��#[<`�[:�^R��h�1���K��cٚײ���p��9H/]�JҮ������=�9��&!��������l��z�Ov����\�����6�Ji�wu���9r�C*�k�lW�g_,�-;����C��HN�= ��+"���%M�q���r�o�[�\NXM���ߪ�'�)H��q24ZM
�ER��F�A�%�] ���Q�R�k�D��Z74����b�� ����P��)�<�P��I�A�X�zaַ|nWm�0�ë��L��}	�B@8.�d�NR�d�髥5)LR�ڀ�%�E3�G�H���k�:I�i�	�1����a������!|0�}���F6f��غ{����4A���L�<n<p� ����`;	l�c9Қp��(�?��i�������ؼC�sE������]�&���!aM_j���?�x�znS�F���A�~"޼8(Jt��:w�^�3�TϞt��]r`ş����>٥��	6�m��n����M�?hB��	5��D-ॶ�^�6��p4�D<+�Δ�E�%V�Ĕ?���x3n�?��>y�v6�L�JX|�ba���-_��s8N���_�X�N�Z9٨L	���U���6wHn��q�}!�(&_�e�.`,l�c#đ=�F���y�ԕ��M$z��"X�-:�!|���o��Kd����Xၞ0��2��E��с���o'�����:h�%����=7���I-D`�R0�`�QK�.m�G���J��_S~�T@�_G2�1#�[rc{�0k�IvZ�
�T����:YN��h�p��8�~�@ү���U6�޽	�� t�X�C��)�ɻE",�[l��o���k�,�x�S���ӃpJf����B���XC-�\��1��@Y���GRV������&���$�x��(��L����/����N���د���V��!�qQ�{|Z�/�"����!������mǾ?	Һ.�떶��..u#��cS�Y��r��;��Fj�$���#Q��~���q��]�9����<�S܉LϬ࡫c���N]�8ΐ����@y�E:�`�m�b��nZ�M�ȧ�[;����U�f��l@4����~HE��T���%\���Z�E�r_Yٴ1~��Z���;�n:���3�h�	�j������uk5����F�M�s�E���|ſ�o��>�T|���Ԏh�V#&��u�C�)46?2���J�K���hc&��[M�Ev�h���@Ɩ�BHp�7�H�SWQ��Ja�G����x�XD�	x�Gd�*�1cT�S���./�fa��}�T��
7�8"�a�dE�Wo�r3wBȂ$��@N���-~ؐ��´Di9p�x-��u1?�ٹ_PŠ��V¹L0��B�,A�x�C��9��Ub��Ǌ�vkm��3U<�^u/�=���Z>=�n�f~�o�ĥU 7A'NP�A�9B�f��(�񆛫6:�;/xƁcT�P\y��^l"o�-�vI�mO]����:Z�OMm ��V&c2�������ȼ�����}�g���(����>_�� �sm��31K�t`�ܡ�4�ȩ���\�������"!���.��lG�����y�X��j
�e�ȫ��������U�#���� @�~�8�����*pKm�F�3�vo�������/S���2�g�a�|<�l�Զjf���Ģ	S��F��VF������$x���zg52->�M� v� C6V�N��̰\�#�l;��NrnL�U�c�Lf���S���FD�B�qZ3�˜X��S�k�H���>xg�P�~�R
��V��.X]��f�.��#�c�ۈ�p��N�/WK9&}kd���̷�>]q�	؍�f�qB�.<�2�Vt:�g̅�Cvb����PQ�)( ʘ*߹+ݫ�wyD�n���2�����`�� �˺/c7��,�<)jڔ�bb�I�H�e2}�E,��`0
�vL�9�?M~�k�j�?(CE� MG����nz�Qb�@`s`C�x9v9Ö8"��P���0�֪IO�*�l&�A�!S��=Դ(�"X$�9�sd�$����|��:*B;�V =��؁�_�v
ˍ9b)��$8Tf��tܙN��t���ݗߪ����Z��`<D_����!�+~���^Ԣ����v]� ��f�aiub��>���7b�N�"eNS�2�=��x��&/�F����[r���s~���1Ģ���P��]-��$��/�|��z@ƒq���]�U������zհHx���.�=�������-|�f��������/Z3����r^+���0����)v����s����T�WeR� �j�o�C���t{�C���Ɗ�ZKm`PQb��ʑZ�)��&�>��g�Dٟ����igR�c6f6�tƮq�9��N-����Bc����,�{�*E�xB��Ǆ12wI�GS�1�:`t'8�o&:n��os��'�r��Y�ۊ�p�:�`�a?����Ld�����&�� Y�)�uu�����½*y�\'J9O��7+a�!zM>8������\�ŧ�a��|p0����;�zd�H��=����ސ��đ$
T|�I�4�1���MG����	Bڌ�����4%�'�2a5�~R�;9�Z��fp��D띢�(9�=HAp��$�^!�q n+��7n�AU,�F���z�T\+�֠B/	���%!�w��S�<�Q�wR�+M
�s�(��?*�7���f��y}�`�u�iGq�+ Z���7�16�����Yk�Paǡ����c��m�N,�JY�,P��^[�W��)@n���*i��8:�<�;����R��+҄�HqY�FM����j��z��vsI��ѱ�"�eCd{�	�nu��+��F@���i���}��o'dNv�b���z�j�N�;�w���{3ڸ ��m�pŊ�r-��%�}V�DYУ��N����E;4��O59P�wyz5Fo�Ʉ�ˍ�ƣ�^\�/�����ޙ�<{ި:|YNR��S�l�I��Y[cԹ��'�Yp�M#HJ^�JM�,��E���$��ą&Ⱦ��^��g�O�l1�D\�;P�O�6 cMi��΅�l��rL�=*su2l���_��);�FZ��)�H		 ׃2"u��� gq8e>���Vb|��CX���W�'qz&�\��4�������\
A�*]ڀ��줖�#��F�D�@�7�a�Ժhbe c���k����j�+J�I��5XN�ֲ(}n��\0�Zi��i��:��ߢ�s��dyR2�_M�D�5�m,�13��E� ?2�����B�߭�:�r���r��%,��q*�^�M!L��0�WU���F�t�{�'�׈FR�j ��X�<^����zy��˽�~S\��np����3G�a����3���.Q���C��7]��������y�b�x1�5G�S�6*� 5h~��S�F�Y��͖�sɹ��3�tӝ�r�D�����y�S�����q3�ɛ�����Z.��d��5�Z_��A�@b^�.�f)����+�n���5V�Δ<(�s?fn�٧� x�1;rL0��Jӛ�b�o��ӗ�s3qe�h���Y�X֛Z�C�'�m�%K����6rx��]�u�ї���_h^.;�l:db�,E�F��yOoӕ[|8$�-"��X:��|
�o�V}K_P�e�X��D0�_2;�y�p���}�
�Q�\��h�����7C��ZD@7:��x�[B�Q��m��+�i���4Y�)�T{yG�Ip#��pr��j0&eD�c
l��Է�Y���h{�D�*`~cԟ@���jЭ�ޘpqN/)t�r��>u1)&5E�	��vK���eJ��|�,��z���Ju���3�]y���P�7t�1G�@����,Vr6�w���A����Sn9�c��L��G�*Ǻl��	����O��������O����2��"4#h�Q5��29��CXm�|.	4�u����8".����he�cn��W�.�@�́�$`3�������R���xʂ"�����ĕ�GWc�^c����V�󂻐;f��H�Eie�ڮ	���$nU�@��b��;�8Η'p�f�}����x�@��~(H�Q4"ͤ�_\AZJ��r:n��B�E��׃�����D�����h�Dj;�@��)��&[Ȏ�Fc�����db3�to��>��B|�a$�)��VgÉ�S���4�j2z�6JeaP��9��{r[����hO�j@�dBì��Nr��3��'���^��N\xn�_�$10G�x-���T�~���.*%)aW�"}`at7��
�""�x�dV7�W
+b3r����Y@	"ּVS�͝v}itm#x�$v�piĎ4�P�Ã�q<�����q��,II���5>�h9�J]U�����,���s���KT<�qW/[���hZf�j��M�ҶD��<U�0��AblPq��4�!fs��(����qp���u�\���/\�f�Y~�}R�-<����u��9��s+����X�QUg2U7𔾡���ʊ�
}�+>X��("�8� �>��� �H�s#inϮ�2�O�m��d�4Z�}I����肔=Œ���`�!�/���� �͒1
L�H�fJ���T�2�lUn���U� �Lu~ԓ�	h���K��s��.�vJ�2b8.������q��7�Ql�|pj��	��}����}���Q7��J*s�@bx�`�z�+f-� �[�؛�V�
y�_�԰��#��p�߇NM�h��t�F`f�}�q����
�D�k�BA��Z�̜�����y�k���Q?�x"�aP��R��*�\�i�ְdP�.��ƾt��Q�r�i˞W�[o&X�?d�3żg�>E�q(�ލS9��l ���2q8�tQ�GggECq{�`��P�(;ߠ*Zr6݆��y�	�5&�%r�%/�`�����}/�:,�j��<d86���7]�I�e����`��Z
���L�?�~� jwi�(�C, h�"vL�IC�Q�ϯ`̎�s��v��k8�_U�kd���օ����l�� �2�!���=����=sʐ7]�N�>$嘈q�p�B��Z �,:؜%���x�,^)��8�Z�o&N$/1��_��%�ܮ��Q�WpD�����2�|(K9[��"�w����ɖ�������\?@�3-��V]�ُB��6e���X��T�s&n&�Nm�ː[�E�U_��m'��Ӟ;���X|��S���=�|�z�1��L��Ԙ3Iǚ�D������Zk����#�=¡��&���Ȫ�f�q�����ƚ3*�ȏ�u�^0i�k���nv����2�Ť	�TGkR(�]jבR�~x�;��{���"^l�΁`k��b��,�^��dVa��+q>�O ֟�d�T�q�.~g�+;6A��t"��Ի�N(━0�fV�,,*�WBj���l��w�؛S��a3�`/K8�

:����;����������6�p�@��{b�?����3L�<-�-*&�nY�u0��K�`W �E\b�rO��+\@z��'8Qi��y<�ł�aa���pˏ���4���(�H@�Ļ0�7e	+��>q$E�"|����$�1��=M���<*�j���4`E}'N��0gQR�Uc{�W�)��xI�}�>9N�Hܢ�����^|CR �^��?u�`�!����P�T���֛��	�~%�27�'���'��Rx�f.G���9*N�S��W��W��u�:I��g �kB�2�6+���K'�k���s��|��Ԩzd,h).�'m�P���s#�D�v�o(ߢ���s<J���f��q8��+��y,�c����1M��?�x3���vn��n���Cܟ��Sn��fٻ�_q����է-edi��b/wz�㑼�H����Y���e�(�p��>r��%�P)��J�>��N�3���w#uT��w�(�FJPÄ,��a�^W<��*�譙��<�:�RjR�'J��%dc��߲��pr7�He2J����T��sΨo��&�K�g��c�0s�Ol�����\����ꮼ6�7�iI@(��l'��Ǭ�*N��l�4�_b׽;��o���QHē �e�"�χ���Vqs�(���(�Q�Ö6�wXã��%5'����7Q�4�#ǌ{����Ap��]�!{�]�ꞩ�!7ID���7K��ϻ�bx>a ���6����� I�CX��X֭��n�0uˣI�s�Bκ#y�F'dvJ�Z��xD5����L��~�D��j1v<E&���:���?��#��WY�9��!�Wo02Q?�#�F��Q/h{�v��y�E��䓖�<��.�ŀ��pn��3�����f����a�n��41���zc����=���/��Z�]t�������P�}���YI��?�S�F���H�~�d9����^u��̇�qV�ʶt�wrVb���̴���5�
���$?�[��u��N�5�3mѺ�
�ۍI^�����ݸ�0+�P��;��Vs��wS�&�n����[W��_0LKf!JN��b���";�>kts.��������X*}:Z/��R�``��<u.6mȆθ/����Y-i_���.)lu����l�Fz�Gy���Bg$��4"N�O:�2�|X5oO��KZ6X�j
DXWO0��i2�p�T���g��L�V���Phf���s�7����4D{x�����V��Q�tmH������U6`�Z�T�]FGh�#���r��0�V���
��3����Y�,�h�6�|<�~�%@H��7�@KEO�s���EtQ2�9R�)`��E�zԑJ��eHT�Į,3���B�ɳ�J�5)s���xcG�N~��Q21��s@�o˾�V�_2ι�\���
lӶ.�%��gnL"�u�%�ǲ;�.����}�������M����!["�K��i��M�޺�5m}Z�	H�O.���.����#$�c��6�����i̼�,$�C��o��5[��堄�����-~��:~��D����|�Y��U�0��Wʐ*�O�68�E�GZ�i���nP���=�#j;�������f�g�����`A~(籬3��_̾\ a}Z�0�r�S�}�A��L��P��$o�X��hD�j�q�k�����)HZF��,�)r�cN���oz��>�J�|H��ģV��+�֥�|�4��2�^�J@�P�+�\�W[	CA���Nh
��@�R�B>^��.L��/ɠ�1���X%�x)|?�?
GZu|j)�TF����.%�Ga��}�KRZ�
-Pw"s��d�I�W���3m<����@��A�k�Ε�xX�i���xc�~�k�厏H�P;[Ì֐Bˢ�L<�,�q����9�9A�LU������u�l������<'��/�R���Z�x��<���&��e�ѥ��A��lP��/�Qf�s�(U���̮�1��7V�-�\�@C�T%�U�-�3ܼ��G��������mO���L��2�6��O�1����F�}�^�'(�"��%�>?� w��s>���)P��*^5��j4���x.Z�vuq��X���<�;��js�߯逻�B�
��"�!� ���W����UI�`�q vԉ~�NdBJؠ:K��h�)�rv%���m���􂎤9[�w���}}lEj\�䂎X��V���LH��Z���Z$x�z]B�-��Cɖ���6�EV���}��x�#��1AHN(p5�� m��Kfػ7��?�|\�D���B�;�Z����Uُ��k�L��Axݱ	P1GzR�<�����D��Y�.�Ev�Qy� ��*�WA�R&3o�d1���>MGq���,���&$7�2Lu�t��0g%Cl�����<Pǁf(Vq*�J�a��y�����]�{æ����`N�d���/Y^%�E2�<�&�+TX�)IB9/e���{"���
�)�LRN?����oj�K(�b8 ��/۵$,Q���`�W�n��v�_ 8�	���Ey��`Q)l\�W���!	�Z=J���X�)����)��$ �j ��DQB��^ ���طܜ�l����)��$8�ߨ�j|NNfcX�{ރ�ߠgڮ�d쒠"D����JL�ײ��0��=X㢋غ����V�>��W5��ش�����D��e�q,��s���n�<&�.�C�[��_���K����%��!��S4Ѯ���|*R@zCԒ'���ӏ��5�ף��F�ɰ�[��9-R�$�=���ad��c��fz�Y�kZ���S3E�R��^����N/�}Sv��<��l��_!TV�R�ŭj�Ӡ���4�ֵ�{Ǔ��}n��p�`��Bb!�K���R�\��>�Ҕ��}i���EgH��6F�t<�l�o�=N#0n�t=	�!(,�*;+xBE췄� /w>�S�1碼k�`ꎉ8���:�,(�j���T�]k���%��1p���g?�>?_L����eq&��Yc&�u��!������\���O0�j+W��zb�8N�8i��;��]��a3R�pf�M��y��05H�^P�KG1�SQ��`$��|)#��4�1Z��M��[�-��ڂ���I�4�%'��L+B�RR��6F	�fl���r�X��9�{1Hw�E��O�^ר� }oa�hd�7�����-GLT��֖z	Y��%��z�B���2�x�-���/��,���O*��1�g��	V����mu[+��W ��3�-�=6��+��k�	Ǘ �W{��N,([�"�9�_aI�x�l�_���j�����^	�r=
��I�O��Aؘ~��k�MfՐ�L����W�vi��=�JИ3C��o���\n��ڬ��|����:��n�\�b�d���b�<�z�+	��J��C����WS�n[���t�p�j�r#v�%yCl�����ٕKN��G��끨29o1wo�HF%�L�g^t���:^R����s�Tw�<�j�:rl�R^T:�����c�W>��Y�p-ACH���JC|��ܙ0�T�
R�&�>*��w�����K�-O���1�\5ô�p_6�,�i�ԁ�N���
B��*)�l�]_��;Ʀ!�T�;H>6 h8"k�ն�vq�eG�C$�LXǖ���X~���0�'g{G��4�#�����A��]P���"5������5D6m_7�"��\b�~� ����1�����I4�tX���֨��nhO�00�У�����Ε��`d����U�k��5Z-�gE������ֶ�l=���a�Ց�:Z�n�:,��>s��`N���!�)�0�j��pXFGˠ��3{��~�� D��s�<PG�ݴ�0�%l�͜��h����;����� ��]��#�ФL���:�C�]O�b�W����x�.���XtSwԯ|Z~�������:i��E
�o	(�Z t	�r�ఊ�T��k��;����2�������Z�5�,+����v)i^���R�u�'+B����9VN�S��<R�,�n�mӡ�*����LfBJ�:b���=L����Us)��	��ثXEDaZ�xݖG���1��QI6h8���ސG-,!߆_^�Y.�{l��|�b�OFu�y����'�$�*"�/:���|���o�"KU<m����Xt�0P�2���/���INƐ@ u�Ӣ��7h!���5�R7Ц��eD�٪�#j@QZ�Q\��m|t�7���W���8T���G�#�TOrt�0�h��Ս
b:½���Y���h�,��wn0~�x@&�R�~��S�N���Vt��R�4O))�>(E=9'Ԭi���J�� n,W��$�t��{J+��.N���mh�����M�1�.@*J��V(����w�s�ݶ	�b��
@L��{� cm"�����)����²Z���L}��J2"�`�Ǽ��h�κ9HmXX�	��>�_��� 
.?o����c�g�M��q���Vr$����.cِ����NT��0Â�͎K�:7�}��TW���J�iL��E3���GAE�F?�PC�3��nK(^���آ�;����f��ޤ�>�v�J~H"�S@��A\;�aZ@�#r��ش��q���z��;���z��[h*�j1b�F���&���Ī�F��fބ�v�ڃ�So�-�>j��|KN>�_qBVI
��t(�t(.4�?�2p�iJ���><x��T[��Vx|h�.�@auB�/���/֑L��]���,����x�=��Z GՑE��T�)S�P��. ��a��}��m>�
��8"N�d�{DW@��3h鿂5�@�o;�IH!�SZi��x���f9���DP�hVç�����'�,����IK�4`;9�o|U@��W������B<b�/����dZF�A�8�����C:���WA�HP�,.�*m}f)le(����G���j���'��\J�7�O��3y�-���!��/���� J|���G$2���
҅�mzʀ�A}�NΦ(X���_�>p�b 2r3sY�vϤF���RY4S�]�s3��Ѫ�,(��s6����C�J&y���
t�ܟ4���(D�U$���9* |V~ʩ��<��[�@K��%��O�v M�����d_�����x��ݭNl0-�j�~��i�U�S̅��_�Gy�� �k���jx/��z�x�-Ϝ��Y��ќ�V����Ű�_�#+Z���4N!����|�fӂ.�'�ӵ7�GD��&B7�Z�h?�	-��$�@k��R�x���PLۅR����ߞ����_.����tMH�ǧ����W� �&!�dl�T��->uIq�M��>�� ���2'ҙt��Mg�$�Cg�6�Q�P�k(qi	*PC��<��y��;�kȔv����	�`	��/ԡ
� �C<�4J��)�S�I���ec8���M@���
���L�%n?��j-�@(t�� �)7	���4,Q��`D��ivJ^U8S�z��F��=��;PX�l�����7!d�	=S9�s�Hʆ���!c$[�@��3���BL7c n�S�ҳ���w��H)9<C8%̏�e�N����.���m��^����cD0d��"�2]J�&��X�\��6��0�G�7�RKjs���o8:�����M�e��g����i�&@/;���[�+H�K�D�����S��q�P�N���	G��`K�|E�z�t�`�L�Ж�����d�y}q�T�ۊ���=x�Zٜ���g'fu���ۚ�` p3`E����^�}����9��V�v��4����Y?T:�R؉j�5����_�q�&{�k���쏈�3`��7b�~�[X��چx��jn>�u��U����6��g�\N6���twhh�
ѯN�#��jl����,7��*��B OX����w�,S�j���.`��8���:wk��E�Y� o���[ ����촠p<�0��%?��:ҔLŸ�c�&���Y�ԅu��7<�V�i�D�\؇bOˋ�+R(�z^;�8�R�SQo[��8�+an<�p�)���톋�H��߻fβ[�愒`$���|Ŀ��dZ1��{Mx���H ������]��4�%�'��V&=+R��w������n�h�3�Z9Ć�Hh���6^2.3 8��#�;�ר��֨�h]MT-d3֑�	�P!%R�B�]�x��4�$�P}�Du��A�*j��"V&�$t+�v�u6<]"�� +�]�(ĝ6ᢐ���k�����27���,�F��bẒ��3��z���e�a��=��頼��%����cQt�\)����ǚ�-7MA����%�KL�vd�|�G�S��C�y��z�n�K1��i���������L,�	�d�53b%�#zv�м��\��vǋ�u���8A����plr�g%TV��C�t�N��q�V���*���{w���F �f����ܗ%�^M������y<���:�&R9�5�g��c��ز8��p�jyH�!�J� �n!4�kr���Ȃ&�e�Q�����f�Ob{Ns�\p�� Rz6�A>i��ۅ	�CV���v*S�lC_-_�P�;��o��gEH:	| (�7"�z�Ց��q�������G���šX9/T�K�'�+���4FzԌ���^�A&;]Ú�=-�ꔀg��Dq3I7��D��b.�� �p������ =��+�Io�rX��֣�Mn��E0��z�8ū�i��p�r$�LdJ#�Pr U��5�SĂ���tz�ڱ"^�$�r����3�:��0��8��Y�2�M���(!�30h�{��yF����wd{-u���=Φ�{�	qe<��M����'ԋ��a�\GᲔ�D���O�j0��`�D�,�_�F���`��K�]*ƌ�������sl�T��f�^S*���ϵ~��T���w� ���ވ���y�@�t$�rLy����*�տk�b� =�������L~��@���D5mE��0����^�2g�w釸0��+/S��1�-V)kΔ�{%�DSn�gs�d��b	YL�>_JD��br\"�x��tn�s$`��ym�K�<X`+Z%C���L���ٸrN�6c��n.C��"<�L_���.��l�$X���FpG�y`>R��-�$��"D��:m�.|��o�n9KPb^� �X��0��2}���
�큄Ę��]����m��h����Py�7�ƥw�CD�ZA���LQ��:m�"��R�X�K��p�T,V�G�$}#��r�T0W���>�
�Ɯ�e�
Y:;WhL�#�r�"~t(�@��ӳmC%A���)eD��Zt����/l�)��E����Ǩ��[m�zr�,�m��(?��cJ��l� �஗1�D9ޕ�jz1��@�΀�S$V���i������ ����e���eLX�Y��}:�:�D�{�s���2 �������"E����0Ƹ��ƺ��m3v[	�_�F`Җ��.����c�=���3��:{�2;l$1�-�g�����˄��+���3����u��{��O��4��$a��`�Z�,w0E�e�=�����nF�����ȓB�;�����Qfr{f�X�����~���b�����\VE�Z��@r�l���էQ�`��Fw��#E��JshE�j�rp!�S�a��_-MF�|��|G��İ1`�op�a>E�w|�t���^bV�'��4��/�74�2�J�b�ym��%j[�����cJh�� @2�kB4!W��P�?����'�c��2kx�K�u�GP�� ��T�p����.˙ah7�}�G��BT
#?f")}hd��Wۗ 3c�
���F@:��'*���.|�i%%�x��X�a���EW�P��u��j8����,�!��/�>9�1�U��i�,��bM.�cS2<�k�/,���Zw34�MD�#g�[�����BA��PBrm�%f�f���(�����C�'i��행@ F\�D�JjN���-mq��٧Һ�N�Ҧ};�>����B��2f�U����(ޙ��NO}\7	F�(�:��>�Q� �6[st���q��۔܍�4��4�nXH�,o(�w-��}����z���ཛྷ��	��1
]c6ȗz��5'V����U�� �� �C�~�d�W���Kٱ���v�ߴ�cL�9��%����M�h?lK5jR�^�D.jĎ�)�N�2�Bʉ�[��q25xJ�zS�J-��y�;��l��V����p,��Hf�#F8o'dMN��ތA�F�[\f�ia���c��_�Dg�B��wZ�䰜D$G��� kΐ�b��xS�Pg��R(�]2����5�u.����i��O~��HW7��&��Rd��:�8��>
��q9g���q8ݪ+�*2O�t۞g8DOCb�.�q��P=ݳ(��i*�[���y0�҈Sq_��6�j`�99�7{5/O����A<c�a�N�&I���e�����Z"
m�L�^"?�@C�z�j���(/ = �_�}��]�QN<5`����dV�v�|j8�3��g�o��������l�����!��=�Ǳ̎����R�ߟ�$�GBCI��hB��g )������b�ɍ�I�)t�u8���`�sN�!`q˃I�ߖ�ڮ9��a�D��?�� ���'*j<f�s������Z�
�k-�����M��γ��*�>�*XT�:	Yex9O��-�Ďd��&�O���[��8���I�d�hĎ'sÞI���d����|`Nz	ƒ���%�I�[�k���+T�����4��o�����=S�n�ג>���fpu>�!}G�Ͱ3{y���˅^�T$��8�TP�v���C��հrTUԭR�
�jh�m�/P��_={�c��3�шF�`�8�b��6���O���:>�8�ְ�3���! >+g>%�6�ճt�;�̥�N,��*�/���,R��*12(B��h���w�iiS�Í�r<+``v8��:��� A�[XZ��l���a�GX�p�v�̴?�q���LP���<�&��Y��ua)�W^��Ԑ���\�Ofr�+M��z�4%8�wUn�>Ꚑ�ya�F�p�$~��c̆�5�Hq�s��u��HB�_lp$��|_|6��1>KM3#��c���x���83�4F�'!X2Reb��8��@���+��`9��uH������^��3 ��'�>��-CU��������T�aO֌F�	!3%f��x0@�(�����v�������*_e��ݼ�?�����umo]2T Ɔ��#:6<ɵ�|��k5�Ǎ����Y �,9��������������Ţ�ı�$dרp�����͘�1<�����Mc��_���`Nv_)��c�9SC�c��� snp(���F�~]�� ��$<��&�d�
�b�,zQ�:1e�ya��̳��$6?�Y��p1��r�1%/�B�0Ҋ�!�N���Ш�^M�<�we�Fۉ��p��2�S^HXJ�;jj��Ԯ<�vn:h��RF�X���RH�c�u���6�p��sH��$J9�2�IU\��!ި@_�&����x�ՀJ��WnO�j0N�"\�d��S6�v1iZ]5��+���8��*��l~$_3�
;��Y�
goH��� C��"a 2�lGq$� �y�"�B��G�X����fL�']���Ȑ�4�UٌL_>��A���]����XE����w^D��7X_�~Ab�_V O�����e������a�I��X���֞!n�~0��ȣS����@J�Kfw_��d���Ki����5�4>ĝ����v�ڌ���+'�����:����e��tuZ���"���Q!8.�0�ͮjF�?`/�{H$��t������D�U<��A�m�����n�����$_�o~���`��߃�����1�%��t�]�����T$�nZ����!�SE7�C�~i���2j/&�˗�%�K���t?J[r�=N�ZPP�eԿ�)���`�5�]�����Ɔv�P�5H~��kj���P^����}�뽙+J����0nVO�(���ߙ�n��o�l�4���L�ZJ�Y�bM��� ,� �sE����	���X{2GZ�-���a�`��kG6^x����ǐ�B=W��_T1.�d�l&�gĘ��Fk��y�R�GS�$��"��:H��|	w�o a(KK�+�{��X���08��2�rI���L��Zߐv����0���h���k,47ݰR��D,�k�Y�%G�ZQD�my�M�m!����}K�wTg�G9X�#�r*��0����0
Xsý@�Yu��h�I�m2q~���@y�����3�ˡ�L�:xSt"���*�)q�E����0�֯��UK,�:%Z����k�J��>�������x���f13�2@`�o�&�V�?c�O���!�{�T��M��O��L�4���ju���_<���G�h{;�X���D����"��Y�=����ƺ/m��	�X��Ȗ�Hb.����T c�3��CҌ��#�m?$̆��
��F�]�>����܂� ���Vܰ�ϳqګJ��f=��ߕO�{�|��ƋE�����W�iY�nA2��J�N;UԗVfMe����T��f&~�l����͐L�\q�"Z6�	r�t�.�m��0���q��5�O�� �h`��j'����S;��ϊF�zn�:2x�P%�L��o�> �i|��(ԕlzV
�A�<L����4�f2fR�J������j-��[����o�h;�O@M݉B�2?�~���z�C��|���޶ih�xZ!w�U0G�*2��\T��w��0�.��aØ?}L�)�fI
���"7dB@�WvQ�3^�т��@���B9
?��	�i`�0x4�)�\��~Pl����d��#��ݢ-,5�k�J*F�9R�U���G���՜�>�q<��(/���^�Z�@����>7o���ϥ�.�AN%[P�פ� �f߼3(�%�2�������Ȅ{{�u\�Ri�EN��-(@��MԺ%��ҁv�� �<�=Q�2�����ez�Co�v�}7{�De(����3�>&l �gs��Ϛ�	���,���O4����i�y�S���Ô��%�u%l��-+��
߀�1��i
�rp�Ru�PyQ�O�U�;�A�7 G+~�?�u����kuK�������v�p�O�������
�.G9�#PYlf]hj͵�����ɘA��I�=;xⶫd�,΃xe�7z�E�-�m�G<�ΑV�:U���6���#a6�%�N�⻌|����8f�pЙݒ���D+P�B-�Zz��;��Z�k�b&����xZP�c�R��8y@�U�F��6.���*��=5���W�%E&���d�(5�Ӟ>%"q��;�?Ĭ�T*���2��t=$gӃ{C]!��U,P��@(�s�*F�Z��%�yk����cl]m��dS`�9�R�B/ʈ��֪�<P�.��4?I��IS�de�������)}
H�\L�j?T���fj��(�~5 Ե����hQ��t`z���_�.v �?8�ư�ר���j��̬��l-I�0!v={\̩���|5'�>H$������îB@l ��}��u�ݮ����r)�&�8[&�[\pNwA���d����ܮ�\�C�Dfs����J%r����֢�\8�5V~�����m���H�)Ʉ�噧�E0ղ���eS�f�1.Dvَ_�&��	�t:�[��1�A�Z�?�������KN�Dl�ѿ�����
|{�Jz�74����Ԅd�������W*ٰ� ����Ɗ�U=.S�Z��4�fk�:�|>��ֹ�3��a�yӘ^rK��We+��i�v�S���јŐ(�TpC�R]�jCY�j-���{�{_ʎ�3�=`גb}��Ҏ�P7`�-*L>[����@2�;�Jg��6�͸t�.\�@fN�"��%S�R��,m,s*�ebB�t�X��wP/�S|<[��ԧ`,8,��:mH���^���a��.���)���p�;_��?;��L������&��}Yt�u�rOpL�ql�\N��Oy�+H�RzN�8=����e����O�a�pwp7�J�'�AzBH,n��<NQ��:f�$1�&|�X<�$A1k�:M�}��~D\��n��x4L�'�X���Rc��g�������dG���<�9:��HH�:��^蘔 �a��Y����������TccևM	j�%�a^�������ʾO�R��zfW��X;*����C��Zh�l��u�1��` azY�r6���7�vk~!�eH��:Ԕ�,���
��pU���&�����[F��qkx�_���C:ųۥcj���X���̹�|mM�j����h���kvZ�gNv����(C�m�pN�nK%o�Rz�Mǆ��$��Փdd���b� z,�O�u���lы���S��o�pL�9r���%
���k��Ъ�}N���e7�c���)w�"AF��J�*%���^CL���խ���<-�:�x�R��<��xT�퓸c�4²���p^2H�C�J�i2�$�T������&�|��s:����*OXz~)�2\�>�Vu6�ˠi�Q���p7$k�VY*���l�		_�I�;��ߊe��H��s ^.."ܥm�Gj�q_�ۀ�;�=�:��:�X�:�ˁ�I'��s����4�P2������A��]��J�s}��ץ�"�D�y7�%r���b��R 
�<����r��I��*XU�h֙dnyQW0a,��n���_��&g,��Bd�D��F����5���ĸ�p�j��gZ�S���%����:k�T�k�yЏY��C7���(k!s`�0�w���1FXP��{c����ݦ��r��Y<!�;���A��yt���R"��J���Z;Z砯v���C����յ`�4ʱ���d]�U��5���>�ih�?�k��b_S`� ���0~D�0�md��K��pzɀ���GtZ�rB/�5�L̠pf���	��d2�d�GJo��쒂�4j5#ׅѦ�7�G�^���-f2����+e��'��V�R4�cZH�z �n��ǡ�6���2L��=J:zb(����d����sJ �/���kX�YZ8KnD��L�f���*6YH	�$�l�x�{r��_φ�.�i�laE��3KNFf]�y����$�#":�%:#2|D"Vo�s�KF՚��[XC�a0S��2s^���5����9��r�#<�hRlۆ��7�-��Dg�*��üB��Qm��m4а��߯�A|5&^T�΄Gԫ�#zI`r��N0�]�q�
�?6�C�Y��2h�q�h�~*��@4���K�7����R,uZ@t���%�)�ӕEnpG����Q��0��,(��1����J<1_&���K��:t��~�1n��@����vV9�s�_��1%���¶�U�􊴭L����=�3�H�]�zP�i��C�3v�'�������"�,���w帹�κ��"m�J	4r�|�֖��8.P���_�c�Iҿ���],M̨c|$g2C�+#١�]��K���Ղ���^J���A��N�T�E����fX�����"6SE\���f��n<�bo(��	�;*,�����f(o������GS�~h|�q��K��\���Z��~r����i2:���U����ҐX��Doh{8�j���p �׮ȕ��F�<ޕ	���gp�of��>���|� ��0��V�W������4!i�2�8�J����/��6�[�2{�g��h��#@hK�B*dS�Y򔑵`*�.�[�1U�ľ5xCg뫮$GF��֘�T2_Ȭ!�./\a�}�����
�"���d}�(W+3Y��Fď@��]h��r���i�?�x�;��Wa����JP'Q!��~ .�'�,pR30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸���p�&�1�#l����_�)��ToڬrN�'|V�xcĔ�MS�'
�x��� J�恰 *�y��%ّ�'=�F-zӬ���	3��t(�ن��Dq]4X�$��T	3A��"<i7�lӠ�7;Dl�ᣄb� J4��@V�|`'Ñ? �� � ?a���#��7M�r}�ҿr��hd�
�!�t��1�X�r�Jt��i�_yR�O�pԫ3�L<I�
.BV�%�q�at��1)Ct�<9T�Y|����`.��|'���h�l�<!҉�<>�J��<X-����d�<YB�K�ܕ'B_�]� ��&e�^�<ᶏ�j]̩�s��A���s�"]W�<�W��?%��ᦃȯ��hs��I�<iFI�(q��@A����P[�<a4J@�Z¢��a��	V�bHd��^�<�C��L���8����x�Z-C&`�\�<�1�B�n�TC+ֿ -��k�Y�<�C'.�(
#�W�Df�is���~�<����D԰��d�ǭ8�̹SA�֟�Z�Ox�r�}��c>Y��c��;u�޴QDU�^�D�;��]"���'��Qe"�U�'� �O��5�2�� ���Y�x[|1�@Z�l"��ɨM�h:�ʂ�9x�R�+އmu�xz�0D�T!�@   �����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   �  *  ?  N  e&   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�%J�L�TM�P������PČP_`��7ju�r�d�O���<�'�?!�Ov�up��O[��S5E\�]KXl��_�&W,X��wJ�:�͇�/|�a��lP*��<@� 	�'��Ї���X(p�1/jE	��<=Ӧ�*e��O����O��d�<�����'�Z�Q֨	�δ%�"���}!2���'�.�!�ϑ�*����M��rǠᩋ{��{Ӣ�d�<�F���?����P
�m�rbj}k3�P�\.h"� 
��|$���?��`�V ��'�(�#S��'m5�E�qb<r��
�n��x��*��M/ `Fr��㔛p�ay2D^��?Y�����}���z�ŋ_V�
P��4���O��$5�)�S��p��U��EG�`	O:}�:C�	� �ؤ�s,O�c��u�K'2��Yk�ʟ\�'��T�t�mӬ-�ah�O|��H֝�_d��5!V��`r��ռco�����?y0��?1N>q(�剚m� ���'sx��`s	U"@)FOv�"��ֱw��,y��׻�h�H�S�\�I*�a�Mk��I�x�N�?���I�Ov�O��)GY�����M���D1,O�\���N��]�6o\�`���y�a�5��'��ɸ�M��i7�' �����x����*�0z#�d�5O��ħ<!�b�?U��ϟ��	}}뒊/�� P��Z�|\�%����'�j1K��l�y��6]˘�{e�N3frY�>�!
�YX�L`Q
4vO�Q2Q�(Y�~��Ǆ��'�v��S�g�I?PB����$��%���C��NB�.W��	[W�#yѤQ#fϛf|n�'\"=ͧ�ē^�P<�uչVڎ�J��(��u�k�R7��O���O.ʓ�?)���t�"O���!b^�~�@Y����>C��G�#(D�Q��	-@�yrk�
l��Y�#�)���E		��rd� �BYB��Эl��yr@�S�ڐ�u�ϯ-��0�!g� �J,9��?I����'?��p�C���4Eʲ(����0�]+4"Or=���T��vX� ϲE�H���Fz}�U�d�5i���M�g-���M{�Ȁ�2�uC�ǧ
3`<1��Ѹ7�"R����ş�ΧB����2�F+o�Ig���4���Ӏ��Q�4�w
L�8M�]K��'��3iQ�X���*��G�U�fy�b�H6�XL"��*,O���t�'^����mvWH��ЫT%��3��'�	Οȇ剢b�l�)У��0���8VB�/�\,Xff�H�ܭx���,������O�ʓuUp�hg�i�hd���'������0�c%�9{�� 
�'..�� �'6nĸi���� $^(n�#���O��K��L ����[�5�h	�4�^��{fms�o�	h��q�O���(�@	�k
.(�v�8
l��aQ4�xj��?���h��6�C�ui��G9N&�+JJ�*HL ��� ��$S�{ӊ� ��K8�������0�����Ń%=V`�',�r���4j�@����?�E�c��m��?!��蟴֧� ��Y�nQ�&�.��g�(T�`�����A�w��8�AZ�'�\XI�p�ƙx��eJ�q�5� 扁U&(Ѣ��L<���V6�,�2�C�;NP:t�C3�b�'���D�CY��,O�6M�7>`�}���[ � i�I¹T��)�ēV: ��K�I� xcc+���v̦O��Gz��O��\�P���LFʬ�E�R�(��5(9}��U�{��'"ɧ�'����'̄�Whtes��ʋs@��������83�%I�
ZlȆȓ(�X|K@���t`�W*��xPl-��B��e���:�CÊ�aZ���"i����ңv�,����˼ZI���=�����v�ć.Q/�����V�F�r�@I�i�|h�Iy�	П"|�'�L=�B.C2v�Q:�A.���'O��#vO3+�E�cM�=?.eB�'/�$��)�F٤X*�H=1zH�
�'�� *����-�2��-�
 �	�'��i�o��C�6�Jc��aҒ���*[B�'��Ë�i�6@�N�!��F7[U-��E	�"��h����4��I\:�Y�  ��R���!�ΰB䉓x��pzg�$L����/W��B�I,]��@�6��3OM�C�PC��,K5jD��M	�xxs��&l�.��$I�'��]��l�"�x97�F58*C�'0�ʈ�4�����O
�>q����Jw<5�$�
�rąȓ:P̙u�˒7��W�J���ȓ��� f�8mV<"I֥r��ȓl�r��m���9�呸g~���4���s���3�|���e�)��ťODGz��4,��~N���w&ыV�(=B���hR�T�Iݟ�&���(,ID���3�N ae��iH~T�"OHh�3�$jWc��^;J-""O��[�☏���(a\�1iC��y�,@�@cX�	W�R������@�y��W.,d�ƃT����7m��'��#?�1�쟐#�� |�<�%ID���+9�?�J>�S����;_͊Q�O���8�s��	!�d
�]zL{�@.?�FQIьs!�%U�}�A	1�$@�C�ÚD(!��%�\R��>e����Œ���T-}T�T�Էx���gS�"&�ํ��:4Z�>r�4��=���۬�b0��+ա�?A����>��#Ș>Y�9��͚(@M���l�n�<��H�>%��	���/j��89��U�<1�A�$��k0�]2tN�b2!�T�<���	!Y����`�`G��*���S8�� ��Lu9"3�F��z��r���R��G�J=����T��I}r,��>V\!!B�w{�m��G͂�y2-x4���J�>�Ji����'�y��L3Jh<(c0���5!��!���,�y���>O�B��r���~�4 i5ȅ/�y�	
�P).Ȼ�
�-*5�T.��ɫ�HO�ִP���c��Mjwok�ĕ[כ>a#��?)����S��3��� ��WJ�4�7X�NC�3hq�[���#�,\K��ި-��B�	�6��}1��4Y.�-A�(����B�	��JI��a���'(_ \y�B�$sE����gѴ?ҡ��2Q���x����WmbO[$`���iNr@����M���t�D?�d�O>˓,��,)p�	.v�@�2E#<=��D�$}�\WےoX�|���E� <F&��3 Ә\Bh �ȓ k��aP�	V��ɶ�>p�E��J&ꬢD��Kǌq�WI��:&2�5�r<G��l5E����5jG�+"�p��L�4�$�OV��� �ً��@?2�z��&e�-��7"O<H�a�a|q�0iEyH�ʢ"O��yGiX����
-8[�"O¥ ���/��lB���{*r$��'@�<�$,�<o��7i�@pn�����x?��@���$�'�P���ƌ�u6*�ps���Ͱ--D�Pj7E��iR2=!ŝ�q�l����,D��y%�$3h�@0���g`8�`�#8D�D�s�ܽ!�,�x��*Bo��c@7D�h�"�]�,�r�Seϖ*��6�/}R�5�S��=�rU�"
	*$<�A\�/��O��­�O��D<���$-�?E�(A�s��8(�̌�C���y"@��r��\�raV�7�$aK��T��y�
ԻQ��0�DB6:�b���f���yd�,X���F��,W�a�"���y�)Hw���3���!��c'�T���'�."?�"Ǐ؟԰u�ɝ8���*1�E��	2UeN�?	K>9�S����+�P�bŠ�Xv�#�+�
�!���K�.��!�^��[E��$�!�d�;}��Ҥh�/%o�a�d��:.�!��(�~��b�?9���Fh�����+m�x�)�!@�e�^]��������8��d"M��>� �07�
E�5c�?[^�`*��?q��Ӱ>�]'S�%xd��5[��P�X�<ae�Ϊ|Jl���/v`�P��Q�<��F�:i[m����D/hL�WoV�<�������AWu��$-�]8�q��d�q���Sn��4�ƨ�U���p{��	!�����(��a}�l�/�ҀI�)Y�Ȁ����y�DU��"�:ĉ
���1��A��y�,�9_90`�B����e(��y2c����:�KO�8̩U�Y-�y2��t~��+C��,.@�ZP&����
�HO���R%e�Wvt�I�5J���>7�M=�?	����S�%9B#���S���4(� JpB�I�!�V��U�ֶ�n��7JjC�	��FTbNо�Q ��ǂU�PB��`M|�Q����s����C�I1Iz |`�)�d�y1Vo7K�v��P��$�b:�n�CQ&����|�-��͘*��d0���O>˓<����Ik�.��A&�~�V��u�di� �
*X�`x�E�?<����'2^���n	<�
�7.Z�n��ȓT>D���j��O��3kV?X�2i�`�R��	ױa�XY��*-��a�c7�cn��D�t�R��)��Q�bBF��W��W*���O>���ڡ!)J��X*@�`�r/Ǡ`8!��9ª�be�*�nP�$�ǅ'�!�dӣ;!��pF�	!´k�D�44�!�0�����:�:��e�z�x2)<�S
�́��@��F%B���
E�H��c���Gx�O���'U���g��#�슐9�e���;?xB�-�z�臌B�]�����ʒ�f�"B��F�,"���4'���
>A1�C䉂z�,�˵��*��`�d�9��B�I�ws�i:��˱ulv����;j
`�'&#=��@���tA�<�6JƱY¸��FK�D��K3L����O��O�O�B�Jq �xz��Q��8r��a�'�}�Qc�+�d��Imr��*�'n�@y �g� ���%0�b �'�a�5�T�_"谙�c�= �ֱ��'��!�5�D!H��1(��7��Z�{o$�A(����;Dx��K� q���Bj�Y�����?E�,O��1�c���8�nL�i�x�Jc"O� ~���j��u@�Y3$��!9�"O�lr�đ�gnМ8��-p7�E�e"O݈rӴ_v��؃���]3�m s
O���`�2 ��<y§�bgl�)��v�'an�c��I��9���Ce�8�j�;P5��IȟЅ�	B�h���A��D�F�B@�Ԋ-SzC��'ZyfLk�a 4N5h�h�\�C�Ƀ�*�ñd��$*�D��� 7D��2��+*���'5Uc�B!O�UGy�k�/o�*`@��9'{�	���8�~�n߼�O���O
���>�f H�!w��P)Ԩ-��A�x�<�jr��9���"*��8W��G�!���\q&�jRƌ�jN�z�!͆�!�$�?F�&)�ӫ�=mF��$��<Q'!�JN��Ab�Ɗ�D0�4�+|#�jƑ��?�Sf�aC�A���B�6��|xB�.}J^:Il��'pɧ�'hT��	�ҍ5ULl�1*F� ,Rq��!hj!P�ħ7R��"��M�
�����$��l����
� P�A7+ �ȓ��][�`�<�A�*8H6��ȓ{[�l�r��Ljx�4e> ��L�=aE��I��d�o$�zC.��9���S�U0���Id�	�"|�'%�4Ȁ�� "�"�`1,�8v���B�t���>u�|P���3L�`Ȇȓ
���C�M�o bP1�C1':�ȓ:��q�-i�ȅ�Ƙb|�P���IĦߨu�<-0�,)PΡ�b�2�;�pE��-G0Fx捳�� p���!O��p�d�O@��D��T�\]1�N�`�hC��L�)#!�� oJn���&� Mb�<���ߩp�!��$;8)��
(2�x��*B(�!�$N�N5���"		$��H��I���x"�7�<e��Q@f�%V��E�!��=&@z���M�LEx�O�"�'P�I�K��)�VK��uh�m����/Q+�B䉧u����pgB�e(����KHFB�6 �X����(}$��0�cP'I�B䉕?�xe��ˈL����&E��e�B�	J�у�W��ժ%$�/g~J�'Q"=�Rwn�&�y�� �x�!B!��Y��ޯ3���D�O�O�Oy��{�OF��5�2f�5�>�
�'�2y	'��"P1��")Q�Y�'C�#�a7|��"��?j36D�	�'e�����V~�A2҆�c����'
`u���Z#+��	:QdG�S(�a�{B�>�5�����-�t����	��88qƇ d.�}������?E�,O��Jd�+;
��E��^(:쀳"O�4ڄ+J4=���b$L�qo���"O�`���
I&�aq�N�.WhCw"O ʵMI�BR��Yä�0R� ��
O��ƭ�	�`h:N�^��+S���O4}c�-/L��m��^�ȩ�M��s������?i�=���!�Ɇ1a�����t�9��@����a
�ڐ�!��F;��t�ȓN*8��dO�*��)�eE�5͇�� ���d��5C��K�8��-�㉧�(O �*AfΊ��U���7"�)���O�Is��i>Q�	şh�'k����e�K;�x	�ʍnx�
�'�q@n��G"и��M�h���A
�'�(���Mʅ4pX9q�H#m��D��'H��;v뜬*���A���.�@�z�'�*�;�ɝ|+D r"ǚ��D�L�t�������a��Q��*Lf�
ܒ�b�%e�M3���?�H>%?	�o��6.�m(�I�8Z:vy(v-)D�|(ӣ�1dP�My��ئ@�8{dF+D�� ��$C��7�^�a�-���r"O�}Ӡ�K��l�ŉT�S1��ڒ"O.�
R�Ks�� �")�
6>�����d�'�:C�dD�x$!�[�^�o�=$�@F�'�'%��Y�����ޚI�Y�$M���񃡥!D��0�m�+'>Qd��,<�h�c$!D������Y�x8pM� �F����?D���D�C�X�>j4 ɶ@��\Ї.3����-� l���"
5�lC4�M<�Q�,�W�?�'v�p20�ĺ4J��J�a_)z��`��'���''X�B�.�"r�f@���>:����'�����GJgL���#Y�-ؘ���'��u���Z+X!D�ी�V,R)
�'7�		@� �-G��"�B�S.�b	Ǔ|�Q�\���?
(�R�R�N��4�W�'&ԧ�����Ol�2�9B�H�GR@�����;��U+�+0�]8���OL�m�n�g≉"��"H\�eơ�'�P~rNP���*�;"�'����!9�3�P����@+ � YV`��|�=��|~���4�?�'�HO�p��I �LyR"�ߊ�,x0V"O���f'�ē�!ZN��y��>q��i>q��Q}B���c���;֍�
]N4P�]�Q�*�9���	�$��O$P\�`�o���pҁ�8e��)Ә%c�ى%O��|Pt� �'3����5�L��I�V�j�+�F�"	�6�"��Г)�B&�'�0M��K�3|>�#j:h�`�Y� �$�?���hO�b����W�Pnb��5�������.D����Q7h�&HkeQ"C�I�2I-��.�M������'t��O�V���Sl�I6�A6BzdL(ϙ1�T�Ĵ<���?Q�O<L2cK��&u���A�C���w��I�pE�Pn�wk�r��]q8�,�V
��^5 Vl�@�|��܊V��`�C�d�q��:k �xR`��`�	R}�i��3�`��Fg/0�(�� ��#�'a{��I_��X$f�w_H�
�Px2K�/M�����)��gv��#H˗�\����'�剞vb ,{ٴ !��K����'�u����lHі�2�P�)��Ε!H����ONAX�.��0�� ��Z5��Uϙ���tW?�k��'o��d�FÄP����'�L�� ���^�
��e	����|B���J�X�'�	�>\9��S��1<^���O8�}BشY����Į�!��=��D�q��[�d`�mԁyi�zV�F���p8�����䋸X.��@d�'�|Ƞ�I�CF����4~�v�p��?I�m�?9��ƟH�If}�!Q="�̑��G�vhݫ��80>�M"3mP�#���	)K�0b�1�3���*��Pz��RM���(X�\������F<&����X�f���xrkD��>��F)ńE���Ɓ�t�"��%?�!�Cӟ���>	� �A]���R�W�G����t,PA�<�W���D�h`�`��@��e�����'~�I�E��T�m)hi��g+��(���'/,�Z�'1��|J~��)_�!�$�pd��,�����*�X�<�%>Sx���hɰ�6T�<�aɒ;-2��׈0[�時��g�<a��ҘkyVu���]�j���Zi�<A!۶���)%��5���P"��^ܓ"���tB��O�9�(PǮ!��	�6�v�(d@�ɟ�&���)�gy2m�z\��;�f�T�t�҄��y"���P�pi� ?HL�${5<�y�N(J>�RW  <'Α��� �yR��T��Igd<b���� ��Px��*�:, l�6MGl�����r_|`E}�A��h�����A N��,r���5;���B�럀��fX�Pk�㔻��}C[BX�$�<f$!�D�o0q˃틛o`1hFkJ	!�/��8 |�@�@@U'�!�$� kr�L���Ӽ~8DБ��"Z��x��,ʓ#cD`XdT!H@ya �� �Lm�ȓ
�*� @�?D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  5  �  $  )  4  !?  J  �U  _`  �k  �u  �|  7�  �  W�  ��  �  O�  ��  �  s�  ��  g�  ��  /�  ��  ��  !�  b�  ��  ]�   W � � � ]$ D- �3 S6  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9�ӄ1Z���1.*��5�����)z� B�4��E��c��q�B�s�'$Nݫ�%�a���%䀄�r=�
�'�P�1A��BC�a�M�z�l��'��yS�H_���R
\�wz`A�'R����,'3��:��^f���'V�s �^r:�r#�ԓf*%0	�'�6}�Wʈ���¢G(M�Z �I<Q
�6����hGy�؀AK&�z)�ȓj�B��m٩���2a�(
��ȅȓ�]:�L�6�ZA���f#~8�ȓ������#'*XAc��Eb*��ȓ>� q �IH�p9�U1g�Z�Y�)�ȓt$]��_��a{p�ӆ-��E��|�~�w �b���:��k��'��}�ˇA�~���W�@Ġ 遱�yB�L�	��R4�U*P�(7�[/�y�F��M$��W�NK�����y⍄c��#��ChʡE��yb( <�*((��݇py�xI�
�yr�'[�ЙS�/��Wy�U�s��
�y§_&M�y�%, �LϜ��BB��ybk	.^☽0#�/���8����y"A�2Xɛ�,�w�W2�y��Y�+.���d��<,:y�F�O��y2�˪P�$��e"ٙ3Z���U��y�'�4�����$�J�R��S�yr��dq���V�#_�m�fA-�y�L��LY��LI�1ch܋a����y�GV��ac'턖:�x�׃��yR�߫XX�di)\2��tc7����y���[2���E-a�nq�Y��y�%�y��8Dc�WӸ]6뇑�y�凖B&��)tFZ.7n�a���ލ�y�J�.n���I�߼W�Vй�b��y"��Z�,�"3�	K��� ��y��E�*�����P'H�Yw�H �y�	"u]�@�ӚQ�왒6Fݺ�y
� ���6Q�,N�L�c�1LiVฒ"O�1Ue�Ji�m�r�ZU��"OJ�#Eh3�4��I�E���Y�it�"=E�ܴ�਱�c������N�XY����?����*lYS��ɒx�l
1ITv?q�xL�Z��߃�9#q� 3�����If���|%�9:���_�r�$�wl!����r��� ���QR�"�&d!�׃���jf-Y�w�����*.�!�d��O��3Ԅ��z~@��	L��'��|2kS�p�\��g�.;��=�I�:�y@֑,\�����i����FAE��y"Ǌ�a�L�J�i׌^'A�$�ȕ�0=���Mw�xcgmz(����yB�Ļ4Z��%a��`�f:Ը'5ў����[��&4d��� ��6��!��"Or`&'_8)��� m>��ѷ�IkX�� ֋�Fئ�	���l7��5�;D�P�k7���������@�O0B�I@����JQ ^��a�ʙ&yJC�I�C��|giE� ;�m��	%r~�Y��R���1M,C��C$�Y��̅�TD���Aǘ&@��Cb�<Ԩ�ȓ(��D�G��8����Z&H%�F{��T�����HܖsT��r᎛�yR�ܺtWd��AڱZ��������yRf�8^n<YvH�4L�p�6��4�y�DJ�g��EԏC�Lx���H��yZI��Ec��E�U��@w���,C�Ɏ|U��g�/j�@��^S�C�	.@[�S%\�\�� i�B�	;>F��T�S����w 9W��B��	�<�g�$&�����(��B�,�m� 'R3p�re8�ۿWO�B�I�H�
Q��u�xI�4Z�	WbC��6� �ƥي�T]1#�"�B�J�(����1Y(]�G@��i$tB�!$�4���7c�ֹh�FO	{jZB��5
kҹa7�:&��鐒��;vC��<R�44;lK>B�<x7E�<u��B�	?�\�P-I��|h��Q+�hB䉐{�
�[�dZ�ڙ�r>�VB䉣6j����h�܅�"`B�ɴaɈ}��e@v��Er��W	f�TC�	.ac��v��9W�l�)5N��Rk|C�I�V$U��f�t&��ZV�Q�1�FC��<3^��5 9Jc
���*i >C�ɦVr~�y�&�?rr�QZ�ƒ2w�!� �v9���ٰA`@���ѢX�!�d��m��	�O�m/Ľ�0��t|!���	/{�Gj�4��AMU�F_!�d�2nl���m��!�n��5����!��݅�F�X�̂� ̌�1�D�	A!�"y��Cff@	s�~�8���*[�!�D6L�y�<q��4*�ğ�)�!�ԄXT�y�����~�ꡃe�j�!���U�M�#�K�#�V� ���d�!���PFe�Q��Vv���7tZ!�W�Z<TZ`-_�:U�u8ፌ�	O!��1��pCV�@?cS��;Э�}>!�
��)��Eގ����H��!򄜅QQ������e��x�g�R�d�!�ز\v,Y�M�9L��8�'S�\�!�8����#�7��1A�9J�!�� ��X@O��L�f<���әDL���"O�(#"��
$���k�{X�P�C"O�E�P�A0Txp��W
�Fq�m��"Oz��a��`���HG��R`x$"O���W�[�h��d���T�y0�3��'M��'��'��'�b�'s�'C����F��[P�	�}w����'a��'n"�'9��'�2�'B�'o�$yB�jd�	sPWn��s�'�"�'.��'0��'R2�'d��'��I���a�.������^v�)3��'"��'2�'�r�'�b�'|2�',���1��M2U��_%� �'g��'.��'�2�'�2�'��'X�����	Fh�S$��J�1�7�'��'i�'db�'PB�'��'٩����@H��h��]�U%�����'�R�'aB�'z2�'~��'Y�'�p�2�*ʘ9��N܅,I�}R��'��'��'r2�'��' ��'����ǯ��EQ�Aw�q����2�'���'���'r�'QR�'��@H�	�<p��	ߊ`���«�3�B�'���'���'���'vb�'����C������]�w|�lBR�J7B�'�r�'�'���'J��'=��[M�l5R��#Q�&�����u<��'���'~��'���'��'6B�МS󴸋���3P�ȭ���@��'�r�'}r�'��'�7�O�ĉ|�xtQ���}|�2w͐<&�l�'�Z�b>�5țF(ދ�,��D�7G5�q�-�7�yRY�lzߴ��'%���?�
��PA��S!J��9r�cζ�?���MߌU��4���g>i�����S�=���@�
�8m�����-��d��c����ty��=�!ӖAO
ED��� �ɐ?d��OPʓ�?���/o���Z0M��k�̢du� ¡�P�&x,�D�O��`}����)8���<O����܈xW(�y3�;�=�08O��I�?i�?��|B��g	4����4v�E��&		4�͓��$:���g��?�բD-e1�N#7�Ȑ���ҟ��'���?1���y�T�<MC$E+���hOz�b���%?��O�*8��f�'O�(��&�?��ɏVf�C�䄙����Fm�!��$�<��S��yrC�\p��8c��a�D��Ab��@'BD�>q/O1oZP�Ӽ3�YH����'&�,T,VMC���<����?��L@۴��$v>=���gj���\-IL
� �N��6�$�<�'�?I��?a��?!f� T��(�VD@l�}a�&����\]}��'.2�'��O/R#�=vr anƫ�	�r'R�]�.��?y����S�'V�R%�s��\����2X��&���M�Of`1�cڼ�~B�|r]���w��0v�҅�Ӓ"vh|��3�O���'���]3/���%�[�p�8��G� p�҉~�p㟌��Od��O6�d�,�
5+�!"�%�¾Uy�8(��q�
����92˦?�'?I��.i[\ѳ��:üI� �N�V�
�I}����f!��w� �	�Y�u>��� � ɟ���ٟ|ٮO�S��M�J>�ƄW(c8�H��1m�� KFO�����?I��|�4�Ώ�M��O��\(G:l�h�`�M�`����fuҁ�#�O�Y�N>�,O��ĸ�c�N""�'A�	JS"H�w�'Q���՟���ʟ`�OJГ�U 	<�u��nY!I�-R�O1�'���'�ɧ�) C��!˂n�<0iAG��  1f+��a��7-ty�O'�����mwz���f����Fi�^�I��?y��?1�Ş��d�Ѧ�R!��q�d�P�ǊH�zL8��o���'�.7-#�	�����O���(��X��4�&%	�}��Cs�<Qs���M��OP�;4�ϳ��wH�<� �@
``;T\Xo&@H��<�(Ob�����e�MI��7b�U�0@S�N�8�'���'������睉s�BH�
_�_���ز��Dbh����L&�b>5%ĦΓ~ު����E��1�Q���Kz( �>��Q�d���x'�|�'��I>b��T#/.� 8��3d����h}��'�R�'��h ��N���S�,¼��9����S}��'���|�'<EҒ����h�)�P	أ��čR�v�p�b�$?yp�O���><��Rde�: �2� �88����O ���O��d8ڧ�?���!U,�DJmM$thna�ˏ��?��Q����؟ 2۴���y[�D�:�Ϟ97��0٥�ф�y��'���'���*�i=�	?0bvUxџ�%�eh�4�,��G\��5�a�;�$�<ͧ�?!���?����?!���|���F1"��t�����T}�'7"�'��O6r+�:+a�!�s.	�-�|���.	듳?q���S�',0n����S�_�  ic
N)M^q!���M��O6y��M�~�|�V� #��B0_%�1`��)=�^����l��˟���͟�eyRL�>)�oM��˓2�VĩW���#������ �����o}R�''�w�"`�6F��X�ۂ.�%lOF���]�ep���8�f�%���2�	��� f�*�(1<����a�#t�y��3O����O���O(�D�O��?9�f`Y�LH1��n��؂����ӟpa�Oʓ}����|��b�TDXH��,�ơ�ҡ7��'N�]�����Q妵�'��E!(D�4>�1 ƞ �倲�T0�F��	+�'��ʟ��Iϟ��	�
�8�X��9 o0x"�8r4��Ɵܗ'f���?����?�*�l���� tUb����� L`��2��<b�O���9�)"��Չ���P��1\CX�8��L�2;6�h7Eِ%�́/O�i\��?93'7�$N�3�\���8Gn�K�!H�0����O��$�O���ɨ<��i��a1癅RT�<���ލ}Җ���'tb�'��7:�ɉ��$�O��$#�6o��c�D����Ҧ�O�$���7�(?Q����%ן@�W4���#D
\>��퓬J��M���D�O��d�O����O6��|�w�4bB`E����(a2��gg��ey��'��O��e���Dk�&8�W�t����8C'��d�O`�O1�0%�im�&�I?T ���fFMX��fd�f_�	�:Dfhش�O��O<��|R��]$��a��$3l��zQ����V5���?q��?�(O:��'=2�'��R�FY���!|�8��W��O*��'���'��'z �����УG�I8T�����O ��E�׷:�D7̈́L��*oq�d�O����P1�$\��dW�e���vG�O.���OP���O��}r��g�R�1�ɋ�-v��/�^X��a�O����O�|n�]�Ӽۂ�ϵh� �X���%�l=����<�����׹UZ6m,?QГ~+d�I�5(i�R��ǋ]�8���"�Ҩ�H>�-O0�d�O`���O��$�O���G#s������F�.]�@��<a�X�L�'7��	W�s��ܐ��d/r�S�k]� ��'����逌>�nT�t�׉&��䨕��!&ʴ�3�EJ#��/��(��n�O"��M>�.O��1��?�DT��)��F��eVM�O����O
���O�<�a^�t�ɉ�2A�%�ԅS��&��8|\�����M���m�>q���?q�9�n����ք,Wv,�6!�'���EX��M;�Ox���O����t�w]���c�+9çĝB�^(�'0�'r�'e��'�Р5�,5Tx{���}�� &�O`�d�O��'�I,�M+L>��英n"n����]7;��]�d�;���?���|R�Ã��MK�O�)z`��)j��|Å	�`�ip��$ ����YH��O��|���?I��[�6�+#��}��{1�������?�(O|�'@�	ɟܔO��5��C�HS�ĉ&(�ޅ��O�-�'{��?a�E"߃t�(�2h���0A�Y^�}k�O,~�������*��|#�+d��dᦤ)l�p��F��O'r�']2�'E��d_��ݴ(��#���6�͓�"�Y��	Γ�?a�p)�����K}�'b�8��J�V����åűQ�ű#�'�B��78(�v���b�է`����<�b�Ei�N)*�;]�-�3C��<�.O����O����O@��&��U>�h��x)�
���B�4�-�����O����OH���d�ަ�D�q��W�b���Ձ*b�j��Ih�S�'[ Ա�ݴ�yң�p�<3)̈vw�b���yR`I�1�Ƙ�� &�'�������I�s�,�*�/�<��)3*F�3~2E�I����	ʟL�'����?���?y�O��FVđ�CK�^�Hf���'��꓆?����1�	�2���0�i$%������'"	�3��El��+���$����+2�'n.��d눸*�1���C�q%�h;v�'���'���'s�>���h�8�6��.i��'�X�ZA8L��-��ħ<	g�i��O�V,u��hච� Z�x ��W�~�'���'ܚ�0P�i�I4��bP�O�\y��ªt�v@��c�\q��g��ly�O���'���'�2j� �����@(y 0
1d^6��I���$�<����O�|�B��t���-
��)��>y��?�H>�|2W�Ͳ|J�<����6<vr�����D��L٦$�n~"�	"{�x��ɔ]P�'��	��}�a�]!�`�vJ��g���	ܟ(��ԟ��i>E�'b�듛?�ЈT;�:�⭙�ISH�˶�ʋ�?���iP�OV��'��'B�K]F(*�b���0X�'O��Ha�i��	�<KVl�����)!��ܵMs��k�1"؄E��.n�X�I��p�	ݟH�������W&+Z��U����R6"-a&���?���?�dP���쟐B�4��Vx��9
D?
�����k�LqM>���?�'NS0��ڴ����Ix����hG�w^��qC[�r���PBa��~b�|\��������I���#�30Z%��
	�Ȉ��i�4��hy2m�>q��?���	��6��bs�[�{��$��,I��I�����O@�(��?���K�a����d�� !5�����>��d֦]����P?�J>��
{��0(L��[�(�A�?Y��?���?�|2)O�ul�!X>��qR�T�l�^��4�l���Iޟ�	�Ms�bʳ>1�l����j��s�>C$
3Έ����?F�3�M��O���'���RI?� ���H�yD��3,C1+�5(12O���?I���?���?����)�$>�(�hp�Y��	�`�ֳ���'�B�'�2��T�'+�cޝAE�-)Dr�A�� *�)X�O�����IM�)�9���l��<C��'J�p)ٷL=�{u(	�<y��F����1�䓇�4�����L�{�CB�g#��s��:G���Ox���O����ȟ���0�HP���R� �?Q��d!K`��s%�	�	�lg��7C\�J�x����A�x� �O���ppgZ�B�ѰI~�P��O����c�J��gͰ:F���2�H|��$H���?����?�-O>�I�ZàL1�lN*Ic܌{�� �2R�I�����O\���즉�?�;}H�My�D�#S(��z5a
�T\ϓ�?1���?�E��!�M;�OLM��E���d�	+z�9R
�Hަ( ��=^��'��i>M�I��������	SL�A������b��$K�!���'G����O��D�	j{`�����(|1��Y�L�(Su8��'M��'2ɧ�OɊ|9��.kn�1��S�І����/���O���K^'�?�%�-��<q��� N3
��B�U�������?����?I���?�'���H}��'�^��N����D�R�D���Q�'Tx6� ��:����O�ʓ-T>���@�P�.T�e�ٸ ��]HSCB��M+�O <Rw!��/=�����8�vBI�3�aB�ǝ�Y+�d�:O��D�O����O��$�O��?�@A��g�����P4�F!���ʟ�	ϟ���O�I�OUmN�	�U�X��NTK�.i� ��v�vy$���	��S>;���l�H~�a�5��]Ȕ�ɻf�bQ�d��iel]����D?�N>�,O��d�O����O^�#6�E�8~\��s�� .����O���<	"_��I��	]�D�M����V86�r�)D���dKn}��'���|ʟT�h@�O9���{��NL���.4���N_�r]�i>���'�d&�(��R�S*͋�"���a����I蟌�IƟb>q�'�J7�͋M�� q!
� ��A�H\�R��<�b�i��O�A�'�C������kԮn��1���I(��	�>��o�K~�)2`�B��S2M�ɞP�l���ʃy�!��m���{y��'���'���'Sҝ?-
p`��|wR{ ��%z�v��n}��'O��'���y�u���#A��Y����:rZ��@�E +�<���O$�O1�rlY�``����25�L!�Q͚rp`�B���*�牢u��!W�'� ,'�������'J� {%f��yi�	=q�����'"�'�X��H�O����O��$&�v�(%�	f�e��b�<`´����O6��OԓO\�@U`BE�&8�qO��h����Ɠ�DpF�^�l@h��1��*lE��˟����S7j.01�fA*gL����	ʟ�	���	��E��w;(�2s˗�@��I#ǡ>K3�t��'���?���B�f�4Ke�C�C���rЭ�M�L�Y4O8�ĸ<QcW�M��O�ia���beh�x�<`�Ů��K�d�K�I��?4ĒOn˓�?���?����?A�
�����)�
y��� Y�sd$�)O�M�'�2�'����'Ķ�PĂ.i������T�3���>I���?�N>�|���D
<T���&�#^d�A��I�(=��<RB�	a~��Ql]�IB��'n�I,1�9� �
p;u�P���<�	��X�	��i>Ք'�.든?1�A�k��!���:���A"�[�?s�i0�O��'��^��� �_�؂���>�ƴ�KQ�5mZm~��!,ol�S� ��O`woC))]�	V�ԓ>�4�J"����y��'��'���'��	�[*½S�J�o
<�[ǁJ	k����O��$Ew}T��Cٴ��<�8,�4-�H܍R�/N?cC�a�K>Q��?ͧ&3|�iٴ��D &K0�*��ߎ~Q��� kL�.CȌB��/�?�e+���<ͧ�?���?�0뚴<���2)�4f� 4�0�?����$�l}B�'Zr�'��S�T����%QVuc��?Y������ߟ���[�)��2D�9��̘ot	Bc�[�*l-���M��O�)S��~�|RaA�[���0 .DdR�,�c+ ~02�'���'���W���ٴf߰��G�!� C$�ʗ9r��?��t�����\}��'�ܤ��*�X:L�Ab�;Aa��?Y�*�6�k�4����������`y+O���ƎW���"�iCYQ��P?Od��?���?����?�����O�wؖ,�U��"~�*(���$�>����?1���O�$7=�$������QRd�!"�4sN�O\��>��	ՃK8�6�j����� ��*��O+�B(�6�x��"o�%��d �d�<��?1��.?�})Ҧ~��D������?y��?i�����L}��'�'k��e��;tH�<{AH@K�rE����o}b�'��|��K����2[�`��	���1��$�f���(�(P�f�1��� ��c� �䇲\���H��R�Y�̠^���D�Op���OL�D#ڧ�?'cT�W��J0#�%Q���qf���?�qV���IΟp��4���y7"H.A	v��Ѝ�.K
ͫ^�]��'i��'�fL�f��l(ԭZ a���  ��c�U<'�����9}�n�%( �ļ<�'�?9��?!��?)��K;B¨0;��Y������$`}�'��'��O��`�=<6�3���&�D�5�		�*��?�����Ş�U� 䅅A�2hB��Q�N  @�A��M�OD�K��A�~"�|�P���4�Z�)�X=��h�.ɒ�D������	͟��By�>Y��G�	ϕ.G7��`f�PC@T@�J��v�D|}��' �'�.a�wE��GX�q6�N,o��1�R�ql�����I3Ō2K�Q>��/Lu�I+ͩc8T�5'Z�P�������	�������}�'9J�i�$��i����b$��}P�����?��7v�i>�I�M[K>�c@m�L��Խ)r^]�D@	>�䓙?���|�E�ƫ�M�O��d�l�1Z7`�*k��	�Fթ*�$��'J2�H�BY����?�����o]M�ay�h�5鲜�� [�H�	Dybŵ>���?����ɂ$:?�T�#B	_�"ͪ���{���O"�'�b�'tɧ���';��8�h��wѾ�Yp��0i��9)v�H��ܕ*��������1�̓O�x��ޜ��0�ЭJ&�.eP��Oz�$�O����O1�ʓY��H�;iN�0�whԩdm��"g��y��'��x��⟄1�O��$�?g��<���
�!�	ȓ�S�L�r���O�H�~Ӻ�;O��˒����OU�h��,�1#�p�`&��)�&��'���ٟ��	Ɵ@������Iy��!U�.����v/�	�pp;"AO�.2��?���?�H~��V|��w��"W�p���r���'r:̉Cg�'`��|��t@mM��5O�M)q*/	�c�&F$`�ܑ�=O��B�[1�~r�|�]�������PBfZ�S��<�T̝&e0�!I�-��������I^y�>)���?y�l䊥{�b	�נ�A+^��N���rH�>y���?�I>����%?�9�ef�%���� HJ~���Kb 4��e��ΘOk"$�I�NRr���hGΩ C��!Jr
p�'㕏:{��'���'.��s޵Y�'�]�np� ���9���O؟X�O���O��lZC�Ӽ�� �vi2C��aP�R��<��?Q�s�(��4��d/�����'E��y
�C�>�l�G�	sl�h� 9�$�<ͧ�?���?1��?����%�0���k��TɓF�Ĉ���b}r�'��'P����1!�i�F��I���� 
}}��'�|����f�����6���ANҒ��0��i6�˓r��x]�~��|�Z�0��I:7`\1�Aꅃ*gJ�Y�����Iğ��Iݟ��wy���>I�]�8E�"��g�]h��^�#	J���-����J}��''��'��Y1�\ z��aq��(,����"3p��������Ai��+����,x�S��|df%:����nE�g:O���Ov���OF���O�?!JFHY�AXGf�� D��⟤�	ǟ0�O�	�O\�oZR�	67&�z���c$��êӀr�A'����П�j���oZx~��߀Ip6���l��dQ����7��F�>�F�D��䓿�4�n���O`��ɋ"Y�B�
=:~����S%5���d�O�˓W����X�	͟\�OLI1S�
)k�N�a�K�|[����O���'�2��?!rD��TwLi���R1<�ة�U E"G�q��"՗x�F4���I�˟4A�'�軶�'�����NϤ�ܘ��"v[G�'�b�'`2���O-�	=�MۥIP�t� ł"�n̤`�$K��<Q��?�мi��'Q��>���=M� `���G�=H�Đ-6ȵR��?������M�'���&E�f1�#���D'4jv=[�n����%kD*R�w>�D�<y���?���?9���?i,�r�we҈I��Ɋ5�:C���K6�P}�_��Io�'9���w�"4Aq
֛p� <�e�J)3&� �`�'�R�|��dI[�&:O6��WF��B�̛�*�2����?O09�`N<�?q��!�D�<y��?	Z��"@cT�ú�̐���O(���O����<)ES����������$��u��2J6���b_O,Z��?��Y����ڟ�'�����ضP�r� �&L ��$O.?q�F�lV	"f	�1��'nX�D���?Y��`�"T��ʆ�O���Q֡��?��?���?A����O�ՙ�mڗz1�$�ec��X��g�O���'a�I��M��w�`���&�UN�A1c��S<.�(�'���'7"d,ϛ����%�
,�$�C�"�Yh���X�t릊� =�!'�x����'Z��'���'�~��jɘGg��£�ܫ��7\�X��O����OT��,���O6p!�i2{+:���Ō�!l6d�s��V}��'&2�|��$*f(�0p(/�� �U�!$Lh j&�i��	�#���1�O�O�ʓu����Q�	��EAч�3�x1����?y���?q��|
+O�4�'�r��0 �c�$�(�J�vaV>�y2�bӐ��Ox���O
���y2��zAh��2(`u�Y�<���t�`�f������J�L~���j0��K��0<���A �!�L��?)���?���?�����O�M�`��\�SmB�+��C�P�p�	����?�R�4��s1��c�.�u��%C�R=��<�����D�H 6-=?�0�s�? VX��C7�4��e� �4��5�?i1i*�$�<���?���?qQAw�����_tȘKw���?I�����U}��'n"�'��S~��Q�81J�[� �\�P�nv������	`�)��/	��Qv�܏+Sf1r�;Z��p3m��C��-���G����[d�|��1������V86��I��%Ȳt���'�"�'d���\� kݴmLiu��( ��y`A�W�����?��]������y}��'eva��
:9"Hx"d+��@V�'0b�=�6��Ĩb��q�$0GP��0�{&.��qH�"0<O��?��?i��?�����iH7{Bщ�	(���"���'T��'�b����'�6=�� �+:XLjWJSNF� U��O���$����Q�6-t�03d��<&m ��3�\Q",v��c��!u�˅P�Iiy�O��`�R��4��Ԧ4p$��H�R?��'`�'F�ɦ��D�O��d�Ot���$(Y�L"���?
^0�$�7�I$��$�O �d=�����yST�IgƉ��*V����΀c�O5T �c>�kG�'*�5�	�� k��H|�dU�'���l����������h��O�O��H0]Npa��,K�ֽ�&N�(H��g�>�.OBm�_�Ӽ���]�Z<%['�"����<����?a�$!�U0ٴ��ą�lŬa��'s�J��K^8e��\��F��y_�d�ŀ$�$�<ͧ�?)��?���?qė�	��X�e��� -�f�ؿ��Z}��'���'z񟮽�6+��
aV�h�bWx�
8��(MZ}��'�Ґ|����V�i���v�4t64�`q����S�id���s�Z8p�O�Oʓ�����5R�J��fwX1����?q��?!��|�(OBA�'�+�)SN���+Ɵ�X��3�['D��/q�v�y�OF�d�Or�$I \T��Ja ����S��ܴc�R�w�d�s�%���?a%?)���)��l���η�T�`�薑	������Iş���ޟȗ��OCع@$m��O:����^�Z�^,��'��'����|��BG��|�,Bk�(�8B1j�Q��K��'*������۪yt�星0�0��=��r3Ȓ-h&Ȫ ؿM��x�C�On�O���|b��?)�	FH2���k�J� �C]+(�f[��?�/O¤�'Z�	�D�O�d< �◘�rH1��ȕb���Ol��'@��'.ɧ�I�2V��i3��T�y���Sud��7�p)��W�'��%�Ǘ���+<J2��\�	�
^<3�RA��ˢ�ٰh.nT�	ʟ���㟐�)�Sjyүd�����z$iBcS�1W�Q�3O`���OR�l�Z��K!�Iğ !EG�/ ��ٲ�B�g���ʟ��I�w��mZ~~��:l�|�����t3m��B9=���ɓ�4���Wy�'���'w��')�_>��GE�:n�ӁJܖ[���cM����O���On����Dܦ睺r�q!JbI���ÃO�,q���	���%�b>�2�Φ���b�:��'ƀla�*ߞa��=��X �r���(&�l�'���'��d05��	
�rJR	�I���'FR�'�BY��)�O ���OL��ؐ�EN'����3>��ģ�O��D'�ɷ+�%�u`�&tz�����%5�M� 
�F�9'K`�L~R���Oj���xxx�g��8Op�j�OY3'ٚj���?���?���h���$���|e�e�F�q��`��2lT���PZ}"�'r�w���]�\�u���'�z��ѮX""}z�I矀��۟��jB����uw�X'#z�䡛�O�L$:�Y�@T(=S!H1rl,&�,�'���'���'���'��i���S!rV��b��J�P��j�[��i�O��D�O
�D*�S�h��(҆��+�D�S T<kQh̻�Od�$�O�O1�܌t�II��kr �gTH��TN�]�.6��hyR*\�r�j�������Q�{���i׫��H�� �pn������Oh���OD�4�vʓ0�I�����<���+&ƥS��
ŧ��8�۴��'0�꓋?�)O:��w@#l,���"��3"��5&"6N�6�4?JјK������'ϿC���	z��ӇiL	��(�J�<����?���?����?��tkT?��uP��B��P`�$�]����lèO�I�OHl�t�#[H��j�[ne���iOm��&���I՟擙w�ʵm�t~�Ȗ�m��|��B��5Le`Bh0ў���
W?iJ>�-O��O����OL�Z���+"f`��#\
���.�O:���<��T�|�	ɟ4�	`�#��>�^�qC$4ݠ�I���D�F}��'�"�|ʟ�0�`+�?h�P�[�j��c9@	����%��	�f��`�i>���'�:(&��k�*�F#h��;ixbb�������I�b>�'�:7M�<o��$�^�*�������<�i�O<��'B�(
>f�T��
ݶJ��. #Nn�ɶI�>l]~�˨.�����`��	�a���HκKk�(��#L��~y��'r�'���'��W>yZ��&J%Tiu,ͩ0���%$˫����OH�$�O2��J�d���|���!��(���0` ��K�������&�b>m�Ц	�S�? �h(���5(��@�C���L�?O�1��b��?!�/(�$�<ͧ�?���[)> ��_�Ti�3E���?����?����YF}R�'_B�'?v9�eZ,
�r$m1K8�H���P^}��';�O@�A�P�x�
���۝�a�P��`�,�uV8� !�Q�pR!�ß��uĉK�$��%��"UxT�
RhDȟ��I͟L�I���E���'�u*�HIw�:f�Ӕ�t��'����?��Q����4��1�
3\��(K5I���077O����O�iD"�@�i�i�4#_����j�5=Z��KA�W8���ݳ|��X'�����'v��'���'}6�)F-
�vK�,ta˂$���U��)�O����O���)���O `�eF�S���GY8pBHE�"�E@}B�'�|����ύP�8A����o���`ĊʮgNa�&�����G'ژ��'ܰ�O�ʓ��(�b%��R����B�<x0���?����?��|B*O�u�'%�*��|ּ�[�\,򲥉�M��2X��D�W}��'[��'x �R��[+�P����RĨLJ�F� C��&���2,���t�I���Yנ� = .�1-�q�e4O����O*�D�O���OH�?%��OD�= ���a�&*X�Gß�I۟�B�O�l7���|��v�2�e��b� `Ь��''\�z�(�����'NN�a��������D�B�6��k��q%���\H��|RU�$������	ݟ�Z��(�έQ�i�fA�B�����	OyN�>���?y�����A��t+L[�T� 
�lt�ɷ���Oz��S��L��L�4\����B��q�͗z�9���:�P�x�S�_E@P�I"@��l�C�tv^Q�Oݦuʮp�	ПD�� �)��Dy�v�yd� ���B��&D��T6O����O�pl�Z��s����k�털(5V�ّ�u�|d�Ռ�ߟ����y��m�b~ZwoV����O�|D�'C� #wنX���#���H�'���؟���ٟ��	ϟ���p�T��Jl������O~�Y����j^듞?i��?!I~�aJ��w=THa�h�z�ء� �@D�� ���'.��|��$�i՛�0O�r��Q�]�Hؠ!Px�|�=O��%��?Q��(��<ͧ�?����VQʠC�>���A��˪�?���?A���N}��'���'����c+ t�&BbT  R��D�E}�'��|����(C5�ފesL�;uL��$Ƚ8�P`W蕄�H��zh)������M�H^88��Ԫ��}Yb&;1�����O���O���)�'�?��/Y�̠�B@��EE�<u]*��� ����O��ě��?�;:��]��˦�ڙۄ#
�����?)���?�`ҡ�M�O�n
	���I޵],�:��!|
�QL�!6>�I�O>I-O����O�D�O���O��"�㏣e��\3¬:Q��SpL�<Ir^���Iݟ���_�ݟX�r�O��>��+�%̭{Q�����O��d<��i��3����L*X:v1�R���uԽ6 r�4�ʊ8�n���%���'3D�£�>�$MF��}������'f��'^���DR���On�KY�������� Z�n��m�I��M��2�>)����$�)�>��" I:_�|��L�gr��!�n�l�}H�mQ*៪H~Z��?�T�؆|Ռ��fʁ06zB���?Q���?����?�����OJ:$�ebֿgE��{Qc�_�؀i��'%��'F�S���z��O4uI�#Z2PZ���1;�P�����OP�	����4��dS�??�:�@C�x�\Q �� \�ȑq�A�*�?��.#�į<���?����?�SJB�\�֔�T*3���J�?�����$g}R�'T��'��S�ew�h�F�2j��ȇ���Ơ�;
���	F�)�N,~��`\�Jk��:%���p��"Bk��M�]�擔Z��2����&ls$�$?�4yq*�<Jx�d�O.���O���ɺ<�c�i~����2ul���L�:��,
�'���'4�6�6��"����OZ������+`F�	��Hڕ�楹<��O�
�M;�O��&��1��<GoL�#T~����G�,@�Ti���<!*O��d�O��D�O0���O��'n|� ���hT�S@˝�ͮy�U�H�	��	O�SLZ����gG֓qq�x�t�FjбB"����?���S�'h��T;�4�y�,H*���H���!9�>�S�e���y�
^�T���s��\ 9*:})�k�<�)ƯH;��ur�#ђ�> API.��� ����Ā��T?y�� �H�	:3�i�b�~��т�C�@���@�	6�>O8��E�S�����C�!�}��Z��R �K�Oy��TiϨ7nQa4�$䐄T&K�K��<�a�EdL��M׌f�9��1!����GW'�\}���M�	.��"�e�q��AJؒC�4x �
+8In�{B\�E�b�1�-ʠt�r�h���)3jٯp���H��!_��pqfFZ�"���g�Ó[:�hӎ���O�u��-G6Js����	��I�������	H��������.)�I2��K/ӛ6P(2�[�)�L7��O���<����i�O�d�O$���	/\H��ٳ�߆}b�93bm[e���D�	v�v�IR�~be# 1)�ԉ��bR�k$� [����'�ny�~���O��d�OR ק5���0�bT�̟$��i�V���M��?1�R)��'q�� 6�����>�"G� :&>]3��i���h���O��D�ON��';�ɴ8[�j����l�@�9t�g
�+شP�������O�5{����*�ReqKN���iJ� �Ȧ�I���I՟ 	�OP��?Y�'����"�(y�8pH�NL�2�qX�}���Y�',2�'+B��/]P�C��/u�X!�-�o��7��Ob�$�K}r_����J�i�M�G���6tH�(���(�>9���8�?I-O��$�O��5�4��8M�<��Ʋ6�DJt��/�M� W�8�'>2�|�'?��ֱ�.q�glʜN�P����]'$�a�|��'B�'��O�"��n�$��+�.@�����FN6DZ7�<)����?!��f��'�<e�'���)�/s;�Y��g�	����O0���ONX&>Y)��F��RF\�RF�x�Z� f$^�&n��D$�H����!�lɟ��O��P�Ѭ"��#�"��D�>)E�i9�'����3�����O$�Ӽi�ڑɢK�x:�2(��l@O���OH��r�9��[:w�R�.=(tx�`�pB�8"�a¦Y�'��qӖ�D�O*�d�ON8֧5&A	�vC��#��	�y�6��h�M+���?ѧ��'q�\}
��N�QL�-e���X��M��6���'h��'Bʡ>i+O =q�E�-���7�Nm�Z�12k�Ʀ����U}����OS2��6w�b誢�T�t�Н��Ŋ(N�<7-�O��D�O��$Kg}�\�d��^?�1��L�����+R��H�6�Z�	L*�HM>����?��C��ӍA!�;F�C���)H�it"�'/NO�K�ɝnX����fĒ����ɘ\��̀K<Q�����O����O��O�\咗���O�T��C,� S�!۴(�'��'R�'�i��P� �H1���`y���h�R�ĸ<���?����'ID���(��9gŞ\� l�H��lZ�I�����g�	xy�O��G�?ڶ�ר�T�� ��Nq�O��D�<�.O4�'�?I�MZ��A0aS�Pf`�V?ߛV���O��/���&�p�P�/$ hK�DY,N�[�x�F�D�<�(O(ʧ�?���?�1l��'��u`<� EA�>�&����By��z�O뎂>�UW��P��-_�'��'�����ɟ(�	����u7cYCs����� ��Y"��*�M����$�63j���	)�Hd�[� c����W�t����p�	ϟ��	gyʟ��+�	�H�a9�&�0��0A,PX}����O>�a��\g}���Sn�|U*:�N��M{��?��?�.O�Sa���PfRݻ厔2)S2�HWO�@�lEx��'�S������h�'�{&���Ƅ��N5��lZ���	ryl�~���M�/xZ�HU��p�,��z4O�����������	N��Śx&�8���:�ARA'ހf���$���O�d�O�ʓ�?i�Op��Ң�
Ѩ�ÕǍ�2�&؉۴�?1(O&���O�����?QG��+ [J!�T�2v��*n2���'@�$�O�˓�rUl�	�ε���
����E-HN�듖?���?y���T�1��9�Z|h@gƧ-�H���Ѕmt.�nZ۟�$�X�����'��hu��1a�I2�:I��1m�`��syR�'l��:���Ok,\2a&�#dN �T�v��V��_�'��I��k�s�֝�w�Z�3�F�[D������&G^7��<��	��6�'�"�'���>��\�<D�p��\h��!��C(dO
�n�ǟ��I�N��ICy�'[q�����E��zU��b!��he�p���i���j�2�$�O���O��	�O^���O}I#GR5	�@�@;�A�͛Ϧ���@ٟ ��ay�Oe�O�r*�7/T�y��X��x��2JL6��O"�d�O��DVɦ��������ϟ��i�]�G�5 ~x��b�,${�U�Bp���?%�C�<�O�'�R��#x��rI��k�@PL"1�6��O��d|}�Z�X�	`y���5ƫ >/g8I�dH�w�$ٚr����d�9S�D�<	��?�����/B�R����
��=~'�%��iT듄��O��?���?y4�͝E�q7�����ua�\3#�1͓�?����?q���?Q/O���|�Q�ҧ>���6LY�=N�P�Ǎ��q�'�2U�t������I�yjx�':�޸Z�ˮjD�`3Ǒ� dl�۟���ڟT��Ly�O�X�'�?�1%�(�ChK�6�~53uK�)n��oZş �'���'2O��仟3v�PcBKO�{Bdѡ��N�gz�7�OR�d�<����ҟ���ȟ\��'�G���ǯa��t������O|��Oj���=O��O~��fi�Ebc�����qP���7�<�eg���'`r�'�"��>��3��ɕ抸QT|��AH"��Ho�ӟX�Ih4�	[�Io�'N����� �������i��4o�ҟ���4�?���?Y�~�IEy�DF��6C�*C��4�B7k�!y�7-�(%��\���h�;b��4x�p���EK�k&!D�i\��';r�'|������O���=`r���	#`q���1J�&k�7-�O���O<���2O�ҟ���֟��� P�CF��{ �#WXvLb�i�r�'xx�����O�ʓ�?�1):N�˴�!���G�'���nZ�pB
h�h��՟x�������F�\ce"�*$M,"5�P
�y� �ߴ/���';r�'��İ~".OL��ݵc�|]�R E;�Ȑ.�>O!
��>OZ�d�Op���O���Oʧvś��Z�b���ĨS95R�M �-�y[N7m�O
�d�O��D�Ox��?��B]�|�.���P���0���`d��8@��F�'�B�'��1�Z�5��⟸����)�����i�#'�ݡFN��M+���?q����O��<��'�!�W�q# ����a�hр޴�?�������O\��OJ��'nb�Ԛ�4$`&lN2`s����(R�I���?���?Y!E�P~W�(�'q�q�c��<~�9)��K�z��mby2�'�7��O ���O&�Ka}Zw�Z`��V+6�4y��"�'9Nt��۴�?a�;���Yz�s�t�}:�B�$���A�O�/ajr��1�@ۦ��	*�M���?!��?�rV��'+�ɈPjQ/���c@�W�!��F�l��6�U����<1���'�:��T�}�"�C�������M��M��?���?�#T� �'qb�Of�IQ*p>x�UW�|��3�i.�'����i�Od���OP����)Ov��e��gn��ԀӦ���ş�x�O�ʓ�?!)O���� 9E�Ьp���P	?��aRV��@c+?q���?����?�)O�N���D� ([LYx$Sz����>�*O����<���?1���ܹ�q�ÕO�:+G  ~F��\~B�'���'�Y�擅��d�C?��}�ԦV�,o��*c��M+O��$�<��?���Yא�ϓ3~�� �`F)x����ïAZ2@[��i���'���'��i>]I����d]D�8)�؇Pl�`��bz�\�d�<����?y�7�4��>Q��Y�kf�� ʊ(�0�� ��Ǧ��I�@�'r¹~����?9��o� A(�)��7���SQ��+>q���TS����ʟ����KvT���ĳ?=���opЕ�_n��PC�f�\ʓ�?Y0�i�R�'q2�'���Ӻ۵bZ+5!0h��J83�8�j�KĦI�IƟ�H);?�.O��>i��H�Y��-hC���M���dtӮ�d���a�Iş����,�O:�kE��fbI�B<���ʍ8]�|��G�i"|dӞ's�'������N)" � ��9����L�D�mП��I՟�������<a���~"%��Q:<�$x�x �4i	�Sw")mZ󟌗'��J�����O���O���kR�B�l9�@�E��*0��m�䟼�ɮ��$�<q����Ok�>d[�E��ٴW�(`&��	-�ɗݤ�I�D�I��h�����u׬az���3���9��$��M\���'+2Y����韨�	!z�auI[�d&D���J$ܾ��c�p���	�����؟ �	Ny�O���++������w(9�T�V�3q�6-�<�����O��D�O���6O�	x���"�:5(
{}�����%�	ҟ���蟸����k/񩁴PQ|�cA�=,SFP� m��m���L'������X(�G�ȟ�O-�g�v1�2ȕ+r��,; �i��'V�����K|*��?��<"������U�Ȃ�	�#d�'%�'0�`��Ĩ?��ŋ�#e)��f��u��j�z˓�?ّ�iL��'�?���a��	�r53G�ֵ/��7"\4$�0|oZğ�I�����G��cܧi�\��˕�[����U!��F��]o���i�4�?����?!�F�'�R�
%9\Ir�/��Ra�b8||\7mGQ��*��+�Sޟ qt�ĶY��PX3�J�3� ��M����?Q���?aD�x��'���Oh��\�0:���"d�p��i��'��T���'��ݟ���ҟ�6��S�AE�
X�y�C`19+6M�O��p��?�M>��G�jPr6��v�����0\���'�x�S��'�	̟p��؟h��29��:�4}"��qL�Qې�iNdO��D�O��O��d�O�`҂IRn8����Τ/@� ���ӕP�&��<Y���?�����':T��"< ۢ�3V` HDc F�	ן4��d�Iן0��$�"����R$!֠��#S���b�\.s��2�O(���OH��y�S��ħ&�����&�+U�iI�CT g0��i|��|�'}2*�y>���� #i�E��` "�<a�C�æi�I��'�� ���O8��� ���X`��
=�	c!�`�'���Iʟ8�e����%���'c���B�FN�Q�f�����s��ho�YyR�'�6�v��'�r�!?�B�_�h�Y��Ia���gHG������������$�b?��0��I��5�����jcr�J�ĚզM�����I񟸨�}B���?\(D(։{_���7n��L�۴D���2������O���=L� �c���&'G��B%����7��O4�d�OD�d�~�џ��J?�ŕ4J�P �J�8@��W|�#0j��M>��?���W�`Aa�e	�j���pBD�#�	Z%�iMR�'�HO�:�o��e�˔��Œu�Z�Rl�%����}~�-Ԩ-Vs�?}�V)0a�Y�u��0�w�L�%q�)�DiȯQ4X��	�cs�$:Ӆ�B���
�Ā%���Z��G�	) I��oŵ:9��0��_��%��!���G"�"<8�ݣB+Z@���� L�t0Z}"CB�: ��q��P/?h�P�E��A9�O�g�� ����ԥ`�:�C�R�{����-��w9d��(δ ¥js� �*I�T�ۻ\�����_�8d0�r(��[a"5��V%^Ȃ��M�#�s��Q4.^D1�̷}�0�"�eů:O4����ۿ2�p���/6W���#�ު"�%�AJ�V)��X���R�_�<	��?1�m�$%e�
�+�	'��>�O��˝&:��K�iT$N�,`y���ȍ-�ά#�� [bP�}�EL�T��)�*%sr�b�
C�'��0���?��t��0h��@&U
MC�D�6���y��'۴�HG�	)��0jӎ]�&���/d�'N��[@�ʆ}�  �4L>�R�И'�z�$�>������?���?1i\�ar��:P4���j� ;��#�.@�|�*VV+�*��c>���e�v� ��^���Yє�ZP!�OJG(6�ZaK�{0r��)�� �� 4qQ��qb� 1�ʕ�WC��SH��I՟��䧃�k:�����68e�ķ\vД��Z�:)rЩ_�=�-�d�߶$� HDxb+#�S�4N���<���w�N���N�9�R�'�0��f�t���d�O����<A���?�cX_����@�\3V�¸��ng?1�c[���SdD�A��x���'�UJ��0x��������~�M_�KZA��	P�<P��P�#T,1'��.���aߣ���I9a���'�ў$�'kV�'6g 	5�%|m���
�'�L�a�k��LHl3O�r*�!�$;�S�U�`�˝,�M�E�9p�����ݢJT��a!����(�I��'���'����X^��MУT�v�	�Ɣ
XH�hU<X@�\p�JC؞��D,ŏ<Μ�h�b�-kQ�
'l�v�-��j�tntd���^��	�%
u��0sA�k��K�L	b�'�џT��@Tj���C1�B���$D�̢�H�0j�&麔��)��1K%jp��X�O~˓	��h�Z���Iy��E�Q��������³�yb�'@2�'P��
c�Ȍh�р��T}*�t=��,��U�R�11�(���g剋$Ҧ�����E��@8��4�^�K�p�(2*��A�����(O��D�'y"����S�D����֮+:�	X�6O���$E) 긡!e[�S!4��g�J�a|R�:��	F�l�nѡX2ի�B��l�D��l�����h�埸�������N(l�a��+��V�����k�=T�(4�eLQ��ē��)+�9OFuq�E�7+�J'��M*0 ec�N4ȑ����;D^TA��n�"~�I�?#B	�bd�?	B&�����?�:��#"�����i��&�';?�䊕��-A�T��T�E�6��O�˓��<�G���nB��(?lQRL#�ÆJ�'ě�`Ӿ�}B��J}��k�!Q�0��2S�B=�?���ȶ�1�ij��'��S��ɟ�z���=80�c�(����i�f~�����,L��t#�K3LO����1/g`�q �1���;&oR�*����&V3f��"i��P�����4b��r���]1ഁr�«D_]rv���4�N˟\�ɰ�M�gy"�'�剓�lIZ�*F7"�&ಥ��1R2�C�	�t���#+�>�ta�N�vX"�Q�4�?)H>�,��ʓ
��̻�������pj8l�%��t��)���?�����4���v>��@�=zY�LZa U|�V�pt$9PS�;��|�E�:]�L��4[
e6!pal�;krD���ݠVnJ��	v�����O��Q �(U�b`I� ڀ���i� �O���<)�������L��	�/�&�ޭ`�IU:	�!�d	Q��H�ޢ�.���G_�k��D������Ey2����7��OR���|:�.��WJP�2��cwH,Z�.I�<!��?9��M�L���Ҙ��g�0�"��t	�$M4J�Q�\�G4��.s$���h�"��)V�1�a�:��e�Ig�OxX��Z%�|�ah�i#~ �	�'tq¤�G<u��P��
4�z���bX�'0�i�@㑼>G�@����(y0�'�jL�b�o�@���O���B���O����a��u#FU n!X���7#>�au��O`b��g�'j�HQ�?&*8�1)8R*�2�A��"Q�"~��68 �Il^Id 
�C���
h�cZ؟��<E���%�����=f�� �@a܂���'�:���կ@�{��/Fm�h;��DR`���)�)2x����
��uhz����0v�v�D�ON @Q��Ц]�I�D��Myb��y�'=����� �
|����{4�U⒉؈6e|4PK-�h���O���<١/[��� �tNU<y.�P�OH�9�p���|��E�Č�k�\��'aQ�(�vb�����	���R0t��"��x@��O��&���.'�&���O��*��Os?��S�? ц�OhZ�� d6n>8��Sg���	�<i.��<��`��8-
�㚢+���3DC��?���?9*Of�$�O��S+0�D�OJ�I� !_������9cY�5�'�'�T�p-O����?��q�� �+H,��J��'�"�����?��W�	����� 	����-�:�?������O���'_W�$����=9`�������ȓ\��{f��i��sE�Ip�=�����'��I�"s����	柬�O}����cށd͊�:��t��[�'7r�'Bf֤Cb�T>-[�(Ps5�}[
\�Q�\x�C�(��T�F�Ƈ����ִ�б��"	R��Ē!%d��.5%��V����"��8,҄B�ɻ W��cG�m�V��S��kZ\���Kc�	 ��(��ڊH�0p��C�
06�I�PxЩ�ܴ�?����'�?	���TQ4X���w�\�9�R�JЧ��R������������7�@�K��ȈI��U�׃��6}˓��e����e^8~�����~��԰��B1DQ���'�1O?��F
}8�9��/2�����E|!�ď~/�@*Uf�&x�V1@����k��Hj���?!��t"���DX���5�6D�(�i�09`��P��5z�-�4D�@�VȌ7=(X��	�/4�.]��-1D�jA�*\��Qcu���_���.D�XwN�x
D������i�c9D�<'k��I���TDJ�Y!��/9D��Y"�x�� 9у]����[u�*D�I����Dy���ș*���S#D�4�S���*e�rgX�6������ D�d���a<��h�K\"�,��s�3D���)�;})��8ǆ�'\$��-2D��!7���d<���+)+(Tc��2D��:28v�2�K_2��h-D���v��tO�4qW`�6>BX5�M*D����l�'��(a�ܷ9�\��0�=D����lǫI���� h�X���:D��)& -\B�!�kU�r\�p�:D�43����cU"��qhX{�J�1�G:D�tӅo�.B�p�`��k�.�Q�@5D�y�У|� ���݈D�@��1D�@�0䎌qA&��SN[�zd�O"D�`��K@��r�0�L[)9$����i:D��ת@$lL�i4/Y�u�H5�:D�ph0�#���!���5K(���b:D��J����XՒ�C�8s��!�j6D� �� ��&-�%@`��W7���$1D�D���"u��9��_�$8�|{w�-D���Pi��2�5yQ�ݑB>uia*D�ԓ�E��6|ꃨ>Ts
��qD)D��sT��%$�F�����@���M%D���YexBd�$�@������#D�x9���f�,prc��e�
�x4�4D�|�._
�t����� �oc�<�C%)~`𐑡�TI�v��'��V�<�2�	9�m=�0&Km�ʀj��V�<ad慍Y�0�Р������U�<i�̒0(�J�	�369�����RK�<QR,�XODx��E�O���P�GND�<���,|��X2�4�!#1b�y�<����r��� EQQq��*��^�<9�JT�3��)��K�(9l��LZ�<��T�w�"��M�'�h|���Fn�<郮L�%��b��<fE�Qp$�k�<��3��b7h�!�$P`���g�<y�'C$t�`�C�EH�"DjT���d�<!��Nl��@T#*H`z&�`�<� �pc�ڴ8E8���ET�`2�\��"OZ���d&��ݨEK�F0���R"O�q�E�֥�@o�p*�ܹt�'�#�	)������X�fT��	v��$wAC�IT��Q����N�����j�3?C�'�nQcsI�|�S��5s����	C�ִ��mV�Cl����~t4�D�ܹ[�4�P� M=ZP,�=�) ��@�TH���E�.�D �DM� ��$N( O�9R��,	P]+`m�!On� bpĞ!�x"	_;&<�kǬ�/y�xP�M��<�W�X[�1Ox-�� ُ5<Ҙ.˸Q���"O&� ��;W�^؊��
���"O4�%�J�J��(نl��:�D"O�H����ZӺ��pl �]I�qZ%"OЅ1a�C�*Ĳd����^f���"O�i P;p�r�1#�M�Je���"O��f�3?案g`X?TR@� "OJ��a��-f bjáěTL��1"Oa10a�*8j� y� �A�(ʥ"Oj�xF��
�H�5.������"O���ҫ#<�h��O?���ۥ"O4u��.�z����K_{ܠ�"O���ICm�"$�M�\���C�"O*tB!�,Y:� �ΟͲ�@"O��!�?J�<�V�O>Vbe��
OJ��M�#h��$��;W2 ��`H�\B�IH0�qbñ�H�P��{������S��t�{�[ #�t����[�IN�q���=�yBb�#��!g��H9�Q�(>��D�
r塈{���H�~�ę�+�8tb5���9,�!��X�u��a0���M�4�a��5Z
1O4�c���p<y��S���	q�[�{Z�#�J�|8�hjцL
s޹��념q��aJ��ē7i��
+9w^	���.a~��|[�-�N��$�5.F�O�����#y��Y0b�.$�H*!�?`s���QT��	��.4���t(D����s�~�*7�� ��1��O��{)z�s3�F�2SP8
�,G��w�"�X�A���h����-��'; ��nL��p���b9L]�K����Mk� ,P�R ��ۃ6	��x�'/z��qAP���)�;~�,���`�|DH�k4���
Bn@iJ2��H����P��2��#���d3���'-$5·�R�zO�c'��!E~,�O>a#��%a�~-�SJC8{.4���^~�OÞ�e$дFۜ���.ۇ7��	�'�l�2ȟ!D�(�0Ś$F42�QB��6n�8  �+#ѬH䧘Ohe�<�|D���.O�R�ӲjX,^e8�8�O|h*6n8B�!�c�C0]n��0d��<I��1OAt�sˀj����p�'�.��gO�����!��v�F��ӓ���Wm�3#|A�s�N#DN1(��ǥ
��Hƃ4U#:�2F���|]�h8�O>1�Ӧ�Ńv��آT��Md6(��D�
�M�&�/b��ԟ6p��D� 5񄸣uB_�!�XԐ'"O\9��-.�F, �C�"��1X4υ����d�"p�$)�P��>ia�`n��*�`�	HP��I��ƉW��� D��y(��	�yKq��?�XԄ�<��%���X$hA3~�� ȤkPb�'w\$�U��'r������8�t{ד\b>}2f(��A]��s�LF]��]��,@��iwkI�I~���Q'�p�� `�'����l�a`�j�4#,���{2M�1VI�آ��Ɨ ����H3��ԟN�@nD�^��-ڷ	��y4��0T"O�X�� s����UR�8��䫕șha�0s�H�u ԉ�g^��y��)a��6�:C h�u�];��ӑ2D�lkpm�*�(�0"�O�@��y����FW��.c��5{L�WX
�i�
?JQ�t"MB%q��YB�^�_��D�Ǐ.�O���C,�>�:��"�_ VRhL�֧��n�T�b�M<yf�`!��.�
��
�;�bL�e�>1��=6�SV�F��>�P�şQi���5M��uz��X�$�P?��jF��BM�7��P �i�p�����zǢ\R#+I鶹z�A��d�s$�%�����f��7�%+��QƟ�|�{�? ̋��ڥy�XL��i
!><t�"OBI����t瞅W���|hh�$�Lߛ��̓0`*��k�/MM���HO~�2�	��2��t1�&X<�R���'A�᳑��z�0L��Jr��9��ߊ0���
2Ĝ�wCd9� O�cJ�����R�F
�7*_�͛ �'����@��B��9�5�/Ծ�3It����p�������&"@V#ĂCp	pC�	72 9�!.��v_h�!
�j�$q#���\bB�h󍖰_" }�2F"�矴QJP+,V��	��?�}x��0D��`�/H$���'6*j��� .�v�j����'8:m��.]-!��9��C�BV2�8�'�:l˥�/�R(�t�4Q ��	�8Z\� �,��L�}�'ޣL5dm�G���V��3���0<�%c�e��"�Y����@ ���*(Wl܈��H�F���<�*xx�@ڹP�4A�II�=�'!,�k��-t�=9OE%O�I9�t�'K�Tl`G�@�l�2G'[��Q�ȓ�h86�̦b<hj抳  Л��'C�m(�ȓƦ]s� ��Om�O2��&�!Guj4x�@!=5�O2�Y��-�e/ǅC�9�!�ܛU���D.�"~b}zP&�#_�μ[ab(,O^`� O۟J�j��D%e!�S��'Z�UHP�_�`�((	����u��@��؊ N�1q���7ذm!e�0 �B�	�1��2яЈ<�&@3���/B:�9�S}�ʧdO�O���o�:��60�����*͌w��qض�K	X-�B≉1�� c@���_ � ��c�!n�e+�}b�K':Y�x���GC~���L���Z�(�����jO0��0�_8q3�qE~B!(ݜTy���	}�e��M�gm�fX�1`�+?FTqiŎI�~�F���c�%^���gL�lay�.�� t� ��=F(ƽ	e���yB��@0
�a�j̻f��s�&����O��H��"{��pŨ�D�&��ahH<	��>$��@�%ʻ,S��'G� ���AV�d�'ߢ��6-��8Bp��;
b���Ǉ�?�NM��.�"1��	7QrcՂ�<l���J�Aj�;�$3-���P�����}��i�/>�J�
V�o��0Ѷ����07sF��r�(+�Ҵe.9�a�q1c�
wB�`5 ]f���	r�  8����\1�G�"jj�cc�7�̠�U�j��(l�pd<@Bt�	N?v�;�ܕ.���z��
O�\�ɑ/`�uPd�;��y0��_;΢=IN9v(@�AukB�� �ᐇ�McG
3�~��$��'���dC�b��]�!a�.p39y�	���6�DzZwE��4K�"`f�ݒk�2�P!N��!Y����a��B�I�L�Th۔��,(�  Sŀ$<�T���$��d~0�Ҳ!�
�PIC��?�AuӐ�svL�'8t���D�Ut4�2��'����@�E-E�4�0�;OD��ȟv�A�'ű<0��P�i����^Ht��:�fx��T8g"b��Ma8�@3��#lO�h�&8(��y*�#d�Y�vF��fl��m��8!�ORh<y�L�P�<�b�d�`�d��C\�A����pB��4�=���A�82զą`���$�X��B䉢F]>�Y3{�e��F�=r(h���E1 @2�oIf?ٔ�>q�g�?,ڀ*v�8J��}h�DO�<�dJ6�=��Lx� :dh�o^d�<����(��!��	�xH*I����W�9!��I�~k8C��$!��)�E!
�_u�U7��B�ɏ�\8"�ر��@Ǔ?0�C�N�	��޼rL��A�$��B�I$2Yb8A�KJ�1c���F�{P�B䉔}f����ء_��#��
h��B�ɧ~��w��hD��4�=HĞB䉼!�� @,S xg���!&`��C�'a�N��)]#y蘌:%�@��C�I�1�H�R��0v�vH4	�<dlB�	gw\�ר��P�*0����`vB��B��1i�nO/
���/ҝ3EdB��D��ҵ���Y���
�x�C�	A$!h�"
@Q X�B�W.�8B�??x͚g�^�5��|�J�5d�B�	�r"mQ�UZ�0�eK�&F�B�	+U�Tٰ���	���H!FѢ.��C�,�V����ՃG�35Jl�B�)� ����M��	��ʕB���v"O��a�J �����LQ}�*)0"O��bON�K
��A
�m�r��&"O�<)�<y�2i��B

+��Y�W"O����ÂW� X�� y=�0�"OHQ�Ae�'��}� �/s�૒"OVPi]��:i��Y9�8��"O�1��NQ��� Rg�=�|�	�"O�*��ΐ�����H�Ӷ���"O$��e`��^�&�i%�@��AA"O�G" �!(`d�U��a�j@j�"O�l���$���9WIZ,S��z"OBu
���SL��p���C�"OBM�Ц��e��sGM=!����@"O��R��(*�t8�(� 6ӦP�D"O�-��F)n\<�m�s�z���"O����O�x�����.��͋�"Oj�ˡ
ÖO�j0�נ(�\!
G"Ol�ڗ�Կo#\� p��2ܘ��"O�(�b
�i˨Ec�_� �"O�|j���s�Ρ����$_ r�c�"Oڱ��X�d�VQ2��F��"O����B/O(�c���@��C"Oؼ�ᄗ�3�H=9�&IG�
���"O*��I-5� Kʏ?Ѵ�@"O�@jr,�!Y1�QCv���ҘM`U"O��U��z��W���B��:c"O��R��H<,�$�ڴn�x ��"O z5O�|���c.�z堅
E"O�ّL��)k�	�k2�z&"O��YS$N�S�293�̕�mJ��
D"O����.� \�dٛ���V�]�5"OP��F�ET����P� �x��"O��T�t_d�x`��9�nU�"O��PcHOJI�L��-
p��A�a"O�����]�~ь��/U�1�����"O�̩���N����-K��Q%"O�`W#��y�pHc���=��"O0�*���GI���«��e��Y�V"O��g,2>��A��G�g�t-�u"O���s��4-0�d�I�IL|�"Or}���V���(���"���h�"O0k0���P���B�ԭ���"O�,�qGV�a(.dK��͕2e^�q"O�l����K�"�	R���ITFPsU"O��Thݢ:��!rɅG�Hz�"Ol� ��
V��ѻWI��c�
k�"O�	�@%P�cF�=�r�J5uV`�0"OT�i � <�+��ɻ^ZLJR"O�ea�"�ZeT�G�.�naA2"O@̢T��6� ��3%��Q��"O@���?x��(�d,�e�*uk�"O�,X&�����i��9���a"O�8����IH8L��h�1���D"O��r֭t�@A[��޴[��Z%"Oĥ�)�k��9��9
��¥"O�@h��$ߘX@�d :V� ��"Of�[uᆅ2���2�^�ntp+`"O�`J����l�^�s�F#s�$�k�"OV)�B �,g0�����*ġb"O,x�Q@<PV� �����J5"O�5
 �D�p�
�i�!0����"O�h+c��c�p��!���� 9"O��+�/��Q��%s�D�������"O� ���a'S�h��X�3b�@|Y�"O��1!��D��({S�Lo���0�"O<��CƏvl�\����S�R�"OL��f�7�.Ay4,؀	��M�4"On���
�'�f-�J�0�x��"OJ����D���J�)����E"OT���ʜ�Ǆ��)�_�N9����\�O�aS)��CK��;�ڲLӪEj�'��Ce�Db�b;;�"HӍ{��)���_� ���#�aRJ$���W�Z�!�d�U�� D�
�=G�)s�
~�!�2�Е����w6a��f�&+�!�$�&W��p��l#`)� #ʃE�!�%tpB�k�`	(s�Q:#�@+F!��^�~�s��|Ҥ"e/T�w�!��+vi��.P�	m�PR. �!�d�8J0@�@N��N9���E<h�!�D2Eĵ9��#$�)[�%x�!��1y��@�T��.e�A�A7^�!�4
K5B�$���� i�e[�'�(5-}^���b���l`(HPN[P�<�0�1�:C$>P��hY���L�<ْ�ACᶥV$�!��)�D��G�<�w�Me�5J���N�F��H�'M�x�-)F0�啂0̃���0�y���;^(���@Ȗ,wJ�T�c�Z��y�$��5���o����(�y"�='�uIw�N�m�����d���yB�\)%Қp���X�`�]�GiT��y�o��l!)��Y'ef8�j�C_��y�b
O�2���.Ͻ*�|�z��T+�yř
M��)�$&J2 ��!)����'�a{R@I�?RH�ӠAU(�������y�K�O�z�!��[hg
4�BI��yb��+7�BU�d�g��������y�-��:�3C��5\��m&�yRiZ�o���I�ԓM��#���y���J�pKc�ԛ����FC��yR=Pu��(�&L�,��JU�P\�<I"+E�+�����O�>l����&�c�<	�ۘU���:92��vʅt�<�E�O�7^�1U� ;Oɪ$H�Et�<���$�јG+�-k:z�S�MT�<a6oQ���S�-�.H�3��j�<�3��`��*d�˶1�(%{vO�d�<�`/9mq�͈���18-����J�G�<1�*��a��q�����؉bd�T[~��)�'L� ��2��q$�	��%�;t��[Q�1閯US��ܕh�`��ȓ<�P�	�˙P��j E���݅ȓL@8�U�X/R7�`���nx�ȓs����"��7c�j4�FS�8�~���_����e�A2P]I���)
W�y��W���ٵgo� q��yv=�ȓD����F&��)�lH����Y!��ȓC����/Ń:� ( �> �04Gz��'I�dC7G�6�8�'�J�d�
5��'G���b���� Jf�%%E<M`�'�f�Z��:��4� D
0N~��`�����,B;B��E�.t�}�ȓx��]���&c,��q�'>�Z��ȓ�<�������'�� 8�bɇȓ_lH 1��؍;�jT�QAV�*�VX��@<9
t�Ҿ�!��J�ΰ��S�? Δ	r�Q�7���.E�x�QAP"O�	�S�@t��$m�,O%���"O I �iR�_�jt���ˋ(	|���"O���Q*�0BZ8�C"`[�D��"O��3 ٤A �!!&��]��I�"O~hz`�Z!�4ˀ�^���[U"Ot�"wτ�y���Aʐ�` ���0"OR����=/!�MkèB�/�|�"OD��%lEG �#�Ɠ�A���`t"O8�	�F�#q�"�^�k}�bs"O���e�� �.H�6�ـ5�d�y"OTL�"E��"W�)Ĉ�&x(�"Ob�P���9Rܡ������"O����J�7�J` ��Ϳ`���+"O60` ��i��Yz@׻f�d�"O�D�Q�Sn2�a��x��y��"O�A��k��y�ڌI$��N�T%c"O����G/<g�]��ؼ~�uaR"O�c�l�q�F�Θ�/u��+E"O��
׏'z�V�Q��Tn
P"O���G��r8r5p��;bd`�"O�xڠK^��a�p�ņIf�\y�"O����K��N�9���BO�"O8Y͒���s6g);�m�"O���#ݜ	���W�[�K2���"O�2r�V w�	�#��E!&�""O��ɄC� l������h��`���;\O0f��?[e�����2�~���'d�L5�!�,h���0դH�2�P�ȓc[����;�2 ��5&z(��IT�'P�x��8sE�A�d�L-޶���'�@�i̄YO��˴�	.O����$9�S�4d� Y��MU/B&:�0�݊�yR�H�
ҘU�d(S�"����Gғ�HO��=�OÊl��9% �j�D;N�0�
��	)F�4��FQ96'�X8�GQ!|P!�$�,w��(�1�G�-p���*:!�$S)MQ���O ��Apń�#!�䘮Kbl���M���	۶U	!�d�3F�X�
0���{!���C�Z�}�!��_���@+E(�����2�Z	�'>�|�H��)���>A'D�7O
/�y��#̆�)-.\Fإ	���6�O�+4À�)������ON�r�"O>H�CR�6�p�i���#;�|�"O�Hyde^%.|�r��� $��)ң"O�л��֖VXɣ���Pd-��"O�j�e��Yj���ğ�T�P "O"u13�Z<]D��17��0?�=:�"O����l	TQ��՚|�L	�"O����D�Rug����=S�"O��!��+����v�'�4���"O�����Y�> Z�T�- 8����"O�U���ո#�AB��h,�0�5"O~��Y1X�I�I�1R�B��4^�<!��@'lr�D�7R6Da �XU�V\�<1p�spĸ��{�4�'��s�<Y�ᆒ-���H�̙;��}JI�D�<����	>9��>`�����ZA�<I�H�,l�a���@"<p�N{�<U�oOƘX��Q:C}�AQ���R�<!2a�e�0e[���7M�^����\P�<a%$__3�=[㢃-?``����u�<�c&��X�
T���13�8�(�}�<� "��@J�d�<��F�2�d�I"OH�)v��;��)��@Y��"Or��Q��&�90��t�G"O�����M)G� Q�詪�"O2LZ#l��=r2��K�	z�����"O�Yo�>�"��䗌ax�H�6"OPԉso��/B�q�1䛀l0 �"O+�!FR��e#�'o[>�ps"O��hj��.o�tpa��Sd]B3"O �
�������v�o�|�"O�LAAM|�`�0���:=�4D�"O��	�B�"J-
ŃakY�h{*H��"On-�1)�3�f���)ӆ(����5"O�<K1��LC�͋f5=����"O�к$��o��D!��J�mt�Ӈ"O:�́�,���tJм7e0 ��"OD��ƟSed�ʳ��?��a7"OL���CƦm(�b��X)@��9"O�A3�KRi���tF�1O��\��"O� �f�
"m3~@ F��>q����"Ob�$��f
|}hXI¬b+�i�<	5' �&��=�e̞�XO0@+��k�<�7�8yxб�b����q� j�<�e��R��Y�.:7j�:g��b�<�&L�_'���4�H(�lt��Mx�<!q��4)�� tE�&y)��kW	Tp�<!�*��[�*�@'�O�z]l[�i�<�S-N��Z�Z�cUI��lS3�l�<� X�NTd�Āx��Ȅ�R�<�4(EM ��h⌍�%�֤����u�<�恟�_4�p�я`��]B�+Z�<II~�(F�.�bu:D�~�<(�!�"�(̏+�h��@GR�<�i\$��\Qdɮ1��NN�<�#_��ԕჁٻ��Ѧ�t�<�s*N�*��mH����iZa��Ur�<p-֢9�@%
�׎y�Ԝc���p�<A�eԄ?�� �gϦ3���hk�<���"ޠ�0��./&�1�Mh�<Eɓmf0�h#�P������b�<q��M��"��Q�Y$�Q1�^�<aR�<�ػs�� �Ɲ�@A�p�<	B�_nHYgCŃx��(� bCU�<!��/Z9���ـJ��1��*�Q�<����
�v4}�dhG�UT�<IC�X�Z�L��*˱Hc��!#H�<q6�E>��H8 ��)��X"CQ�<	��f1�s�N��@���� R�<�Q�� VH�6RW^�����d�<����(�z|#r�üYh��U-�w�<�g����ؕ/ 3l��y���
H�<90���Z�ls�n�'!&>l`R��Z�<yVʖ�*eĉ)�~��4`�'L^�<q���/�����H�?-le�#B�b�<��K�6l=���N�7z�a+T��U�<Yb$Z2k� ��!(]�72���W�<	� M̾��p��2���!��M�<��ϕ�=f��ǌ/?�( r�I�<�e�
1U�-��N
�I-4��%E�<9�@��1`c/�&L#(㓁 z�<�!�O�5���)P��J�.���h�r�<	Wnܺ;_, G��q%���#-�r�<I5nC=A�%�����):������k�<i�e� ��`��щ40a'�@�<� ����
��C3��g�G�Z��=B�"O���uB�85���S��׼y�2��w"O!96K� on8�"�ۦ3{�b"O �8B��t2ꅤykf5 %"O��珇;WD��،4W�y�g"O ��l�q����-����b�"O�إ�S��L�Q�X1�4k�"O ��&�>V��a��
�vOH
d"O�P�j��h}�E�<4Tz@"O4P��@�C����N�K,�0d"O�Ŭ4PHJ`�#���d�ِ7"O����������ʎ�Z��V"O$<B�b0X)�	�8=���2"O�쐱(Q#S+�͠ B�O<vt��"O81�*@��VYH&���I&dq�"O��Rk��G��� ��@��e"Ob��N,�&]i�xBb��"O��s "$dK`Lڳ �R�Ip�"O�pr6*�>oR(9� ��ҍx�"OB��f�ǂenФH0����M��"Oy!�,&���L�%��<�"O�I'd�8�fhኻd*x�"O��8��	�T��I�6�.-�"O�3�T*l�LT񠬄�N�4%�"O@|��N�*j|u@J�}d�	�'��Ę��ո_�P�Ë�a��
�'�Ph2d��3[V���BT<+ߴ�9	�'pl�y���"�\�Х��.*Z���'�(��/ҪjVZ���i ��R���'b�	�g��8E����lD��'�z!a��@-[�l���'�rA3�'�!��D�F�|<IUW�����'�氻%��0��D� ��z���'�h� M�\�@�D�^oR���'
h���A����ƭ�"S8��'Y�Xa���-&
Ԉa'��NI8d��'jd<Ѐ��"�ER+��G% ��'��Ń"�W%?�"I'/� U�@�z�'��س'RS��V�I$�M��'��8&��KHZ0O�$AY�E��'a@Ѓ\���)ZGJ�"8��Ț�'ς ��/H
f�6��irQJ�'/>����9O�����ظYv���'�>��p-R,Y�.�Ӑ�E!]�b(p	�'���N� 0V��6�
�Y�V�r	�'�.���&H�g�nI���0R�B���'���	%�6_�,1���VE�u��'�"�б��/�~�+� 	3f�$
�'%4h4��B
13WI�%P%��'���G !^1�C�!In*�Q�'�"�b�,s:�Bv�B�A�x@��'��'��uk���`�ڜ5���!�'3���c�"kd�LhW��-�|Mk�'5����Ŕk%�q�Nʊy�z<��'���J���Rh]ڰ���r�PP�',�y2ש� ���r�'@�p� �'^�����(� ]Y�*�M�����'@���$��3� �e�;Bo8t�'��jׅ��C���U� ���%�'\���1�����z��ع-E���']�1Bs&K0�	є��/t�e��'e�hz���6^d�ӌE3&�ٛ�'L�]A'��LݸV�
Ј�'�԰��(�1*E M���5~DH���� "="���f�~�E\*	����4"OH�I�%F�R�!�>G��:�"Ȏ��X�B�*�I��Ӗl<a"O�@�D�s��!�ED C�`eI�"O(��%o/\Y��k��U/ �r��"O�5{�ˮ,���	"#�7�h)�"O��0��%�܁*0HZ����"O~U�Pf�<p$���g۸&��M�q"O��#4� 0R������&�`3@"O� #��ߠ]�rl�Ҋ�<Q2�$"OZ)�ˎ-P��a� �~� ��"O��*���(�vU�7�ƧEb�h�"O&E��(�:��;U�E�i��"OD����4��¥�ǆ<"<��"O�L+G	���+ж\�D�Q�"Op(j�.�,�Y��;Pր`Hq"O���&�W*)c剧I݀a���q"O�u�4yl}h�j��W�D��"Op���H�j~fu��A=sD+"O�0���Vnf��	<CFx��W"O���`ë0/^h�b��+<	<	��"O�����7��*g��
��0#"OR9C1��7me|���oO>A�"O���3D�bХ�s���	E�E"O���F�R�>��=ÑmA�j��Q�"O8QpA�W��iR��="j�� �"O���`�6j�d���5Nn	��"O���W p��%N@1H-� R��E{���~ԉ3H3+תՋ0�#Ly!�d02���Fŕ��V ��ai!�ɘc^�M�Ů�(Oά-ڂOZ�}u!�$�^���pA??Ѣ����`!�$��^�Z@�+KϠ���^�Y/!�FMἼ���	Ġ�JZ�N!��a�r�%��0�d�I�8~�!��Z�"PA���Y��A
��֛�!��r��Ȳa/;ll�Bg'��)��	X��D��m�?���	8~t��#`�:D�\�N��q����l'(��4�R,;D�����F&fd$ ��n ;�ڭ�e�&�O"��1��H0� L�"��I�@	��I{B��t�p�P֪�P�`�h��� 4B�ɼu�$�d�W��`AB"
�-�B䉾��]3.�<,~vS�*��{w�C��>/6"�⡊���I	��-'�C�IK��Q�kW!*i���QM�|�B�ɜU&]��Ȇ?�(M���2�XB�ɢ)���q�_� ����!^`�C�	����Vd�7%
��ݱL,&����ɥS�上�lZ)]m�	�&g�{���d7�}��L�e�_"s�J@[��Z�t}��5n�X���X�_�F��C��"P��ȓ�~��/�F�.��Q�"H�R��ȓd����-vG�`r�ŝg����G^�(TN�j�^m���"~��� ?�	��c�Np����A��̣t��T�<�H���,��!H�Sb��j�<���	�a�d����r�~%:�)�A�<�B��2W��,"��H��f�t�<B� gX<�D*Ӏ@�4�E��I�<�Fn��/"�IVL� f��%����<��	&K�J�ڄ!� ��l��Kbx���'��Y5�^�h����<�TT���Ib�D���-qe.�`"!۫����A�:D�� ����ݖ<��2S펃-�\X	G��2LO|zg/�}fx�Z��ն�r���"O�A)௉G-zqSs�g��l�"O��Uᇟj��3$K���8�S�"OZйń�4i/r�x� H��8��|"��,�'�� �u!	�P6�b��I����M��6� ����a� ��ȓ^^=���͎W�
,	�ʞ�APB��'Ra~�a��R����� [4I����y��BPz�aBT��|�|��/���yRe��>py�Q�)�~$
ů�8�y��B1���"$�	�$��1�q闟�y���5�r��	#PZ�I�h:�y��
8�$X�F*�@%Hs.���=a�yRL����,!���)����D�4�?a���SJ#pظ#�T�h�dIX��,V����O�mI�Y8J�B����/Z��y��%�<�g�]�kG8�قEE�d�����JT�1O�{�jQq�aK�]�̄�&N�����O�|�"���Q1���A<5�;u�}B��[�&i�ܑ�&�|�<�A��1*�������<0#b,z�<�R�
@��ըW7���*�l�[�<�s/��F�$K=h4f8���~�<9����)��MZ�0X�=h��O�<�Љ2yp�����5s�M�T�IM�<Aw UaZQ�3KN�NN����M�<b��
�L|�Dυg�����DOH�<1�=X�zm�5k\�	����(�F�	E���O�(�� �	�"�r�7LV��'[��!1Ç+q/Ti���Dz����'~ԩ��
���mS�?,f-	�'t�\tBS�4c�}���ʆl�p{I>9���	����]1d^�z,�Hz!mI�E!�$�&4�M�El�WC|��Ն7I*�'qa|�HO$�� pꜱ?\�������'#��'0?�x�$(>q�y!�B�XҒ�9u)3D��S�Z�5Ś��t��%�pL2D������=p5l��b��>����D1D�Ȩ���[�Ɲ�)[;dV�H���"D�,p0
o���A�>:l�̠�M>���d.�'/�P[f�¶U<�;�H,�F���.�4���'�g��J΄Z"��ȓ��"�`Q/��jg�4����h����8L�
 �O�r�ƥ��H��u:��u,�%A`O�YbP|�� �����O  I����
���FR�S�RR�bK�+�R�S���>T�B㉶eO��!�e�S!�sc�'���F��S4w�x�� .V�a�ᘳ	�f��C�	�t4#�핌>G��6ɗ0j6C�I_�j�:A��4X�"Q+��ֹ!�C�I�24���؆�D�c�eU"*�B�	 wAlT#M�s��q�œ0��?!��iŒ[��0��H?}�%K;e!�$G�r�)�� A�A�u�ӏS�"2!�D�$sF��@ˏ[�"����q�!��ޓ��Yq �nt����!�d�Z�r@�㔂!�	sVS�Pt!�	\��x�Of���feW!�䁌7erh�c��t�~m ����!�B�fsJ��F�
�t� ؖ�Qm!�ě�p
Ɖs�.��4hu�̏B��O����|z�@�<HNJ "J7�d���c�<� ��2��H�"pf����H-���J"O�0���m}&�x���b���#A"O60�"��,�� �@I�X��'|,�@��l�|`a���{�p�
�'�
Պ�mJ-,G�!"�� �eL<=2���'��p�.ĲP���bc�ҕ����)��H׹*[\0"�\B��4-J����O��Ex$H="��a��B�	��*R
ţ�y�@J
%A<$�����5�����y�"��<���OV�qF��@ l��y�`��gF�h>��2�+ �yRFQ�[��$甏k7�<.4 ��'�@	�b֠M�dY9��:ig����'�ܑA(�����s�"D\i�`!�'�9�/N��H�C5M��h;p}��'2�,A��m�L��,>a��}j�'��u�DA�iv��i��^�Z�Z�'�:��5ǖ&��- �Z$������O�"|��	�I���Z��`IFr�<��E̝ �\a�D�	M�mst  q�<Y�Ɓ�r����TF�7�(H3�In�<�Ag�8���`���2&d�bDHDk�<�o�(m������s˔�q���R�<�2��B"Ȋ��ń]�~!�p͝Q��d̓��Lq�
A u����ϓ]��=�� ���I�,Y.v����uӥچd�ȓi�@	ꁣS�kN�<�&�١cw]��If~�Z�0�-�pE�;$���!M��y����dÖn�Zt��LR�G>�I�'Hp��!��.�3h�=�j�	�'J�dy�MN?/`T	@�_���#�'w@�J���=�b�9��P�E�.����x���+� �C��.�z�+�F���ybk�"-b�V)�$�T`��c��hO
��DP>9��C����&�.���Q�T���h���0uڵ@Iȁ�άq����=D�L���u6�A�!�]���R!�<D���%"�1z��-�N�;k�
ǌ:D�dJ�$ٿqnji%f�$vHL��E�O��=E��l.vH��K��6�=��+�y�!�$�tH0�7b�=��ՀE뗎�!�$Q9I'�,�1�'7Y������'3!�$U	kW�=�&��=&W�L��%�f!�G�;t� ���O]0��!���
8��e��
=�T���g��\�!�$>0����xͬ�b��YA�y��'�1O�,�䔨sm2䑰��LD�(`"Op5�� ݾ2�9�� ;�Hrt�'�ɧ+�3�$�"���Vb�=��1��OMy�@SN@�����]4��"O����G�\�u�<IV�� "Oz}�օΜw ٪G��>������w>��#��0^l��#B��M�ȹ1�1��?��	O:C$� ���vo:�(�,��Y�!��X��ႁ�̴��*0I0a~!�$�';$�Xs@�΋Q�>�Z�'Ң(��O� ���-�HI���0Qg��Y"O�X���׺P��)� ���[
a3"O���I��RR�D!Oa���"O���F#�5$�]0w%�@^6���"O�M�Ǧҏ[���
�EI6v�Q*�"Oz��`��vؾ�k�j���t��"O\i�3�?N��l��ő�@8��"O,��3@M5pgTp1Q�0/S��y
� 0!��1p�P8S���"�~e��"O�R�ovR@�`�D}Nr��"O��DJ[�}�b ��>�tT�e�'x���BG	m�Q��)�H%���*D������1Ai�l0��W�\dj��(D��bi͢@Yʝj �ٔK>�C#%D���vhJ1L��R�����^;�8D�H��a�~��`j���!	9Vp��k5D��f�J8M��1��	39N��.D�X��嘞3FDpz��L�4�4tʓ�>���?y����Q�\�
]HX��b"�>P!�ā�y�E�F-\
?*��h0Gُq2!�;hВ�Qn�]��Q6��$!������Ń	w	���D��!�d��}��=�F��Q �P�bC={�!��]�z�Dc)��͆�R,��'�6��B �zjrIB�NGZ�Ty�'�����L�?.~�ԹR��R��!��'�Z92�!JB��!LA/W� ���'H����_&�b�K��P���
�'bD��h�-���� �U��u�
�'�fthb߉J�];�D�Mf�i
�'��i�7�F�a�^L����5�l��	�'E�d��% jʒ�י6�&`	���'�� &��2}/�L�'b	e�<i�/tG,�{�͘�p@ÖK�<qpȏ�O���Y>5����w�QH�<E`LN��)�"�8t���EaO�<9�l��;
��{�lC�5�ś!m�N�<iQJ�";榙��[���ۢˆ՟�G{��IQ�$�\Z�B[�E4Z�b���b5��,�S�OC�E�禔�e��1J�H{٤�i�"O|�s�61O����W.9�$:��'b��'T�a@�B+x��)�4K:#Z��D1�S�O��a��D�&e Y�բӬ&����"O��Q�@�<QJ�ؐoE/!<�89�"O(���n)�\�*H	�D,!�#"O�y��7*�^q ��B]
LY��'�!��yZUJV�ڪ7Ȏ�JY48��'�ܴ�E՟i�4�j�a��1�' čóۺ/Db��),ˎHy�'�\�:#EXR��R�a��v<XA�'Q����S�9��AWI�s�����'hJ�e�7 �u(��� �v��
�'�jlk�b	>&P҇hH�t߆�P
�'�F,(�����b�Y�ky�D��'i �0ڃT1���F&�Rq
9����hO?�@,	�&r��X5���}:�Lc�<�NU'��˒j]v_�*�,Uv�<�f���o�Ƒ+5��d�Q�O�v�<)):��@�������1V��Z�<�T�8�����+zNTu��YW�<���D+<����B�o��}+��L�<�m�w�x��	P�J�U���P�'a����P"d��F�֡V�ڭ�5�A;��D=�S�OL���̽/�ڬ!�㊐WC*�(	�'Nl��!W	@ r-9�+s�9��'�fu2��M�8.d��v��%ll���'{�<#u�@;	��=CQJ����Z�'5��y���r�ꭈ�֢�Pk�'�<لa�u%���� '\����'��)q�ڗ\�2A��� |+����'�`̣VF%zPJ]9s'�}�"��'���2�n��	�h�iK�Y8
��� t�J��=]w$��e��X梨�W�'31O��cweB��VQ�2O8h�*TR"O 1J�� �`@��[��m�<"OpY�U�R,��1�g��%�©·"Oe��%�#;�P`*J�n�1R!"OB�y@�Y�֭a2��u%�"O~=�F'H5A ����Q�"O� kTˏ�1����4���r"O�s�*׆N�P�q0!�������"O�t���L�@�>u�$Ixe"O��ap͐<��[�Fϴj�9�"O����Y	I���jF�ұfOxy�P�\��Iov� YfKF@����Q,�C�	
z�A��L��$HIi�zl�C�	�q�$���O�7P��� �G+
���D~��iv��8g��@	
A�B�2�3D��S���3�Tt���-��sd2D�k�%�x�|���E���u�n�O,�=E���:M.(@��<��Y��m�i!��2	b�K�e�F�����E!���"p���� ��I{� s��A��!�ʶ��8	�Y:BʜC�,�P?!�$��r�T53!"O=S��1'-�8,!��X���Aǝ�$)VK@�m!�d�1V́�LہD�v!GI�7j�Iw��(������}����F"�M��DR�|��)��::2� t&̍W��)��6��B�<G�r�1�G�5s��p����/]fB�	BVx�񔅙�(�9�`��M����:�	1`>�*�,Xdy !�j�1Q!,C�I�ߒA�5LԊMe��2cΟ7$��B�ɒR����1ŗ:=�}J�A�8�B�(`a� �B���z:��	���?wVB�	-6��3Qj�'r�p 
U�vB�	�h� a	� ,:���3�b�wHB䉋Z� u �)�LL���4}6�=��� �\�"�ُtt(�Ӧ
�fP,B��$�6�{#�SzJHW�HH�B�I2$�Ŧ��7#:8��@F�A`�?)���ǔ[h�h��A����ۭJ�!�70�Y�cR3 &bC�H�!�©H|��7�+K�A9�/گvl!��,B���i��{�����ޮ4��2=O��b�._2��%��V�Q�"O���/Gv@�7�
�D�v�r"O"�EOƩ(�����:l� y�"O:��ǉn�Μx��ҧ%��2���|�rA�I�%������ضK��9z4�'D� �fJ
�_��C�-˲f ���2D�H
��'NkF���N�{��iB1D��"2G�x���Qစ$Bf1�$�-D��Lߍ@�x�i!l_	P�|�F�6D�� ���1�bqA� ~J勓�6D�L��߮{��YY�.�E- ���O?D� �����x�bvl�1E��� ��"D��@����x�HQ*�+R*8d\��?D��Z���DJx��E:�`��u�!4� S�&��I�!��b��k�#�G�<y��Ь,q6�S�iv�m�Q'�@�<A�-�aj`1x7�ݿ�����|�<����h��+��:�Ľp(B|�<Yu'Ew�����J�*�釫Q|�<ɳ�ɂq ʸ"R��1*%xbO�@�<� �ً94�"�%�#>*�C�O\z�<� �������yQ.�1a�l�#@"O��rD*	�C�}2m+鎅"O�|���!OF�|�3��v���B�"OJ�`�JW� ސ��C�&ӊd� "O������H��[0�˙?2�)� "OJ�Yr�C�CJys�'Y,l	��"O��sv@�>[8��g܃}(�TJ��'z�IX~2�K!D��@Dǚ�6(ܥІ���y	A/Q�$u�F��+�BUi����yrI�.��!�OJ%O�M������<9��d	�21BDQ�&8�M���B�|�!��FH2�I�Oѹ3�(�Q��Y.!��s��y+�N�+���K���/!�0U�P P�y�*��C08�!���M[�C��Ϩ`g�к ��'�ў�>�w�'�n)b�l���-�4�>D���Em�9Z��I��"� !S\��H D��[���'6��X6CK;���g<D������}���[�a�/w��5��F9D�ĺw(E�_��3׊P7l�|<VC䉖J��|rѣ�/���o)z> B�	Ӣ�r�X�Q��tCWM�2$��C��I�k�ۧ_�����Nҵ��C�(Y��!ZR,�/���IT��D�C䉲qf	�P�m�:�KՊ<Rk�C䉏N-���*Q�|g2M�����Y�C�I%�\�C%��!���aaiO�v�fC�	�V�f��҂���ʉ-p�b��d0�I :A�HY�h�8/�4s�K��,C�I-l�a��B�J��<��gO&`C�9s5f� '-C��s�BΚ]�NC�I�?�tHs�o�rJձ��+��B�	�%����AC$5Z�V�%pB�,3�.��5	٘h<�h	q� %لB䉅W'Zp��H�r�zĈ�k8S��x��H���4+,*>e�f�65���JB����0>q0�-h\��BHI]R�!�VQ�<�G���\���R�_�@�`aC\u�<	 �!('�@a^�vd�V�o�<�a�R<љ#�XlډG��j�<��*kD����X8؅Q��M�<)G�Y�<��xh�%��J)pQ����I�<�%J݇�b�U��>�r|���G�<IU擫�<�)��"{D�Rc��z�<�֧�!��Y���Č+�6e�T)Pu�<������`#@�Ҟ{���Eo�m�<9ө�5a�8�cU�rA�tC]A�<b�اݔ��v��5@�����R�<!�)�R��B�je2�����d�<���V�_���W ��q�,��e*]�<I'MJ�ivh�w#K2hL����Y�<�#�R䤁�gOdk�"*��B�ɨcn��1���8Nu�4��3PC�0���Vˁ O"|�R�Ɨ�5�$C��3l
>�i�.c�r8h�&�7-6�B�	��Pt���\�  ��%߬b�"B� Ymzْ�B=Q`'�.^�HB�I�t-@u���" �Q����E�DB�ɘ4Q>�z�-��?� ��S�G�cXB�Id� �˷�uŅJ�̜==fiQ�'�4��q�0#��h���~�J���'T�c�I�d���Q��9�b�a�'DQ��j����n	����'� l��C�@�D�zG����i���� <�҇�֊@4Y���M�fܚ""Or�r⢞1�h���w��AX "O���A�`+N��莆"����|B�'�Q�!��m��a(vg�	0.�p��'o�T��̂��@�T+P����'��X���h�8�b�̖�N��83�'�|[�b���ʀ�PfUJ�i��'�f�+ub�
N��ۄ	�Hs�%�	�'~�,Ɩ=Sv��N٦.��+	�'�I�6A !��4��?�xZ�'�8$�oǨ�5�t�X��L���'B�|��Y.)��y�UCY�L��c�'_�m����.���6��3��d�'O�؊w$)v�<8��Η*�0�[
�'�6����ˉZ�x)���L�|��'c>1!f&��D7������栓�'L��P������4	��(R>1p�'��51"�8]f�#��	vq����'��5�' �q�h�`3�J�d���R�'q>� kJ<���SIA�^L�P��'J�t���֌����g�X$�'G�a��I0�5�d)��I���j�'p�*��E�ZTD����Vz��(�';(��)�'�����ʘU)|�����+O�M��
^�z~���cT��r�)�"Ob�K���70�$�S�!{�)e"O�
4�ە4.��`M� ���b�"OR5 �kW!u�a��L�iwI��"O���TlI�z�ڸj��FLwL@T"O��1�kV�iCH|8#�
�#�"O�����K�~��р���:v
�2"O~\ځm@�'��)+D�}��<��"O��Be۟}jh�"dD=Ab�Qa"O�m��͇92C��-���b"O��c�u
n	��ŭs���I"O�)Sp,�x��<��gD���"Or��`�r�Fix[��eH�.���y�[�L2����&I+��A�@��hO����&k������V\ݪ����c!򄃳�)�&�G���4%Þq!�$�H�����K�.k��c�X�!�D��?`P��f &U�M���ŋ}�!�
�[��I�t)��>D(tR%CH�*�����(c4��Q�ـm���{VB	��y2Щ�n�;�.ЈR4�h����'�az�)�>M��@p M�9���@��X��yB�Q&V]b�9��ڗ4���B#[��y2�	49�x��B�(�:`�Ò	�y��[�x�ʸSu�P�*8�02�$�1�y�[�H�\0$�!nB���(��'Wazb�
�K�D쉗͔����q��y"��Rꨕa�I��/R,��]��y��+2��<3�@�6ቐ����y�ƅ�dhXg��7s*�@����y����N��Gǅ�-:�������y2��1Nb��J��%F�uZ�A]�<��'�Te(Vf�2�b�[��e$�@�/O|������`BA�	t��"��H-(�!��;2��A���G��Dx` /�5~�!�$QE�����Z�+u�1sm�;:!���X���$ .�⥢Q�
�!�!�d��A]� �ʈQƸ���D�i�!��(��ҭ@D�~���L�!�$��DC�X�F@���u2F�/�!�� d)����
i�@�a��!7n�� 4"OբDKE%F�n���E;Vh8�H�"OF�	e�7; �[�L:�=;T"O��KQ̓�jHS.ϕU-k5"O�cS
�/0�!����@�(3�"O
E�gKV�L�r6-Սh�<t "O��I�#I�+� �X�B̵\��r"OjАce/'�i5B�4CM��e"O���,�6/â�S��X3�Li�S�������CI4P��2 ݑh��B�ɦ.̈́��bJ�?��9���9�B�IxX̪b*ƻqs�ա�L�J7�B�ɎC��gK	
C��Ě�Ĉ�`��B�I�T/���Qi�g�h@�.��tB�	�*&���G��<t���k���<B�	:�6T�Ћ�"I]�Y�6R�R�B䉟O �d�'(]�n�#�71B�I'G��P�-��D�V�
�j�o��C��:/���Ȁ�8��m���9��˓�hOQ>!��E�۰dpL]>�^��Ai;��S�� �C�ύm� y��[$���@e-8D��{4'Օ�F����7J����F:D���7��-�������0a���o3D��6+��)�8�����(R^x��R'2D�4�@-ֻ$��"�.ū��ӈ2D�,�����3�y�*�9Vp@�'3D�R���@ca�Z
Q	@}�S'D�|���ޡ1J�->v�:�� @9D�lZ�l�)���3aI�"*�I�7-<D�t�Q�R�cbTm)�U
K���A�;D��{fGL�A���	6*S�hD��rC�$D��I�-�(�؈e�O�],<�XFO#D�+p�9��9�(��
H|���!D�$��G.$�5Б執!�h��$3D� c'��P������E8�aT�+D�)�O�1+����}�*D�A�(D�X[��ǘ�LLʅ�U��H+:D�iel�._=z�!gO��]��h���4D���4)�Fq��{��1HƼ
�# T�\����,T{"T*O˓K8�u��'�ў"~BtC�+�R���A� ws�C�l$�y���X���F߸~��AZP���y���H��J�fH�A+�mB`��#�y�/��#!^(9��
.k��aMX��yB�]�h2��XW�Λ\��crK�/�y��#.Bz�0 �>Iz�Ѡ�Q��y��q�̰GD�+�h������y�FܷAjb��p��W�,�l��yB��GB�ٰ��W�},X{�	
��y	��$ �k�o�x��L!ţ �y"�Z3�H��U�p��!	��Ǚ�y��F�yf\����<a�.Q�s���y��A��X�!̆.�r���M%�y��"����֡ۡS)N�!쉃�y�!�o�d�� 9���bbc�/�yҏ��;� (rO���ɳQ*��yrJ��k�H������9���E��y2�W�B���w���d!� �yr!��C�fHaD	�;�
G �y"��8E��Q��҃�������=�y�]�v>j�����_< ��r �y"6S1!�dA�[m��q�EE+�yR��)�\��sfN�j���� LS)�y��ë#��<@���_�LiW�<�y
� ��Yb����4��)��)��|�e"Oi��ֆL>�0���8���"O�L��èyDH�'�!�(Ar"O��a�'ؙ#ڮqh�Ǚ�[_$R�F{��i�4w� ɐ �ָU��ArŌ3!��H=6\s7��_98i�A�s�!�d7J{��4��{���H��!�dՙT� B��ަ'~��h��nf!򄐃!������6�%XG'X�mS!�M�Fx@ds�ĕ8٪Ո4&Z5x7!򄒿Y5��$)ǘ|�.dd؀#5!�DL H�P�	�*��#$��Y�!�Z��ZD	{��9DC�!�$�D:�a��F�B�"��ǳ>�!�D˿+��Qk�)M3,A�T�И}�!��o9�$�cLɜUNdu���k�!򄕜�T�Ѧ��&����*U_!�d18$�\@5*W��4Xjb�6-O!�$A8!{��
e��[�V��ֈդ^�!��[�M� �W�. ���6'M�!��M_Ba�7'�\i��U(�!��.>� ��Ɇ\W\�2��x�!�Q��B42�NA�!"~�!�d�&Y׎����78xZ��ڇvf!�D�]��D��U�"	Q���$/!�76���F�Pw&T�7�U
!��;�$�HW�G;}\��r����!�D�7;���c	�,S4u;`(T*!��m/$��w�!H~e�$�ަ~!��8K�� yA�M1F�,dFL^�!�3F�A�!W�
r��spJ-5�!�䁥[}L��!�L���HE��(+�!�Hsi� H��W�ش�ul�>=W!�$+f	RmSP�W&������_�m�!��:�H�zc��B��8���GO9!�䒇(������ P��3�!�d��Y:�	���'y��8���'2�!��K�Iۘ���K�,p���� �B�@�!����հ�=�%6�P��!����� 
�%���(�K�>�!�D]�O��&G �J�V`�1�!�d�\"F�붏GG��y�2`�4*�!��1��y��I�+�"!p�NY!��-$��8��GnrlhD�<�!�:Rp��`1�ΓFm��Bׄ��4�!�ɀ;r�0X�OU�c�ĩ�VA�.bj!�dǣi�D]	Ao�7�t���L�5^!�߱\R8h 1�B�c��V!���K��y��剅0�*ٙ�A�OL!�����݃�j��+�6CG���!�R�P�LŀW�,��&E�!�d�>�17-
�<r ɘ%��t�!���C�	fE��VO�E �d��ig!�$,F4\R��
(J��ӗ�O�>^!��6P��mq���n5F�97>�!��G!m2�c��� �d`�1rA!�d_n|~�A��j�d�C����4!����*��N�Nm&eY�ɺ\�!�WE���
SΞ�%M�k�`I-L!���'��Qy�R����	{ !�D	$3W&� �K֣A��$��G���!�䄟LHS�ŇC�te�sL��v�!������t�prr�r%M���!��ڲu�f�d �KlFA;�L [�!�� ������%aޱSD�
�����"O����MH�gP��G�Ѥl���"R"OBUZ�!\F������S�?��ț5"O.�1e��X@�8x�׷mb��"O��YUÎ�#�N��FK��_W,��"O�,�	�"1gh�r�	�+e�@A�"O���)�_-�L���N?����"O���Cf�'��i9eH
9.�S2"O��&�H��~��F�c��P�"O����F@�R��9¦B2���B"O���1E<ntąӥ��ղ%"O>d�v�ݧ/�@<�v�E�'.�A�"O����W�=�(�1�熴 Xd��"O�8i�a�V}*WMJ�B��x3""O��3j_l� ��Eӈ.ؐ�SA"O&0�M؋Jv����Y�l�rb"O��1'�	QS~܂ň�;�N��"O����7_�b@��@G��P�"O�L�c���}���k�`-.���0"Oʹ�.�3k(ڠ��G�2�J�"O@<�Ah
�g�����>����w"O�"w/��QY\��-�+�̽�A"O�<#I��'f����Ӟ M��S"Ot�8%� 29쬉��ЙS��U��"O�T�Ӌ�V�� ��H�p=��"OPKc��,}���i�&�UZ
)�"O��#�څ4�9�3E(lG\u��"O�t�#��b�2%e�{�����"OJ�H��G�5�0�a�����"O,����0Ƀd"ͬH/t��S"O�}���ՐXn�:���\��u*O�H��kD�*r̻ ���`�'p�kqd\�����+6�4��	�'�
h��(
�fW a�!�[���	�'���Wd��f���W�=J�:	�'�F��'[�_N�LX��M�]�Y	�'f��0B��;��0j��۵Tݪ�i�'5�E�Z�y`\���F�5���
�'İ��ࡇ j�\�c(�5ΐ�8�'��{WZ x:��3��#�'e�;���Z� ��RQ���' �$C��:�EPGBԞC�d�@�'���q[����	!B`�%oYc�<�pNت�n5LO�Y?��!���`�<i�e['l���˱R|u���cO�]�<����F?h��N�Fx)��Z�<�c'�3�*�����+��]W�<��"��p�`v�ˋv�
���O�T�<1�&Ǐ0X��Fop�0��K�<aԨ�~h��󉍔F/$���jMK�<�U�T�&WZ�!Q@��B���[�<i�8��K�a� ̡����c�<Y�c��1:�g��p����"Ni�<y5EA�4�~% qk_S9Œ"H�I�<���K4�j�{!�/K�!���q�<1$Q-
M�'�V�#�ʬpLj�<�7��{�QL�-���X���l�<Y@��>�oˋQCD�3 ��B�!򤕓DrP�E,<%N�CQ.�$x!�䆹CrZ8�L��d��jk!�ă��%)EǒiT��sl�%pN!򄆎3���B��G�SL��A!�$4}����SmٿC<Z���.�!�dA(!rH�R^,��anW!�� f�y3�dVfi`􌖐w�>�P�"O�nQxd̒�ī	ΰ���"O�|y���	Z�!4�ɖ���"O<X�%K�%ISN�{g��.�2�s"O�hɒo˳c"pD��]'n��"OX�+B��k�ΠC�+��8�t�"OT�1Q���E���3��88�8�"O&��5hĹLul�r��貢"O�qI�鎜/�2Tj��@�j�ҩq�"On��(bt��oěw�T���"O�!q"��	n��#�G?t�$Š�"O���C,�XSV\{�ŭ3��=�D"O��ph��iB�-�U,��k�$h)"O�4�wș!Ke2���k:;����"O°Ƀ�U�2X,�r�@0qc2!3�"O�����ޑ&(�PM�9Z��c&"O68�C
�$�a�p,&�!�"O��3���
���P̆�N#� 6"O��Z��S�W� ؠ���#x%�q"O�{4�O�F#L,��, D�"O\@�̏�+S�1Y��64;��Y�"O	�!i �����ʕ&Uꅂ�"OJ�,[�c<6�S�ӉbBn��T"O�H@6mΡ]"41Jv.7�I�"OL��ޯ#��Xi�ꀌ](@y2"O�	�iհ<��Y�/�un�"O�0Z6`z���Xw���3"ObD8cO^-��J6C'�V��v"O�e���>�M��ـ?^<�E"O����)�c��1@�O�br=��"OT��ڼ2��ٰG��#k��}�"OaЗ㒕U��Q6L b� �8"ONEapf��!�����z���KF"Od��A��<'J,��Ζfz�j�*O|�0AB܋ ���pL�3)rxb
�'x<Dz3
*,Dm��a�D
)h�'r�򒏏Dt��;�����a��'����Kq���	�,O�O���)�'�|��d�:g�(�q��G���
�'юE�4�j��F�<VD�
�'o�1�.��H����ԇB��:	�'����쓄
�J�I�$8:c`���'c\8sO�Q�X!���4�ZMA�'��/۬G:�Q�-����'�Xz$�7/t��U��o5�	z�''�a���/ruJ���"Q
�')<J�L%QE�pa�d������'2vxcr�ىo�$�ݞ6�Y�
�'��ݡR�Ɛ @�Qs�gHZ~	{
�'�@p��x4=���
�En��
�'Rr���1DaZ���; *��
�'�Xy�dh�%!�L4`F 5}H@@R
�'KjI	D.0Zy��)�}�Vu�
�'������R���Q���q/�l	�'p����`D�:fe�D��S�T���'��Q�R`�$t-�4�@#R�4�x��'�Z)q�'%V�z���&ߟd���3�'�,���H�p��{W`�e��'p����!tM�]����c�4A1�'.l=� ���[v�
�ݞ[0���'��X@�ִ*\��B�S���C�'�|�6aM�$C�	u�<^�H`�'2ĩ�ҍ�nJƩ�d)OXҀ��'G0PSN�d�H�(�%>"�~�A	��� �-he�4��d�@OT��5"O@�����J.	�g �kCv�d"O �@���.~&�`���!LMȤ"O�	�E�B�<�q1��y9�"O�D�_<3Xv eQ��\�S"O@��T_�uV}b��5Ϛ�J"O��p4O� w6,���K�$XleR�"O���T_���BiJ�%`�؀v"O(d�/��q�ͲB�L@h�!%"OhYub�<$=@���D�X��"O���%oG2���!�-��"O�P�f�M �<�,�w1�=�"Od����:Rz�Mhg�U$X V��D�x��'z ��'c� �� =��X��d>����X��p�A�Q�����*?D�$��B2[�PR��Ά��i��x��F{��)#�,ͩ�KQ�B� 9�ՠ�?f!�7Knm8�h�>K�:���)M�-<�'��|2��F��B#�^7�f;�	���y3f�d��nʁr���D,�p<I��$W�k�DE+!��*)X�#Ɓ�8P�!��ڧ+�F\�p�E�5"=�MR�Q���hO񟢁YG�C��Ȧ�H�Ȕq3"O�HyvhΑ-�<���Ĺ���s"Oy�A�1>��j��y5��&O��1�,ōf#�Mr�jPac`0D�<��_8#{P7 Ň;��H�$WҦ�'t�܁����@u#x5�ɔ	��E��-,a{��$r�@H�@޺i�K4��B�Oڸ�牓PV���5��*��cp�O2�8C�I�r���&��o�di����kcb�'3a~©��7�p`��'�$�H�!�G��y��ݖ;��q�sKQ?$�(R�[��yҍ�f^l��		)#�F����p>qqɐv�VE��c_�V`(�Q �zX��Dy��>�PIb0�Բ�<�"o���';az�d4] |b�E�l��6�L��ē�hOq�"��$*	i���'� j_����(D�\p����hv^\s	�qW��c�d2D�x��ˬ4n��@4F��M9&`�=,O�,�'߉'j�1��g��PЋ�
}�$�K�'|��QG$�U� �A�A�`�pp��'H�D�C^��Qʣ��-d�50�'qb,2����p�f��cI�:Z.`��'6 Y��*+�u)bo��Ph.�b	�'�F�J%�B(�b�`�Ț{�D���'�B@��iʤ*7�@��C.���'����
���Ȁ ۠�\xu"O<� v��Kx���oD8.K!A�'�<+�_-pq�	9��ܜ�� �=D��y��X�� �R"�g,:E�7=?���ᓪ9gJ�y4��>�>���l��_�C�	�j�cʂ��8�6�2Th�=�ÓX�"\@��_cN�#1�ʸ1�݅ȓs4���sm� ����	7�dE����0 �M>zN���֮{���j���d�-R� A�F�$�.8��O2��ӏ*oAH-�7!�k�D�Y%��#�	R��ON�i.Xo�P��՟���D
Or6-�	93$m�1
Ƶd~xMC�׮"W�'-XqFy��?�$`F�8,�����Մ&��W��84�^��d�k�'7��"Sϟ�&Yh3#A�E������'r�u;��T.`���8b��#�
E��'�8����:�x*7T1C�l\j��n�L��|���� ��JQ��,a��mÓ)�|^����'���C�ĳvQ�(��L�1O�T��c�ODC���H1h�+�E�,�����I˙4�c��Gz�I��+��A;�mV��(`�m��h!�d�%�T��a�݅u�jq�7��I��'�j��	,'� �@��m%���4�S(3Q"�����M[���7U��Y�m�xr箌i�<ңB1\�(�e�<�B�qg�h�';?�;F����	S2KGm� ����3D��z�%�6r�\M��kуr����#�3��hO�S3\���p����r3���u�ݹTw^��%�L��4r aE�`>��gh�5
8��ȓ����U�)a��1!�#<@e�ąȓ^�xɳ5
�r,��`w�˾`��0�	s<q���(<R� .�<k�+n�,��y��	�-X�E v�P��l�R���P[�C�	�ECVH;Ta\�2���X�K^�B���O�=�}���O�y�`�nAy�&�����_�<�》(�AҍS�Iܮ9�׏�W�<A����T���@DFN3grH +Ć�VX�l�O��HP
?Q��ۥ��p�\x"O�Ȱ�9�%��K)gP:,��"O�9��ހi�|���	�B���"O"�;󋇶#C���&$�ٰ=O��=E�4�Wh��@��M>��A!�yb�Ix"���M�D-���L��y� �+@j)I�*��>�\��a#@+�y�"D�%�L���`�;I��y2DWO�8�1�#NX"2������y��N�G���2�ߴK�Q#�N��yb��5{ȝ�"!ٝrqه����hOq��l��j�
�xͪ"N�P�L�)�"O`H�������P��G���d"Oj��Ã�r����FH�U��0�c"O��(6a��&�Նm�<���"Ođ���g|�a ^���"OH��n�*}��EcNԕy��AҗP����	>�����,,�Arj��,b��G{Zw��9�N@*�χ?"���,?6K����i� � t �7�j�1��8��B�	Q�QR�g!]���c��%�B�I8"�Ja�Нv�2U���[�^BB䉰0X+�E�dd�K2��}�LC�I,W���pa�� �N)���p�B��?��e�́yN���猹֖��d-�L�q���
�m��~�Bg��]�!򤐚e:�����j�n`R&B!���E{ʟp�WAL�;������,0��M�"O���'c�kl(���U�9��u�"OqcA*��nA{�M[�{e�p��"O�Xz�i0h&�8sp�l!��Y7n!���=P<=#��*e�#׃J%>PQ�P�'�'U�Qu��nǴH���*$f<²���Oz�O^�/1f�H�&� p�L�xǚ�pF{��)�54Լ�Y2M0?�@bƉ��_���G{ʟ�u���	;���0��m޾
��9��4|O*�ӄ�A>S� 	s�Cb��Hz�
OVE#�Ś�U_p�A �&szN��b��y�#�ObƉ��$��j���0��y�-[ �´��L��(�g���y�KW�2����76h.��6�ن�y��̩o�!��ۗ ����.�?�yQԡ�`�(
���A��~��'��Yq׎]�K�3[4��#�OK��HODO� �Q��ڗp� �R�O�}Ծ��"O�9�j�0Xj�	�kݔ̖���"O$A����}I4�J �l�A�$"O���T$܃)�8��w
� fo�(r"Opu�C"U!
�^�C�f·�hC�"O��bFȷL��$HW�E .t��x�"O�uHE�3&�D��ĳ	M�1�W"O���4�ѫY�b���dI?(��eb"OV�z���;aVD�-�"�b��F"OhuK���egHWD3�NY:�#�k�<�ԭ�A��ت��S�\(�p�/s�!�d����c=.��k��F��!�șz((h���P�N�����T$!�ZUҪ�˱O���݃���:�!�DG�$� 5�񦕓b���cW�h!��>Ίɚ7�וMFPIa��[E!�DƌB�d�&�1*�,{5
�#r.!�dF�pt8�7�^�����.[%=*!���.W�]�A���r xfgPZ�!��B"FޢM2!�8{�*����+#2!���4i�f-Pyܔ��$��'�!��N�nPp�yb�]�w��x!"�<j!�:F	�<��%�;�4pAaJ;)A!�	�+!-N����	W�!���"i�vK_?VɜD�wĘ �!�䜯s�`��&�zi��O�<�!�]13��AFc�J���!Jt�!�$�%P�����oY���ꖀS�l�!�DD5>���P�5{�Y��,@��!�ܬb\$��O�ƨ�E:#}!��^����G_e��d�9P!�dҲ�{��7� �RbDne!���,%¦��<@�� L|!�]�B��EӃ��
#�x��D�~�!���M�pR�-��;�m�g-y�!򄒃gBE�5�ea��=_!�$�aδ�P۲;9���~E!��ڋ)̆��H��I�)JЊT/X!������@"�HPq��?�!��[.�>8��*ל7�T����6|!��w �uyэC�����&^�!���;��10�✼P��Q"�c�!�d��B!�Q�ָ="ԫř?s�!��9C�*�Ã݉O$!@��Z�!�$�5<+ԅ��(��q����8!�$]�Ɇ���yuX�Y�فhR!�d�|�ȡ��֟_m�U[���HN��gl�	?a~�A2F���P�G�-�h(�UT�y��U/:h��i�4.��у�U��yr��X�T�	�i�@�ˍ�y"È5Y��������1@�U��y��߉��i1��,[�@j�����yR���p�0yǏZ�	��r��A�ȓF�)�΄�>E�eH�mh}pl��{f.��I��A �!Pq��^[2!�ȓq���&�3f� MAgn�����ȓ`�ʩ���׎�(s��I��H�ȓi	~9��O�.�F�b�#5�V8�ȓ-��,�dD�:|N��"7Y��u�ȓZr����V�X�H@��^� �Jчȓ,u�=Y�� 8�(��U�c�z��ȓ�e[G�$�����٘�\���

��7�I�d$�;gjښ5�B,��5u�����/n�IA��]�^���S�? �@�BEVeh�P��\?��"OxBr�Ќ+4h���>$@�"O���D�ي$ќ��aB-D'DdKc"O�EICm��X	|�C�Jf�p"OD���1^&�����2i2s"O8��u��7BT����ƪh�@Ő�"O�3T�ҷb��A�������"O�qiKѺ*#:�c�
�h8�"O� !�G�O�@��կ\���Tpu"ORy����n_��R��Q�ᘆ"O�}Z&"
�L],���/�!ߊ0��"O� j�L�c>݂�)�p���if"O�UY�}T��Җ�ͯ7�ma�"O��3�bS�H�u�#o�--��<��"O�i��P�tpg��4<��ܲ�"O�����J�
��d��j,x`0"Ov��oN5W0��V!��%��:�"O�I��-O>X�*�1wa!e�Ra`4"O���q%��[��=	��#"OZ�B��N�~��*�M�3��x��"O�yؗ��`2�p�X�H��4"O��i�ٽjٞT2���&J�y��"O�J���<d�Z`�blE����"O��2�L��6t�4� _�-Pa"O,�k�DO�j��@ѥ*�=s����P"O����>�ڑIPJ��A�haPd"O�<�F�-�q��/n޼���"O�AQ��L�G�ʹ��/���v���"OL�aug�1�Ryi��R&�17"O@y����w:�ң́�Z�.u�5"O��c�ğO}��	��ʑd���zV"O��0E�<j\��3�W%Ia �Z�"O��+U{��ig�Nd�h@"O��W�~� 7`�F����"O���DR'|j��� �i+�<�"O�S�˞)��ma�.��)��� "O,�
!'�e`(�@bؚ�b%җ"Oztc�F�2���.0�j5Z�"O�\��NH�^`l��ޜ-�&�@"Oj����T5��D�w��}*�"OXXs�y��c c,!Y ��"O�X��jN%4
�ʱ��)_��"O�,���É"��"�+Vi2�"O4�Is��2�2�� )i�j�"O���b�	:X��T �!R�A� "Ol	[1��s��@�g�\*�D��"O��;�/Cs]�����
�>�x%"O��hR�6+NH!A�7@x�$i�"Od1��Ε�BТ�VU�cd���yR��?@r>���>�~hA��X�M�h�'79��"~nڔ%�H�r/���ec��ȍA��C�ɍ*�T5a�P񨤂��@���	�P@�%��*Y��zB�'KN%XV/�:/_� Ie�=Y���!��q `�B3O�)��$�:L(��ǣ��y�\L��94���c�����3���x�L�v:�	<u\ a�P-]�~���D�G\�'��9�F�͉o�X�ӌ��t�0�'�\����u�ayrn"��B`䀀U^(�+���ލ��G<� `�U��?�Rm=�')���]� Ŏu�LF�&�-9���3)TT���G(<aA��rCl)g֛X���Kl���W���vyv��Ջ�?u���jq�N.sBPY�'�Y��`�]���:L��)��̚%�@5�2LOxj$�}�����S�?:��2���# ����ܸ�><S�f̭OB8*��	�ڕ�����`哰g����%�A1HϞ%�0��2�x�O�-�`lُ6�l$#f�O\%���	���r��`���6,Xt�tl�,ܢ��'OܤP��Ҳ;�Pl���'��w�߬ j>z$�UO�M9a����R ���bIVpE�����O��0�n���� ���t�O�gU4]� k�$!��0ȈHe�B�I2v���G
	tŒ����(c� N?z���(�Ly>p��a��q���G�I	p��I'��-���w�	R�	ۻ:�����,�Gx�J��>��ٛ&�����5BS�o�F�pa臵��]�0��Y/*M���Ջ�jp�(Yuy�Z?S#�"��鍵T�z��eGM�������3�d������ҍM��t+E/�^z�\#+�9����-_�X�aA.̴\T� %!�=��92�faɗ�U��$�ቼ{�ft�DWS�ڙ���C�����gG4Mb�aU�<c*��૞�z�1�:��0K�~�j��ʐ38��*�Nթ1� �?A-!�$
�N���
[����	��1A�A�$M���I`잛g�Y c��M�䅛p�����=K��ջc쓠,�x;fe��RmR�0=)V�X��B<��mK�?�2��P��,����A�P`���R�� M�AS�O���|��'��!���t���[�F���Y�r�p`�6ȧ�'�tl�f��w�ډ���T�<����oy�h*�O���!�).(� bGH(<���O�Q�Ζ�QyazRI4F{N EK��k��	�r��i��XS�Q��Y���ޱ+�$����L5ǸOXX�;� �����ZnhM��MǾM[����6*���H
Ӣhr��̸o0BU2�`)+3�8�`�ʧeLȀ�&��$6 .��BS�'3%q���+?�����-V� �X�z�ܸɲUD
[�`0Z�n	�~���B�,+��� �Dp��ˁg ,$tՒ��'1<ai��$�H1/ք-�4���C�'dt�bR��M���E=[�|0�b>	)��y9�=ʧo�*����d�#D����E�<@T%ڃ�W-DuB$@�_�T �Cb?a*S���R��9�|8��Nd���u�҂9����"O��K:�A�A�,������򰤑cA݅h�������-�D�؇oF�L�"0����tl��3(���ѡLF'F���@wX\4��E�-A��mQ�ۊ�y�o�p��\� �Jj�h��bM��'�Z�9�(�[��EE��R9d���Y�D�7���y�ԗy��#��av����+*�@U`'��,=�'V�>�IlAQEm��7�z�V��9PB��Z�H�&K��c�|��RG�42����k�lxY�*	��=ɳЅ0%xL��H�=Y��`d�R|��г�a�C\8�듼id��Js�kr`,��Z��h��'����W�ߏ@ B��E��^�`t�«^�-�:5��\���:��i�.4*�z�*Ҽ-�z5����
�!�φ`<�a���p=8V��a��d(�����,�ɰ���a�j��s��@"�U*�JI����i�z�E D�d�� �!RJ���T���Id�ö�?��Dp�H]��HGP2�3�;A�y�OL(`?z\bꅶ��t���9G�Qa��?K0��YA���u�ΰ�6�c�(�$�'l
�ڦNz��-Y0�ȴWp 0��$ۻ;+������ħLJ��� "h[ ċ%�
��q�ȓ&�� ˗���NParpꔃ;j (�'�0)E)��V	䠥OQ>qZ���R�ԭP7���j%D��Y"ꛦj�ڑ�#�ҦM���+r�ƛ��%O�l�����L�3�	_T�ܪ�O�;Q ̔��B��N���\\���'Z�B��2�l�`e~%��hB�Nr�U8� j�-��)	[�:��U�
D��æ'ob!�ת�w���K��K�f�;ӳೳ�<D��W�F0ZHrHB�� �>�D)�n??����@xH�8J>E�DmI']�L��c^o*({�Dۖ�yb�;y��е*�L�rD��''`�!Nv��CaP2Wf��FfeօaRk9D��i�핐T�*�P�/W> V���w�4D���"jO�eEl��@��"qd��b$D�h˔�T��a����7G@R�#D����l֩wߘ| UoDC��:D��Q�)NyB���O����@9D����_%g�ڙys,B*�p�рa8D���A˅ t��C1��5�(�"*7D��x�4g(�9��ά)��ٔ�5D���*�j����%S���"J2D��	��*W�){�(�ު 밄2D���V���V(� 	���0g�8{��-D��	"� Nr�� ��\�	v��A��-D�� zT0�NcJ(`
"��P/v��"OB%{t&۞Bޜ��Mɐ��ʂ"O\M�Ħ��$:l���V*��8�"O�pb������@#���C"O��9u��_eZ}�%U���3�"O�дm��n���Bf.A�HX�`�F"O�=�&#����dh��L�9�y�a"O�;�fŢ]�U3��p�tԂS"O�0P��;r��@@ō�\u ��"OZ`Ф��\1$�x��Cn��@Pu"O8����Y�)�����S���R�"O�X��;q�<�itI�t6`8W"OʍB�LI�ry�pX%hK�X� ��1"O���E�R�N4�����-'��˰"O���f�E�!b𣔢ZXw��+�'6���� Λ,���UIGgB��'͐�3a�0�*�b	^!�,(�'����nG; �8e��
6���
�'BȔi��[�q�#����
�'� ��H�+�R/�Hr
�'IDQ�+�+"c�)�A�ۼ	�B��'�X��肎.oƐ ��Tu��e��'�(�IhH=#K�B�K0d�Z�z�'�0a��HQ�H���N��P#�'��r0�DPt�aP:����'{�ظF�Ϯ(�����6���P	�'�PE9�-��2i0l[s̗;.� ���'��+Ԁ��.<vl#e��i�����'������%a��Cm��uab��'����p�9b�H�  q5!��'���x�^2<��C��]?i:N��'=F���Z�UlЩ�t�ԏ4����'��r�J��\�����<$���K�'��!a )S���� �'wM^pK�'�R=�F�>�dbC+pp|���'��N�,U�](ӻ}Y|� �'��ԁPf��\}|���Cːg`����'Ԃ�� ���[���OA�/���'7*|���81W�c���ch`��'�H9j8U��E
[�+�ҥ9�'�(\� ��$l6�  @�3S�D��'a��&�D��-b���%A�L��'�b�� v\���kEt���'�!��fu0��Р�՚D����'!D)�� ����x1��5k�<P��'���`A�E����Ԕ*� s
�'^RP�c�վ3�&ɨ�T���H	�'�H0r�L��Nv���9p�LQ��'��j�"�%��l���[H��Q�'U8����\+Uc�EY�0訑�'�<1�Pn�*F���EjJ0q����'�I
���{�~q���v�B	�'s��N ��T�G��䤳�'���kd���&����F��?Q 	@�'�T��F��N�b� ��)���S�'-D|��C?c�y5� v�B��
�'���;@�=&��#+�f����'F���b�E=��,��`� E%�'��0��eN1�R1�a�4	��'xia��F��8A!���31���'��D��ɦ`�ݐ����{
.u��'�0��sEʸaW� q�p�@	�'� PZa[�1���hΌ
u��@��'z�:RfN�a׸����*2�F�y��� ���eË�s�F5��o|N�`�"O�Y��dȺMz�x�jՊa\	�&"O��K��Y��C��4��5"O���.aU�I�C�W1�`h�"O�Qi� TJx�H!�U�(x��b"O���"���|H����8/��y�"Otq�G�0e���
 )��(�ks"O���2D� D�Dc8		d"Op-�@�V��-9$f 9fS (�"O�M�—',j�FW� N��a"O�Tؒb۔v�1��F�V1��x�"OXU"�c@+u�t%���Q�D/Ja��"OpL�t�� Q
f����\�s&t���"Oq�p-"`V�1�7Å��v"O�q"& �'�dʔMQ'B���"O�p;�
B>�ɱ�M�4�LI�"O>q(2�T�
+�!�lCe�l��"OH��(98��q��
�UL��"O��u�%n$�h�aF�6��L*�"O�� ���=OV�8�N�Q�2I�"OTDY��:V�%x��݈y�j�:�"O�P!�b�.\����k �Rs$�x@"O" q���;P*���aQ�9R��"O��P�aRL�A���vN�L�3"O-CQ�)t�$�G���a�I�A"O�|�����5V�f�8��"O4�@�,�_�\��@���@��@�<i��:u!�|#��&|xST�G�<���J����� �:�k șn�<�"	��q>��&��\��U�Ow�<1fN��ts�U

� ����m�<ٱ�	�Th��xPP~]��@�h�<�e�аo/�PHӏ˅* 삆�A�<A#�_�A�Po5��E���}�<Y��Eo��c3�ܭ5�fEjG��{�<a�J�|��]�CgF%}�8£�[z�<Y0�f#��2����y2n�z�<��?w0:H*��'`@XQ�x�<���Ţ.�jP���ע;�F�itnp�<��*H��@��]�=���X�)Xn�<��-5\�IRҚK� ��M�<�n� &�
4��a.�����U�<��U*ʬ��l��8�t����PT�<!%iP-cD�Uñ��^���P�ÁJ�<��$?W��BF��$O8��gj�G�<��'�7�lm�0��fݴD����A�<���I��i�'�
�O|�e��A�<�j�XX�Ir�'X;=,臋B�<�	׶~I,Q�	���q��Xy�<Ywf�#}\0y��I�;�b(�#�L�<�`��L�z���B�Ԕ�	�' jAr��+hbH��[2<(�	�'Ux`Aⅲ]�a��j�	j�	��'	������!���˭��p�'vI���ͬ�4�S@g��w"|��'�v1ӑ,�^�4;�-O�����'dfM�#I�Fs����KHٔĆ�"��M�F��$�̊�/	��`��(̩���
���C"L����ȓ.��yT���.$qUfź��$$� au&E��ay�쐘O����d����D�5���?�wΙ�3�"i*6DN73����1,۳T����W�&�Px�[	~��{	��d��2�m��'��\�E�[ �q;���qH,5 ��>��h�48X�MF3�z%�(3jt��dX��}� �`�w�O�����3�����J'}"p��ā����s������W�zey�lȂA��!���>y��D�p)� ���F��!�
,����NO�j����'Q�X�sN8;a��2��'"ne����&[�ԉn |���q��O�|�%�;�$ț�/���O���1c�.����n����A@&L%q���m�x�!��A5�m�fAж)8�:�O�;	���9t�O�Y���Ѫx��yxV��׮UӀ�۔��y�ɛ�K(�p��դD�R��;5�O�Ux��ϟ(Ǌf�Ы:��c ��h����,	�f�
��s!O+9���.O�q��.��3D�����nP<�����2X��(F}�)�.?�~Q�̲~�!�5X?ݸ4�4��yL�aZdI6�<��2W�-P�Y<�0<�U��MPt��#K�Z�v��%O�_?���\�
�r�/z7��G�	�,z:����ŧ\8Ɣ�A�?a��y2�±t	lڕ
O�l�JF������KG���J7m�h��qˈ�ذI��@(	��x�ƪ�
����OT�]lr�}���W!R��EJ��Wn����M�(��<��JG:J�n�f�U*n]J���m�~���)�j��֝|��S�d� �Z��TK�u����3�4������O�=�WnR/�fT���߂8I��axb�T�Q2a��ʰm����'�4Tٵ!�P���1��;�p����
�f/�P�*��3h<p���Y#�?]�!N?�i,��:�� ��7D�`��Eдq� �pda��~�~I�Ӈ��~Ve#�O"}R�f����,d��U
��D2D����'�X�!�$�zzR���� ���1��h>�H��'T�,Ę��'a�Kʐr��,�t��
��l���dM=c���'Sd��h�^o2�ͧGs�����ڽky
u��G�:t����-e�d�0��|0�ݱ�㖗��<�r��	T���'���0�G��3kQ>�ݵ(�Yj�C�'�@(�C7�4B�I'2�V��2�M�p��L���]Z|2#�/��3�HN��~��O��xEzoV.]����.a^�a4AO/��=1P&�C��@/v�h� �BJ��)�׏�w~��[G"OPx��[�1x�4`��hp�]A��DN>(⠑��&Ƕ�H�����L�`'��"�Lաgg2�;�"O��y�i?�<є,7gV�(Ủ���Ѡ��AS��8�g?���-
?<djRn.vs<I�&Z�<�I�� |�L�!�Ŧu{��@a�Ο� �Ġ�Npr��'��5"ٸ��3��;�\���:�$���7M8t���+[&�f�R7D�/�!�	a�eRc�Dq���ď�F��O��Y�����<,Ä���+�<b>�R��X�:�@��j��<Hc�?D��iP�C�E4%x@g�$�U�@�ܞ�4pr�p����՟"~����8�� #3������[����y�~ R��:Y�q�Wc�]�.D���'4���5�[�|0�d�,EF{R�K'wh�i�͟2qy��B�#	��?IK%r� )q%k8h�X�3����f��CL�T����D@C����2����ՌWџt CN�4[�PC��$��42LP�f��`�t��5�R��y"*P��d�� A�a-<�ҤH���½S��XP@���)�'s���س���)�@�J� �XJ��ȓA�.�k�`�9G��3�N�V�!2�>9$�ڟl	��{L~�=�F!Ӱ�n-�Њ�"m'Ny�5�Dc��<�&!R2E� �9#-�YeA_�b��]��� 2�aB�P2���yD/�m���"�C���O~��F�<CX���J|Z���">���.V.o�NA���<��`T�Z��`��I�/c�(��w~���"Z��A0�|��	�j�Ѕ¶�I�dC ��r���!�DÀd��3-� k1ʀ`Mƃ�qOB������0<9��)��!S�W�mn@M�q�t�<�k�%Xv�{�n�QL8)P��m�<Y3�xƦ85Ã� �Pf�S�<�bȁ�|'P�$[-O�f�`(�L�<�-�ch`r�	%a'���q�I�<!�@��i�f(�N�E��e���J�<��(�Zb�A+ ^��u�M�S�<�ā�<f3���j�vx8PLN�<	��=T���.�R�|]B�IKN�<� @����,h1���
A�<z���R"O6�Ȱ�Ly�0�b�H�ZF���"O�╢C�+ ��C����мx1"OıA ��}}�]{����t@�@"O���j0C�)j�J��^0ݸa"O>uِ�мp�t#�8WN����"O�rҊֻ$�X�3 �"$�IY�"O�X@TT���R5I�Q�"O.ؒ�鈉X�Bػ��Cl�A��"O>��DU*�ip�,%+n�]��"O)PBgQ�?m8a��ϥ:R�"OfX˄gU�o1H-z�
R32Z$[�"Oh��&��>&�$F�*KJ���s"Ov��e�Ӂx��8�FW�xMv�[d"O����$�%&h)�ˍ�^RT�!"Ova�
X�G%n��JIL��Q"O�0W�\�'p^��2�؋n6(�'"O���'�ˌb:���%�CH���v"O����+�~H����T"�>���"O"�83���L��!�@Υz�<�9�"O,� P@R+3�@=�A�X�Q�t(d"O"���f֙mW��#�C ���B"O�s�c�=5����A�V��X�1"Oܐj�;����BA yc�]2�"O����_1����R�4K��ؔ"O6Gjɬ��-{� �?9��z�"O����(ɔ���Eծ_ 4!5"O��"I4e��1Wb���BX��"O(���N�^O����τ���(�4"O���N�T��!!�c���"O��Z�(ۑ=p�qt�	�<��"O�9R#͝-�v�)T�5�@h�E"O4!�%#٘#�i�N�7#V�j�"O&��c��-ct*<B�MS�I�b�"Oph�E���;uF��ɏ#���"O���O�*��P�B(X���x@�"O��Q5%�\
�M���O^���P"O�E��n�F�3���u��"O�qh��Z�A֩�.I���bt"O}x�a�N���#�H�N�4���"Ob����[t���ǩְwl���"O �]� �B�';H\Ɉ�"O����#C�	V$��\{M�=C!"OJ�8��,gj���'�(�8y1�"O| ��� �0�q��R�es1"Od��f���bٳ��ײE���#"O����N)v�>I��$ƃ6u��E"O*��쒃l�(<��� 5�>Y�"OF��r�В��ZU"H�)�<=��"O�<� �"�L)x�"D�3�z��r"O6Ax��ފ	1��iu��-3�:D!"OZ�*Gc��7�������D�+�"O� $�%*J@���V�y��"O<�����r�nQ����	_��}2�"O�ݱ��O�10Z�sy^��!J�!rŁ��'/8�8�%R2'�j9akЛ����'9��*!`�u쨩��	�?@��'@Ȱ#�h��R���Cpl�$���:�'�p1rn��2˖ cAÄ�L9�
�'�8h��.��#Q�t:�J���Ek
�'T�)S��,T7bY�@ņ3a9 Dy�'�4)d�����d7V[ni���Y^> ۴��}	�Ά<C��sE͈�2����<QM��0��ȇ��[E`�cs�J�N��Y�!8���	�)S�dR0���	��'��� ���@�����!IdJ����0S��	 jۑ,�V ���0|��Xu� �"A�Z-��R$`�)��U��	!?%��#���iO�Zo�K6��$ܔp�N@�E7����F\q}�&��w2<�	ç{䵢�i�0rPa��\�E�^���P�H`��.r��[��O���{&ǈ+��{vnU=�Pe��'BtH��޲q�� �Z�b>˓*��� C67����'�f� \�Rj�	4�pS��������.�J��h��9ڀ�pԇ^Jp	��)�c���'Mw��>�#��
��&y	�b��!<
�����i~���l�S���5h0Z>�rd��9�&(���Pf����V(E�h���킓+�(()%]�3f��	H�j%��r��(����V�\�����,U���җ�ٚy�hU��Oa�E��E�=(T���7��S�^�k_�=���=�ic�������'�U��H�#���b��*���!�Y�
����_1(�Hx��A��?EE��l�=y�ɂF��Od`��Y���Ӈ�-jɧ0|��$y���$�A"8����g.@)m�2k
�f�p�j���D�$���\�D?��ȓk�Xkq��Ә�A�z�.L��Ln�  @�?�   �	  �  �  �  V(  z1  ]<  hG  uR  �]  �h  .t  �  ��  �  �  ʤ  {�  Ҵ  {�  ��  "�  c�  ��  ��  B�  ��  ��  #�  ��   ~ �  _ �% h, �2 9 H? �E L XR �X �_ f Ul �v �~ � �� � F� �� ʩ � J�  x�y�C˸��%�RhO5d��p��'l(�I�By��@0�'�F��L��|�t���pd��46���jɿ���si��w�D�K2��I��99��ӻ8r��"��u'B�]��T�	�~����Ȳy$�2�]�zo�M����;|���� !cr��;��[Z���3�1��ݞB����M����'y��dT@F�){<��e��$�ZRD���	�*�&!P����Dڞ:��7�^3�Z���O����O��D٣[怵9�(_��k��p�����?����?i-O���?a���?Y7k�"��lȲ�1BX
  �fҡ�?1��%�'�B�'�H(��O���,3e�Sgg� ��(d���prC�I2e�Z|���	�*�"PYuj�� ��D�d-Se��**X���%�~R¤ƗLEzv�I6�$	�@��ə0#
9�4��Iѡ;���',��'��'���'�O���1���,�� ]B,~���'��7�ܦ!��46/�	 �Mc�O��Fd�>q��L;�x;Qm�+-ʡ�ە�hO�D��LǮiX�P+\��\�x'�ј��<����_<̣�mN-i1���爚FQ��)�' �%uG���,���û�>� +OP��D�=j�����o c���6��oDџ��'1�f)�K"d����Βo�XH��'ў"~��$�-Z���ng#�� �n��hO���@�?u���6�F��5J?R�%h���O��O���"�3}RD<��M3��ġX>��d�>�y�&Q��*\���G�>xx���y"2�F�:�k��CR0$� �D,�y"��;au.��B��3b�-I@�V���?���'R��N ��xR��	{d����d@>k�?Q!�]2~��j[U��Av�S����IT������(h��Z�&0�(��e(D�A`�ڱGZ�-c# �(Tt���+,D�<8��q�(
���
F��@�T�*D����*��Q+7/�'LV\!��*��U�>]�4"�+p��ĳSj&&�|3bF�O<E���i>�������'�d�{ӌ��Ÿ�%չS��U�	�'�9K 3H�v4��9L���'��#$��YT����IS&A����'��x;У��d2<KuL�.o9T���'9��p��A}6�C �
��(<x+O
 Fz��I�j .�R�I\�����5a�4/��I�6����ܟT&��>HPÄ%��VQ�G/r!��"ԋ�y�iA9o����@�[�`��*Q䉁�y���?TP�w�z@\Y���yBi�> �!�Ǌ�W�
)�Gˆ�y2�P!D�f�#S�Y,AX�Y{��$��>��OҔ �-�馹���$SR�<�`����ޡ�}��_���'�"�'����-.n��D�$ɥo�HeѕExr<'�-�ax"�5��䱈y��T�ȱX� �`O�(��:�0<iW�Eݟ�����I�h����n]�6��w��7+�.��'w���n�z4��)��.�h��1K�2���D���,S!�/nP��� �_J�����O(ʓu�������y�'qF܊�Y�p~��1�������V�'⡟'+H�]*�{��)��?V��v�٠f�D�5�3��#{��D�E�ᓒxr��@N҈�4��A��3X�H�!,%���X$?e�|��� [�tQ��81�}x��EC���T��ɖI}�d�Q)�'<��ihsB΁T��?!d�0i�	0l߰h���D(Ҏo��~y~�I���)�Ñ�?!���P��^yB(�Wn�p�aU i�ұ�5j�c.�'�T5hf�'�Bd�g�V�2��?�d�!qH�0T���7a&lHօA�g�Xmn�1��'
�\�Bި-j����"��ēy7���'5剞HH
ո�'W��UJ��M�fT\���I���':�1㥠 o"
=����(7l(��S����4,�6�|�O��tV��HV	
�f���DǪ 8B��v�!dؒ�؟���ßX&��O�n�
Rl�T��;�ϐ2IZT ��/�x"��f��=AqMY!=Q��dϜ%�"���'��=aQ	��/e�9��θ>fL�wb�.�?�	�'`�pc�U�Z����e�ĳ�'���a��=c̜�e+�3b�$��I>A��i��'���c��~r�븐��#D�oR��1�PG�����d�OX�$o>��Bɀ"�A�OX�Y�.�)� �K!��.�`���a�'O�L��f�'�@�8�%I'8|]��*�2�B(�X�x�dP�S������#�0<��*����	]~�N�v��LR�)U=�Via6*�����?�ӓ R�!��GB6W�@�ӲA6{�����4�?����d�x1b�C���~,������'9R���L~��
��Ov��M{��Zپ�ء�K6NDˡ@�\!�ԁ���?at�]-+f��v$O�tP�Q���	7"@�M1�926��45ʬ"���x~R	B�s�!&�ϱF��@R�3~r����ReX Q����1<�V�ɰ�	ҟ<G���'-"Y"���?`q�ֆ�.v�(s"O��b��K(	 ��q�GU�4������h��(�c����� VR@�/o�2렏�Ov�d[�!���m��?��	۟,�'��5�s���1o��p׈�7S���MP��F݉@�O��6� �1�1O�`�޴\��
��P;�*ܜ8���d+��?I[*v-�#�3�	�z>��bDƇ�S�y�t(ևr���$5?����(������?if�U�"����a��q�����L@B䉗8��0��r���1mZ=hʓ=đ�B�O ˓lL��c��F�3F�yV.ƹD�`�8�b$DțV��I���'��I��T�	�|R#��:"I�C�[���M#w����뚘3�x����I��A��#8�p��A�Q�w��0�K͇spa~���9'�ػ�iE�xM8���x������?����?�/O��8�I#QR*�1��Y�+#�E�)F!$���ca�TRѠ�"�>d�W
1�&��8ش�?AN>1��U����:/�]�$f����H��M�� e�x��q��ӟ���O�-8D�Щk!����Ί�u`�}��"O��犑f�(�%͆?x��9C6"O�T:ge׽T���!%�ƭJ��=�"O��uM��w�� ��"�u��'�|�D
k��T5v�H5a��b]ў��sk=�'5�\ӄ�5��(@�'��H����?��ln\<ف��=1���	@���v؇�*>�9B'K�i�������,�Շȓe�iשK��H�@�	�p��ȓ%vԕ�f��#k��)@cBS�F��$�'R�8�9&��_�ZH�K@> E��%͞"<ͧ�?1����B)�$��d\&��b�O{!��n��y�m�7:qȑ��^�D�!�$G:u� ���
i �j�Q!,!��K� |�T��ES7f7Dp��D��!���E�4�嚏����	ÿ4�	)�HOQ>m���C�n�����,$��Y����<!���?�����S�'1��G�
�����M�}L�Q��~���c���ڝ�r�2-�H��W��ٸs��t�4W&`�v ��r΍��O&���t��c��%�ȓ*����ӣ㌼��$�CZ��&�@z����R��WB�$���
2w@���kI�c,"�|��'L��3(�)�!B�<N2�(��XւɄȓyHLy8G.�2v܈��e�^h�!��r�D���]�hf���0jǐ#�`�ȓ�Ap��#��Z6�Z�����0�?��eӴ�^\c#o�0:�0EaT�'��"��I�r�d�)רHK��1��A�#[��D�OR����5�bU�/e~i#�l?դ���v�$�8��]V����.nY���6��p�Cf�2eZ��k���ȓ:$�H���	=�vTbtc��<�z�F��6ڧ ���3��Q�q�7���T�	��N�$"<ͧ�?������g���#�)[b��9�ӫ	R�!��+�"������H�� �jQ�!�Ğ�U� �Q�[�$X��X�~�!�D�� Ǣ8��ή�J��<�!��Бhj%#i_�~�(�B�U���I�HOQ>�Ӄ O0��3�N�4\�^8ȣ��<� ���?y����Sܧ-��t.��j��4xBBמy��S�? h�+sa�Z2l���'I� �"O�[àϡ"��YP��U�j�"OB\wGP�ӑo�<�)�"O� aj33���b�AB�?��#W�|B�=�{$6l�sӂ%�B@N�>\ ��C��9)���If������O\��T��,��R�^m�� Q"OR���M�GF �!@abF31"O�e����}2�xp� a�J��v"O���q��+|_ꍢ �Y'8K �� �'�R�D�z�q
�*S1{��xsD�{fўd*sO!�'����5 ƪO�Q"'�Ch]���?i	�gl���	�e�	��"E�W��ȓ-%t��$!"O0�xB$cBx����ȓt���� ��~(��)@K��ȓQ�tp5+Ӧy���c@��2���D".*ڧaJ������.l��� w���	C��#<�'�?������K�w�hx5�X?��(�C b!�䊫 ��a�
L���E�E��!���ML�y
$����tJCgP-�!��Y�;ָ��fݧ.�z���À�8�!��P�
���T�in��ǡ[�I��2�HOQ>m�E�ƒxJ��%͍$j��:�,�<�"�[(�?�����S�'3%���sƉ�.�T�R��/��`�ȓL��tkՕvnź���4itp����jũG�$�\�q���)*4��I�|�2%�״GJ-R��B�*���a9�%�s?*KpHbm@2u�X$������F+S�D�ac~�11-I8]M*x#���6b2�|��'��%Ӿ�H���-+[6h#��,vi�̇ȓF0�H��7�浱�C���ȓI,�q�3&̥tj��(E� �N8�P�ȓO��p5�7]�� s�lܠ����?q�*@��jt �������%
;ў�G�?�'x��T�E!��nt��/�Vl����?��Y���1��ݧLA��W�N4�"q���d��얞.R¤�X��<��'�1���A~l��g����]�ȓN4�Y�mύ,r����Q��G��6�'woF��
s�ʝh�C��,h��ɿ�"<ͧ�?9������/��#�Y�O����2�C1�!���h����)����.�pp!��W6���0C�LLF@hZ!kh!���.|3���>tܞ��A�j�!�I��,�BweV�N��+�iӰy��	*�HOQ>��6[�h��HIc��_�dS���<���R6�?�����S�'���  J2~��"*  d
�Յ� $bD�WM�t|���V�aĬ��[��̪�e^�!��i�$-2k�=��)2����˔<�nL2$E׫]��D�ȓ<@)���	<\F�y�.�t��a&� �����4 �D�vo��*H�a���b�U�3H�|r�'(�����*�H_!6���g���x=��5���R �0�� A�P:'�r|�ȓy�(�U��'�J�:� R(\L�ȓm_\Py&؊rܦP0��\����	�?��%B6K�:�lƕ}3�0x��d�'mL�r��	/;�DԱ � ����fkK&@+��D�O(��ė��v�0��@ѐ1"G�S�.�!�Ě81��P�<m:����eI!�HxP͓�C�K8�r���w8!�d�)4��@ȕ�$�1C�'	!џ09��i
�v@�,{�X.��|�4��I,�k�O���O�d<?Yu�	:ݎTYX�
����]�<�A W	e����J�)8��+E�S�<� �`��wZ��
��y�t�"�"Ob�:��'�~ AC'�z:��#"O0����~ĸ�B�ㆀrp]�\�����=)�1��e �L?�ŋe	K�(�2�~�� ���?IL>�}.]N�\3e��)i�x��E��z�HB�	�xm@Ifʃ*A>1�De$i��C�ɢLd  P�.܁�
����C䉝MP�`���%6���0TH� ��C�� p�:��QLӤ
� ��d��O�8G~��[��~"�B�D�i�W�f�x)�ק��?�L>������	6.��Э�M�$����#�LQ��'�,�,A�,ņL�7l_�C�>Pa�'�>�2�'AAqZ���*rvx�'Y�L�-�<~x`@h�;�X�J���K��Н�!���yv
��Cˆ�hO|� ���[�+�����	p�V �	�8��I( Ҍi
�!	.{� :�N�5�C�ɳ5V �r.�(+��	�� �-��C�	�d�1�
���8A��@V�B��+� SEKƱ
Ӱt���/n���?�퓍q�z`�v	���O)0���'�N�@��4���d�O�=�z��n��+`4LX&>&���^��,�Ŭ]�%4����<_�=�ȓ(�a��\H��X�B�פ=/��ȓ(�v�s�l%c�x���ǐ�"�f��ȓ5��F蛷E؃&G)�0��'!�"=E��gE?:���Ȕ+G+(�����ׅ��ČcR����OJ�Oq��y�֏@2�ɔD S�A��"O���,ޣY����7�n���"Omq��9��R�AN3JŮUA�"OV�jA�V�%*�e�F*�>�����"O�]�wmB�Z+�,0G�!�҅!��|��8�(<�� �T�1%E��Zo��avN�c��]�	Y�I����O
y���2��sp+ױ�)+Q"OjDq0��C}�=��V�<�KW"O��
�;4�E�U��#ko:0cw"O��T�� k�-��AY�4l�AT�'��Ē��~��Q"��-�ع���Uў�JS�<�i����-��gTd�S hL̜����?�	�
��P̝_H@7ƈ�o���ȓCX��֎՞0�<��@dR�j���Pyp����<�Z�4o�0/�ЅȓO|�yc���#Z����dW/a��!Db.ڧy9R����wt(y�Ef�b�h��	��&#<�'�?������ԑ�����Dj��@P��>X�!���0P �#�W�Q�H�*0��5&!���1�B��I�:*"�� ��J!!�Ę~�̲�j�]�"5x���F!���0zȦ���ϊ)�2��g"��	��HOQ>����47��0��&O���!�M�<	q,$�?����S�'`� ��;{��A���.}�8Ʌ�Q�&�A���.�椉тJ�c�$���a�U[�#Ԯ��BA
[��Q�ȓmR`�Ԥ*%��ÒnI S���ȓdq�B�M4a� �����}��$�0���Vy��dѣ �|���b�)m���✿-G2�|��''��8�f�9p)ĳ�B�b��S�N����ȓ/~�<�D#¿4R�y�*�*f~<��@F4�t �n����3�.���\
��#��||rU�F4N�>��I��?�c��8~��w��\c�kt&�P�'�����I�#��+�	E�?c.%z�āq�����Op���^;h���� �&*P4��O
�y�!�䄯g@�3&/UF��B�^$L�!�� ƍj���?l�hE/�/	H��Q�"O�<���/[B�H�n2��2���=�h�����ԗ[[p[�/�o��H���'2��B��4���d�O��7�rl1���V��#f�@�9�ȓF/@�{w���I
�y[�E� A��)�ȓ>C"}�����4-R 7g��Ć���B
?$�Yi������@�5D�43LQ�O�J������&o�<���)�'*�ґ!CA�(/V�;�KQ�Jl1�'\Bͣ��'%|���%�adBaS�_�����%Ӧ�yB�_x�`��f��P�])���<�y�̈́�;��h��F�v����yBi�J&d=Q@lR2Us!��y�+�(t
,Ic� �$���ҥEG���[p��)UL��j��X�NH�r'�]r���O�ґ|r�'���c*H�x�d�*f�Y:łͰ}	���2��8j�iR>Ml�<Z3䔬 P����6���$Ǒ?�2��7JU.A��E��jPD8RFXp7ёt���1��|��	��?����{"�H�b �">���%(Xs�'2�����Ɇ�{�H$���_+k��(�F������O����M|L�;4�°OZ ��&�̊sW!��[&3r�8pt㇟pYP�KG%H�:!��?!��q�Nˋ72�
,L!�d�'�Z �'�"l!�D9&��[�џ�����/dnx���? T�q妚+`�	Y(�O�	�O���/?a��A�a���i"�
<FV(�Yq�|�<Q�HU �0E�6�D�u�v�<�,�&��1���5# 1z΄F�<�]@	[��F�S��Pbf hR�!������CUJO���r,Zdkp��'��"=E�Ă�G�,9��đz��e�'a��2qO0��'TnYx���G�$�b� ����x��`(���V��'���'����1�[pu�YɅ���4�����Ϛ�~��m8
�^�L��5�I�f"����դ��ŸS�Qp��6yTTl����H�H�
W���O���&�'A2�iMpG̡T��G{��#"d�p��]����&/���Z���POK��q!%�OD�'A�{ׯ��Xc+�t}��B-O>XPT3O��6�s����#�J-��1a��	dA�"I���ɦ&(�c�`�`�`#QBW��?E��
��Ba�
%(�HY�A��yR��+Vt��᎐�-�45 ���'p� �2�H�i�����E�g��ɭ"h���O>�S�K~��!]�Q�	�A� �Ɲ�y���"�5+^�iS�
%�hO^D���*�"USB�P�)��!��o���'"*K�?c�6��Ol���Ob˓�?1�"H�i��ʷ@����V���sȡ��	�>0p�B�j��_��˟����J_3.��Z��3iN�t�&��"}�n�b��>[����|���g�'�h�35	�:����`X�:p���O�����?A���y�|h�@��u�؀)���kh�UR�!9D����ϟw!�����,wT�����OFz�O{rS�4!��eET�xR��i��%��'�:W��yZ޴e��8��?�/O����O瓿z��Z���2c���� ��%�% "G@G$�2��8��{�ҙ��OZ�óO"fa�ڑ��7r-8�m�$TE)�3膩>�2\�����%�
�G~�(I�?Q��@�w�Z��ŦG����񆛾�?ً�$/�DL���)��)����B�R�ȓ>2�|j�%HEMRt�d�Ks:1�'��6��O�ʓ,s�D�i�����'t�"t��]F�pE��+ϛy�ݖ'e��'r
O'$h�q{�@�1x9(E�F�O�I�'<�LH��Ѡ6�Iq��	}����eʋ?iƥ�g�+Ih�O���u��4�$�R�� +�p����d߷@���'1���� (�.'�P	g"�#R�mq�_���	I����G22����mA+}��إO?�O|�'p��&U�^n��v�n��ԬTj�sgdh9���O���
Z*�[V�-xj6��	�/	(�O�)�$f��NmJ��fW�^��h"O扑��	�m
E$U1"���J�"O� ����1U��!��؊ ����"OZ�Q���L�J��c�ɕaat�1�� ��|y#���<a㮙{d�U=4,Nha� H��O��)�O��,�	w�:)�$ �,��d�Eę?��C�	d�B��&×a���eMA�1�C� c�p�j&�@�2W��x���0{�C�	�Lq�I�`�x��]z�rC�+i�����N����>�_������	Vn�J㇓�?�<@�v��O���i�O���!��6.B����$q4%����C�ɥkBi���?���$�,EO�B�	�#7dd�P"�@�ڂ�1tC��58���q"����HI3�4"tC�ɛw��y#�է'�@H��#d�V�)`�O�0� Jئizg�Hȟ�ϧ8��i�C�Fc���t��]|��'Y��'BIĪIh�s#6�4�L��	�~0zM33hҖJ� x��I�	�r�@��r�'Z�SWꊉ'�L)��F�e�8G|�oK��?��?i����oŶA�١�!~cM�&����?��������uI3�B���#�a/1IN�G�%�O��'.L��Y���	���M��<@,O��O0�d>��f~�CJ�CK�Z;�u��X� X����I���?�r���M�]�e�/���v��M{M<) �7��I�D�Je�	*kzX���ѝ�~�TV�Đ��S��'��M* *F�"pxH��>mʄ�!��;�	5��Iqt�'���J\d�ˎ{B��b"+W5b־�3!�%��I/�~��s��0�٤�%៎sR�i4�9?�Q&�>QC�>�tUJ�D\P�4h�*h��qǃ�&0?h��L��?�f �b�����?A'ƈ�7Z��E��{��i�����T;�A*}b!0}�0{K��sܴ%Y�Z�%�*e��ԧ��h�~��'�l��M�	��	MbVxy��G�w�X)�Z>i�<��3�@�O�s� �$4?�bi��,"6�`�kS!��KD����*OH� ���|y�铞?Z�ّ��$$e*Htg�~�D����~2	A����?�	�Y�t�	�IF���ϝb*��X��\z�ĔӰ?�6(�kQb��(غ�69�iI�<)����=�Tx�*4Ls�|�D�I�����˟��'J�맖��M�mQ6��چjB0#'0�0�!��9�IV�	4���4��6e(\�b)��(@�q�a�ē�hO��v�����*J~�ׁW�Cw�1A�"O�����$T!�aa�+��@�"O�)8��$��X� l��S�"O�,)@Ӑ8��y���:j���S�"Oz�31��uB�e@� ȒPH�"O��ѳ�0ai��q�NN/~S�p�"O~5�P#��h: $u�V;����"O��{�EL���D���;)f��r"O�Iڡ����%E������'P
�9�m�j(:ˁ�ޡ^@���$�O ��O�D�O�A'��T�R% ����>�����ş�Q�	ɟ<��ӟ@�Iҟ���ԟP�I�L��[	�✋�iS�i~X� 5�i!��'�b�'"�'B2�'�b�'�X C0+�%p⎜��o b��a!h�p���O����O����OV�d�O��$�ODeJ�h_3,D����ݲF�x��&�Ц��I����IПH�I㟖�U��Ο\���f��d�2䇉W�PF� *��Tz�4�?���?)��?I���?)���?Y�DX2����u�TXI�.����iAB�'���'�R�'��'c��'�pq�R�I�TM�6��/>o�� dh���D�O��D�OF�d�O����Oj���O�Yz��Wg�Ƞe�e��-R$�����؟�������	��,��Ο����䫃$_H��x��՝�f1�*Ҧ�M���?Y���?���?9��?!��?�)�7'vX�@�]�V�*P��ǭ^��V�'��'�b�'x2�'���'���CMv:�A1GZl$���SG�7��O����O����O����O���O���L��L@񱋖i�:�A�Ć&{��lZ˟���柈�I�@����I֟���(� ���_l8$�@ ���~�-
�4��$�O�˓ш�,�!��Q�<�@�!��8>2<H�>1.O\��<�<�MC�'D\q��H�*Q� ͱ�i(��M����?��'��	w�OD�l�b?���Z%BT�p&ȒH�����d�`S�A���4<O���g�T�0������oNRi���'�IO���O��� �tP�遾�@��a)�nXZ��TA}��'�28Oʧ	MB���i�::u��W�,� 1�'��X���J�O�I[��?A��q��HF���	�0���%{��o�jyr_����j��~�d��RO�u���*G��>V���I���<�"�i6�O"��F)!���B$^5`�	�=r��d�O��D�O�%e'h�b���T������1�
I��,�$bb���M�Ȣ=)���6�S(9c����ݍr ��a~ʓcy�I~yR�'��vi�bAg%�)��Jc��k��Jd}��'�6O&#}��u�F��(�y�A�¹`"�iR� [~"�'�F��	6��'��ɰ=��A��\9=� �+#-IFbф�ɵ���f������wQ��)��2�u+���O�m�|��\J���poZ��?�$�*P��]E-ߏc"�  1��"|Z��n��<9� 2]�:��.Ot�ik�Y����%i�&����ސb8\���O��d�OX���O���O�"| *� pnP!ɴ�ŋ/����N���IП<��O\���OIn�A�Ju��T�ߑ#����IW�{3��$���I����	 7�ao�E~Zw�#�C�#ry��9��Á/E����B�"=��/��<�����m�q�9��ٷg�B�O�4�'�R�'�"�?-�t��xM���0�#
Ԫ��r�<�US�����p&��O���q�Έ�haE���ji���C+/����4m��i>Iٰ�OZ�O��I@��=@xe��fY�H��@�d�5�O
����($� �F#p�T�iP��)D0x��<A׶ip�OL��'��72/ֹ�v�� =�sˋ�V�n$oZ:�Mk�'ܶ�Ms�Oڱr����s�*�d$�|���C� x�>��ßd�'��'Jb�'8��'�7p^"�d%�D����A	�FH�'�r�'���d�'�\6Ma��R����O�2\[%/�
~8q��J覹�ݴՉ'��Ov4�	�i��d,y��ŋ5A�)v���JT��9�2��X��ɯD��'
�i>����)�t,��3퓎1��z3�꟠��şT�I`y��>���?��1"��� �G���2�V=<PUЉ��<y��Ms�|핼��q
�-�2%�HL���\���D6Eʢ)ڇ�v�i>-K��'�(Pϓ<wZH*�ȑM�Ѝ�����j~Q�	��0�I럄�	t�O��ĝa�~�Yֆ�?W��!jሌ�d��)�>9.O��o�g�����F�$Jd�㉀��X�c��	�?�R�i5>7���:7"�]�'"���F���?�sB�}��C��<=P,+[�Li�'<�	ڟ�����0�I؟`��R ʱ��~u��� ���C���'�f��?i���?YN~z�%���2B���v�� �ǝdeX̓�^��ܴ���,��CѬ��$�.F�,P����Y��aǫF/K��	)(H-�r�'�V=$�$�'�щ�- ./�m:bF%����q�'��' ��'��Y�$ �O������U�eN
:�(����*q����צ��?VU�`����tϓT$��+PB�!Gn"iq�BL' �rx����-�'� h˥�I�O��.̗h��T@A�.[QM d� ����'R"�'���'�r�S
e�L!�s�]������c�%�����O��$�K}�]>�Pߴ��'-�(�rT[01Y%M� h-XN>Y��?�͸ݴ��DX�/��D.ydz��OD7Xˢ�ے%�)& Y������4�����O��!,�)�3e�4�AK$�	�0���O��G$�������ោ�O��%8g�P���A�L:T?V��.Oܔ�'>¹iO��� ˺x�/�iV�8�"X�R��ٲ�W�e�"Pc ��L��3�2 �J�I�Q\�(�"C7�
��S�����	ߟL�	��T��m�ly��Of��`�'r��� ���,@,)!W�'	B�'\l7�%�������O�$�r-]�}������q��(��+�O��ě�x6)?��J�����O��>��*$oL�TV6`RQ���I���$�<���?Y��?����?aȟ� IF
�%Q���	Īۇ ��b�>����?a�����<q�i��R���Ը4-U8�td[���+�(�nӢ�&������sdpӜ�	�%S,���gG�R'�P/dP�DR�|��C��w�O��?���a\V��A���YF�q#�X�sD`����?��?�+O��'~"�'3��=`����Kr�I1
ҵg<�O�l�'b6mY���)J<���f�j���r3�X�o'���.O� �*ɗtB����&:��
�?��F{�Hа�Q�:��s�?$z�i �%�O����O���O�}2�'d0h���j���X�Κ�~�q��/ �IJy��mӬ�P��9�t�P��T_K��ږ'�n����ɫ�M��i��7-׶L6m4?��m\{�p�	��R|��0$�+\�	��Q�h�j��K>.O����OH�$�O����O�7��M�84���ur��(�<!�V���I����Ia����Z�+��$d���ߛftR-��
�=��d�O^�d(�4�����OT�enR�[����)�x�vD�!�ҽI�6�,?�A� L� �Ic�fy��ŤZ�Lq �
�I�|��)�ker�'�"�'�b�'�������O� ��0f�0<���˃*]���D�'S^7M#�I'��D�O���T����s��p���ՏK?�Ȋ�M�V��7�%?a#�S�l�b�|��wcz8��o�bH��#�X�&\�q���?i���?����?9���2)ӇX:��e-<����'��'����?������~v�*a�R���E�;�R\��|r�'�r�'��q��i���1\BĹԭ�+Ji�):��I()2�*G�0K��d1���<�'�?1��?���³",A{�kM�6�t���ꌛ�?�����DWx}�W����e�TE�;s��P��(&*���B�I��DA}��'.R�|J?�Q�����)a�dM:H�lpD��R�dL��jmӢ��'���C�]?QK>�!㒆b�v �d�83�Ri���O��?����?	��?	I~�*O���^[�����6+Qj�Z��E�R�x���O��香�?��Z���I?x<����s i���l� h��ܟ|�# ���e�'s8DAv�\E�Ww�-�/�_p�%Z���6¦8��Cy��'Ar�'7r�'��?��/J*s*yZ��ѽ���d�S}�'���'��O���g���I+P���xR�K$� �Br#�	~�����O��O䓟��R� q�n�I6]������S�K� 9AV��%Y
�d�,q��'�'��I��8�ɜ+����o��N�z��,Z1^<���Iݟ8�I˟��'\���?���?��/��j���/?ܽ3뀲��'�t��?��	>�''*��T��a�P$��(]CH �]�,B1��W5� �5?�'�d���y"�G0K�8� j�&3V<�ɐ�K��?y���?	��?ُ��w�"�ǽ',TQ�J<X^�)j�,�O,��'S��'7�"���?]h���8%!�1����lo�y���X�46��f{Ӹ�X�e�^�5��m;������H��:�h-ea�p� �^t�O���?���?���?���F���)~	l��֩֊L�6�R,O��'���'������'�xQREZl�s�
�>xr  �m�>a��i7M�@�)��a� �Uǈ���][�	��\�Rt���X��O�Ф(���O�|�I>!.OtTۢ(�u�f�s &\�&Y@�B�Ox�d�Oz�d�O��D�<�`]�����w$`��&şI�~Y��-�޼�I��M���O�<����M;��'g�ey���rv�-;�(��X*����M��O�8
gi����D4�����2S�ڸ����N�u 5�'8R�'br�'i�'�>����ui�1�O���J%A�!�O���O0�'
�'�6m!打��-��=;�e�v����6M�S��֟����?�hD����'��	p̎-���Ҧ��
<:�[�O�$����I)m��'��i>��	�,��?L�]�SJ=���HǄ��P�d���ןp�'s�듮?���?�ʟ����&�vi��p@G6c;l��W��R*On�$i�� '��Z� ݃1H-��KD2A��E	Ч	����@"?��'E��Ā��E#d p��'j�(�hTG)@<���?����?�����'��W۟��LV��u�G�)<G̀q��O��D�O��n�Y��	���+�M��Ψ3m����1�j3%,ۛ��m�VLc�.g�4�5o,�P���~�d(��ܑ_�<��E�-V���C�'��P�	۟4�I�$��S�D�^ '82����'s5�"��>�����ҟH%?�I��M��'� R��X�}�H �B�9�����?�O>�N~Z�E�Ms�'v8�`G�r*v�3� ��t���
��*����X$�����'�4��I�~\��x��M�v><qP�'���'O�P����O���O���Y�T�<8��$����� �����\j�O�<mZ��M�x�՚Z��fL#<4�T��.3f!�'h�\�c��'|��P!���V���P�<OPXht�ۡO0����,���I��'���'X��'��>���tI�����7�zh�#�,5)�m�I���d�<�2�i��O$�i�iT��o�)j�t8;��+EU��D�OV�$�O2��Ťx�����Պ�~چb�#PIk���t���H#)L��'����	⟬���h��$@��1ycc:ϬLJ���6>��4�'t��?A���?�I~�A6h�r��
v��9@G
��_�D�z�S���	ڟ�&��������
SD�q'�� ��J��V�4,ţR&[�%�'�Ҍ�T��X?�J>�.O���h�)z�ɕ%\�JB��R�Oz���O����O&��<Y7\�H�	((@�����qJ��	8b}�	-�M��'�>��?��'h�x�D	�_4x�5��Pkb�bH�0�M��OF��V�G��(�2�l��Q�fπg}f-*�`�!K\��O����Or�D�O���,�' 龕���@�%��b�i�Z�����ȟ �I ��D�<y�i�1OM�b�ވ`#�	:��F���S�|��'z��'��kD�i��I�@5�����@X�W��)%�U����\��"�Ī<�'�?���?!A�9�iPK "�� Qf՘�?�����J}2�'$��'#���/�b	1��R�>젶g�Y��˓���ԟx�In�)����Xy�����ٛ  ��4�����(��f����S�L��d%��M5D�,�;�"]�p����۬���$�OH���O��d2�)�<ѵ��� �x�s� �tȦ��&̢B�*�XF�'t��'��6-=�I�����O(��l�+J�,`�L6�R;A'�O&��S�R#�6-%?��J�*
^c?��UB>��=KfbL#,��ĩ J�Ox��?A��?1��?�����̩2���,�yPH�@g�I�P��?���?����o�b�ɬ?e<Y$j��� S�M,����OI%��&?-�tl������h��kG`� LBt��R�W�\�I�v^V��'p �%������'�V��
��mֆM��.Ňiu��J5�'���'��R��2�O����O���R�mEZ���j�Ŋ�rn��8تO��d�O��OZ�[�C�G^�ҒC�pV:Ua�M�<aa�F�/�f�ش#�OU�����y�Kءf��$P�+/	H�yק��<���?A��?)��i~�4@1���%/�ME�`;�`��kD���>	���?d�i]�O���˅]�&�����}�!@@� ���d�O��$�OHq��y�"�Ӻ�"������W�"�|2®� 4ܺɨ%�iB�'���Пd���$��ƟH��~�)(t`g$"4K�eXD�'9 ��?���?�H~�b��d�:]�Z��m 6#�P�`Q���	ݟ%�b>=!�S�f?��� ���\j�@v�lhV�:?��̋�$��������D
`��� p��!@MF��3h9h�n�D�O����Ot��O�˓R��	ǟ���]�H��i&n�!Rh�X�Y��� �4��'�^��?���y�k��;S�����ܘ<󜈹k�7c+� I�4���Z�jߎ�
�O1�OM�nD�9�@�
O���y�Re����?����?���?�������"�ō)�Ҝ٤�O��L-{��'�R�'�fꓧ�D�ئ�<	B^�U������7-�ЂA�IE�����şS�ϙ��q�u�D���n��A,� �B�Z�ܽM��P��O��O��?���?��r�*;��$MB�bvB`22!r��?.O���'b2�'�R�?�[�"/0�5�A��S�i���<AbP�P�	֟�$��O)�YX�i՟L���Y"�
Y�z�ЕK&��شr��I�?y:1�OT�O2���@�wz�րZ|�É�?����?���?9M~�,O���&!#���'��#�ʨ�%�@v��<�i��Oب�'���X�9�!@�60*dB`f�-R�2�'u�`�R�i��	g(|D�����" n�A"�@>�I��D���rR����۟�������ǟ��O�L�x@�q]��XT$_�S��B]����㟸�	_�s���ش�yү)Z��!5���T��LY��?����䓵�O?r���4�~bg�BVnM*׎М3���b���?9d%ڤc���w�qy�O2ə�6�:YA��O��ä��x<��'���'h�I�����O����O�a��X�b"�!��� �U+A�(������Ȧ�PܴCf�'����I�m���7 b���r�S����zߖ�S��.?ͧ6���$֝�y�f,*۔��&�Ǿ@ք�;�o9�?���?���?Y���c��Ӗ�D�&�����K1��S
�OL�'\��'��7�!�	�?=x� Kd��c�j)p�R����HП`���
�4n�h(ش���U�\�^a����u�.]�fN�\ö�Q�I�x�����+����d�O���O��d�O�ۀ(�l��SB;\�P	�gA�	�Tʓu��I柸��Ο'?��	�m��� @J�d�P��杼E)��O�$o��Mӧ�x����ڈqsnU9��ڑ|P̫�����]� ���D�']3���*�t�O�˓]0{2�ȘX���H��ߜa�Pu��?���?����?!(O\��'� Ħ.KiC4NW�C���w�U�O��q����O����O���	8;��]fo�U���Xt�X�;���7�t���c٦��&.�>5�;7R*IQD͂t�Q;������ԟ,�I�`�	��L��P�O8�q�S �.�6�z�ǔ(¤2���?��g��Ii�$oӌc�\�V#�FI�":E�8l���NE�	��M㤽i~�$�(e�����p��r|�� -�p�h2��T�`�&�1��'�b�$�ȕ���'���'UJ|���ŁR����A�8諐�'"\����O&��O�0u�Q�b�R��e	�=쌘����iy��>1���?IL>���a��)Q�)S`$��`Ӝ�R�鞽	������d�:��$3�D�%F����3��B�4"��95�����O8���OF�6��<Ʉ�'��e�!�S�%Ɋ�7�L�Ja��j��?I�����D}��'��1�t�!}�>�K`�En�I���'��D�	ϛV4O����1T��y�O?��?qiF\{qA���.���Z�l�6�Iuy��'�R�'���'"2�?�*�K�+_ώ�a�(�,\����y}B�'��'�� m��<a�퓞s@�+4��=%���h�����	y��_�5��l�R?iC'�b^�u��M��t%�����ܟ�*۔	���=�D�<�'�?	�\�P/�ę�D�}p��ǩ�?����?����VX}��'���'��81KտN�D�d��G�������v}2guӈ�n��ēY[n@����X2���+�x�L�����?!'C�8|��Ѕ��N~�O�����W�G)h��Yx�d˨0�Ʃ����1���'`B�'��S�<� p, ��x��Đ�,R)@1�q��'!���?���T9���|�'���bU17�te�5@�{�.�P$ώ={S`w�R�l��MFD��M��'�"��.E����07
4�;��]5R���*'������ĕ|[�t�I؟��	矀�	ܟ(#)]��n0H�$E�`W�1[�I���Ľ<i���'�?q�L�&fX��w���Q&�� ���4�M��i�`O���8��h�m�S�.L�[smڎEj��4,�&>|D˓k;FA�c�O��IM>Y-OP��E�V���Q��n?b���+�O����O|�$�O��<�$[��ɦ(�x ���$r�x-�$c�GZ������M�L>��	 ��:�Mc�i�����Md��3�ï ��y!�+�:4���i��D�Op���c��:'�<��'�yWg,]�����@�
fP��C�?����?���?����?���)��s$Ms�@��dNz�h���	 r�'2f�>!���?!�ig1O4����� ���bC&�����|�'F��'+ ���i��i�qqPf�s���h�eyu��V��������D�Ov���OH��E�c��p�q䁅_w�p)�	Ä!����O�ʓ]�IΟ��ٟ|�O`8[�!Ŋ;'x��3�D�}V��X+Or��'{��'hɧ��FZ��hFa�6V��K�(�T_�����3~3�7�FBy��OZ�����,�Ջ�Y�G�&�A5��\H�!���?I��?��������� ��C�8p=<d�����Z��1s ��O��cě���s}�'`�0��E�-#a�����.3�\�BŨΦa�ݴY��9s�4���-na�����1�H�'_�|����_DU8ԩ&٤2:Y��zyB�'���'�"�'2��?�*�i�Nd���L�&����]}R�'a��'���y�eu���ɪ[��XV WZ�3��)^ꀩnZ��M�x�O`���O˨���is�$ʳC~�Qd��'A����A�%��d����H��-ғO���?q��7+H���0i�L��vj�&B<����?1���?�.O`��'�"�'�iB�x�&��6l1��T����:Hc�O�U�'�i�ON����!+����T�`��4J��'o��>I���zU
�!���������F�X牐%�*��g�F��*T��22\�d�O"���O4��1�'�y�f�h�^@*7*_�.���!�?�'Z���'O�6-?�I�?�3����u��8 R�Z&k��eM�ݟ��I��	/k��l��<q��H�~-��~��N!Ue����&��:�pg�P[�Iyy��'���'�B�'u2��|x�MzC�ė$�<�a`��I�����<�����?��a� �0H�Q���̃�_lqdQ�X��4/țv�+���A�As���q��?
��M֬,i
غs��>�ɭY��t��'1|�'�p�'�8��O��F�<�S�LA6�Yq�'��' 2�'�^��p�O����6]#��І�̛oф��%��MZ��DRɦ��?��R��ݴb���O*M����v8�K����	�iS�N��V���;�E�K����ij�Z�%�10�����˜)�W��O����O��$�O ���O~"|B�G�3>�"��B]���)�7�M͟0�	̟<��Ol���O�Alb̓lze��R2s���iC�u��hH>q۴u�&�O����i���OX<�����\�x��A��ƀ��^ �.���B��O&��|���?�[���b���<񌕢��a�������?	+O��'�	֟�O%"	2kМA4l�9�
�,��)(O���'�R�'�ɧ��1p���%MQ!iuxl����1K��EA�"~ˤ�ƞ���ӄE�"�]O�M4,D�qN��O���̂>[r%������ƟT��v�My"��O�2&� RЩ��a��j!��'F��6�M�Ra�>Y�A\�+'�O �c�%�	|�����?�V#���M��O�B���|��W0/I�}�#�˩{�LP��й�?�*O��d�O��D�O����O��W5pPG�[l��K���T�&��O��d�O�$#�9O��nZ�<u��0c����Ճ �A��������	l��i�S�g��n�U?qs��hjthP!��[zZ�I�g��T�F@W��-��<i���?���~C��a*�@X�³���?y���?������PC}b�'V2�'���ز擁՜�ɇҢ1� ���v}��'U��|�F�i~Z���"��AK��Ѝ9�IOR�t�&�]٦��H~�T��l̓pY�Iyre�(*��ѥ�E�����ҟ��I؟t�IK�O5����<]@���(i���I5 AB�>i��?1ıi��O��iP�9�v02�MA�Xh���$d�d�O����OҙSt�m�|�Ӻ��CQ���4��/C� :�)�� ?�I	�@�(��':����\��៸��ş��ɖ3��<{d�C*&� �F6O�E�'b���?���?AJ~��� ���3 无%�.�Pd��a#BI��Z������ '�b>�HQ��5��X�p��&Iˈ=�ч�+|-�tl3���	�H�{�'W�'���X����%U&�e��-&\f������ޟ���ܟ��'S���?�X�T'��� ,�8��`�E*�?qòi�O@��'0�'e�Q(WY�e�ގPW�4�0 �9*��+��i%�	�xx�$c4ڟ������|
T�b��$L��B�G� x�d�O����O����O�D'�g�? 0d8�-� �a�S��+V�"h���'���'�T���ę����<Y�(�g�*	�F�5_��̹�A�ݟ��IΟ,�$[禍ϓ�?a�F]�1��K�+�T���Ǝx�����꾟\%�������'���'N\�s��)V� q)�b��-Њ��"�'�\��[�O���?�Οr�Pdլ<��]�uAV!_`p�cY�� �O~���O��O�65�����}wF�ha'	�e&$1j3�@GA��m�N~��OE����!W�x�U�U!@d�2E�6\�-j��?��?�����'��HƟ��Qd;��%�" L��H ��O$ʓc7���$O}R�'��X�D�%'Xبu���t���'r� ��af�V���qd	�0����@�l�%%Y�A��AN�J����'���ǟX�Iş��Iß��I���/V�	��>r�-��fܘ3f�	`y��'G�p�m��<�p�]�g�)�Oȇp匙c-�蟤��[��H��H��nz?�R朁Le�H�Pe�~^�YC���۟�4��=
S��:�$�<��km	$H�\8�$�{�UAc�]��?����?����ğa}[���I�q��8��N2A��i���T>ڬ�?�qP��IڟD&���G_3OLigAVQdh�2�\jy�	Y����U�i}�i>a��OP��#*���8��yc�jte ����O��O@��4ڧ�y��^�����O�a%Lt�6���?�4\� �I���Rݴ��'}�T	���8X�Ug���Qѭ�%|��'5�'ӘaR&�i��	�m^THcUY?��5� $�X�Af�2��Uztk:���<����?���?i��?�m�	58u*Q�	Ox�g(����r}2�'���'$��y���j�	k�];.�XYu�^<��듦?����S�'��y
���eJ�$<L�vp���M+�O6���4�~b�|�Y�\�@����,-�`${^�+��_���I˟<�I��x��wyb
�>���n��\sY	�u��.3�����۸�?Iw�i��ON��'�'�󤀁RT� �h�9u�tQP���
-Ď��4�iY�	�M��# ��)U+ue0��N�#��������I̟`��џ\�	� E�Ԏ�&�vQ{�eF�%?`<�Q��?A��?9W�$��ҟ���4��'ߌ!�h�+(�=ȁ�S�M�O>���?A�,d����4�y�֟P��}�5�#d� -�liA��)kTp#��O�O���?!���?1�@��IZT���Y��bo	�/������?Y+O��'���'\�?]�M̉#�n�k����NS�0QF�<ɗ^����ҟ�%��O���e ĕ^�l���ߝ5?aP��/Fѩ�4��I�?�p�O��On�Q��M�vW�E�t�>�0L���OD�$�O\���Oԓ��˓a=bk�#4��"p�f�v5J'���?a���?Yмi��O��'���K
-�vY�U�	�n�Z�ZX~�<*���?�v��4�M��O�.N��Sy�#�c@����G�G>^=c�X��?.O�d�Od���O���O��WW|5)F*��v��p�cḴTb�
�OR���O��D1���O�nZ�<	�aۦxj�qqO  �@@�g���ɓ�����`���4�~Bĵ_t�q�p�I�g��w��?�E�Ŗ��ې�䓆�4�B��T�"Ā�4mo���K�>\�����OB���O�˓��՟�Iޟ� aǒu~h��˒09�0@ a�W�a���,����5P�9�0��	?�P��Z3lS�5I*O�4xD`�&�fM�G���S
L1���<�H9?z���5��-/Z h�3�Q����	��������F��:OZD)jԄD�9�	ˬ&fh)�'����?9��y&��������	0&�=��\-ή�i�I�O���O��n�2;���o�u~�gC�(�˺k�&C�@�#2m�q\ZLAAy��ayR�'���'���'�; ��أ�A�JP8q��eR�e��ɤ����O����O`����) T����%J��|���^�ֽ�'f*7���K<�|��[@k`P)&f lЍZrX�dd����F�����!-E����͈�O�˓b��2�@s<<Dj�T�@�@!��?���?����?�-O��'�b��%
Z��ec�)M�u���{�J㟔��O"���O��	-6R�K���4"�pk�M��h��g���YV�5�R%+�'�y�e��g$�m�k��<�N�1U���?q���?���?���?���K���`*њfN9%l��ET�'��$�>�*O�n�S̓h�~��%Lѯ<����΃'��]$�����P�����l�|~Zw�~�s�O�o.�da�ɉ�U�(�@&����*���<���?����?��N�T�N-	�l�)�@�Ҡ(�9�?�����dq}�'�R�'�ӊ1���NI�v����ӮX�B����0�	q�)�t�R�a�65�գ�/2�9Z��R�����π�M�gU���*T}��+��U?<,pzE�S�<��YH�Z�	�O����O�D�O@���ʓ+M�uV�J@$J��C(��?y/O��o�]��N���՟����N��`Q�cܦmk\�A�ϟ\�IR��o��<��Oi�\Y�ӟ��-��M)��/X˦ٳ��ݛ[My:�����O����O��$�O���>� ��r��F�D@�)&�C+��ʣ>!���?����䧚?���i��D�8t؉v�ѝ<'�`5����y��'$�'���'l��.Z�?O>��s�V�l���1%��� ��OZ��M�~��|�S�d��͟�k�AW1/1TpiJT�_��Mhv,��P��ğ��	Wy��>�/O���[�9�Wd�ה��@̺�㟸�O^=nھ�MC��x��=Ϩ�8��Ǜ��}�q����䛏z7F̫�V?���r�������.�a�wL١v��ZeL�AS\���O���O��=ڧ�y���i��	��A��T����?��_��' 7M?�I�?� ��,	ф�j��8M?y�p���L����I�CD�Lo�g~RNӛ@�2��κ��AR��K5�̵A�W۞y��'��������x�����	d�d)�5P8i��={AJ,M���'�8��?����?1O~��B}P�QEC_��=���΃V���eW�|��ǟ�&�b>�:÷T�*���j�=����,�8i�DlC~rǹ�-�����$^�&�\�S�ʆ=7�����#�D�O
���Ox���O�ʓ#���� �Ƽe�(1Xa�.=�H�i�ן� �4��'����?����yr!U
.t�*��Dc�`�J͌�HOV��ڴ��4$��XP���o�A��� J�@�ↈ���Rt��OL��O���O���O�#|�`�I1�z��Y�8�J���e�H�	����O,�%�F��(~*�"F�v�84�C/K)Y��'�B�'���I� Y�F����!C���H�(|�u͊�p��ak��'D�%�p����'U2�'w�0)w�! *t8� �2�[2�'8�V���Ot���O�D!���[�
���0�EЁ0����Fpy��>Q��?	H>��VYW���
P�RA��*�!�QiU�u.�P3�������|��
�(�OK^�T�FIH%.uA��uk�&Q�'��'����P��p��?.i���C"j>\�4�1!b`�	fyRrӔ�l۬O���EB}R�j�,Mϲ5�Hͨd?j���O��Gt�0�S����'�����EE�05����B&Rz� *!�'P�ʟ��	ݟ|��ğ��	W�$[-����w"��
��*v���	���I�$?���M�'���c��3�`P
Z�*ㄘ#���?YI>!H~j��ڄ�M��'�I�S��"ZI:���	�́��<h)��OXA�I>-O�)�O��p
�.��(Z�Y+%F��9&/�O����O���<�S�8��՟��ɞ��j�X��1 �&�V��?��S��b۴/��V�'��P�/���!��Ҧ-�Â@ɓ\�J�I��i�4i�Ox�xI~��Or� �'����iъ#���c#��8�����?1���?	���h�*�I�4L�aa��>Q��)�%A4h����H}bU�T0ܴ��'��� õ3� ��K"uQ���͕��2i���l��M��с�M��O�0 �)X���v"O�S���SA0Y|xȔl�x?P�Ozʓ�?y��?����?I��
q�m;ҊH�n� ��b̒;j��hZ/O�m�'���'Kr���'��|8FbY [gXthÆ�/��5J��>9вi7-U|�)�S�B#�e��"��!�ɰ�D�~���8�(��>)�Q�'x���փ㟰@��|�S�x0�
�4zh����#�8_��iA��@�	ʟ��	ȟ��Icy2	�>���Eᾖs;0�ia�Y*�ᕨ�`jߴ��'V���?A���y�1�h��B�# �(�� �3X|�rڴ����Kθ�r��ޅ��Ǜ4����FZF��� �O|���O����O�x����%�'m�i��t���"d�)��d��ٟ�����d�<�5�i.1O� 9韧|��#��32�tu٥�,�D���]�ݴ�z�.V��Ms�'��㌶C��X�f�1(�䁒F�w5�}�bJ����|�R�@����	ş�U-�(&Ax����ä��aH�]�p��{y�>���?����IȘ6vT���@�-z.��կ��:Q�	�����O"��/��~:gf]A��m7gED�"��ڵsH�a�"O����'��TmK|?�K>�Ə�D�`�%� 8~�6h�
�?����?Y��?�N~�)O���ɝ~J��M
=7���a:I�h�d�O���Aڦ}�?&V����2)�"B��-�>�s)G u����I㟨y�]Ϧ��'�����ed�;��%2���z�X4�h��a	��	cy��'���'���'�2�?qa�ϰD�z�kU�WC���2cO�D}��'�2�'���yB�wӶ牽|�S��@��v����˦ 6����O�O���6����x�^�I���i�c�utp��H�?��P�!9B�'N�'$��ӟ��ɶټ�b��;p����2���Gx�5�����	��'�D��?���?��3Sd!����,P\-���=��'����?����3]�9PFʹ|KT�+���;��В-O�-!�n{�p7��n�Ǧ��Eh�
]T�yb�b�L:B!�yW>]8
�GNm��M��=(�@86fՈU��Lєa�v��z�#�U�=���	se����)��c�dl�@/^�.�9@����)�WL�R�pB4hT��y�*��w)�ĈEk
�s���Mޙ%�D���]��(�&���Ub�Q��O�?	-�]qT̋�w6����D�
��3��Iє�٧�r���I�K�.�)"臹Q�f$����iJ(�0�n7H��T�@/&0q;�%ƞ���֚E�6��񄑲{hh8l�=h����m�? ��sԨ��|�x!�2��0�0�⡦�1Y�"hk�=?)�c��+v�M3E�H�O����!�Y ���33�$r�qa�**i}��$���Z�V��'8RA�s/��2|�rw��Ӛ��e$̷8!뉄�q������]����2�I�@� �z�`���i�킛$���i׋��]�0 �%�P��1F@�M5��a���W0x6��w9�B��h��ؤ��,v/FQ��b�&za�q!f�ܗzt����Z�F[f�s��Q]���87�߮x� AD$F����'�����$�OГO���O�}�f�Z�^P�a�F�����c]�<	�ښd��D�Ov���O\����ӑh����� h��4�C7X��<�����?���;g�I�'�4*0* �f�h��I�)�ٚ&b��<���?y����'=��Sʟ�q�9VD 0��O�=����Ӡ�̟���k�̟����|�� �	m~��؁�����@I*1;���?����?�cK��<����I�OD�D�O��5�^� ��u04#z`��!�?��O��DG�B���d;�ԟ~ӑCC�Vڀ�� �3�Ј`��'����':Bam���d�O��D�O���'���Z@�ʫ,�>ɠ5bR��q�'���'�����|±�	�bu����,�,�1�ʫgF��{���?���?Y��?i������O���&�h�[��?3%4Eb�E,~��2Cx��y2�lϓ�?����7�1E�5�$��c�x��	ɟ���۟���`y2�'k��'����h+��
����	-�J�I��O*�+bK�O��B�7O:���Oh�D�wQh� W;/�e��N�&���d�Op���v}�W����G�Qj�Q�m�.쉡Dןx ��'��:�'����'s�'v�?�r��!U�(�S �W�%Kب�C&�O,�'��	ҟ�$���IҟȘ��[�;L�a�w@��.k4�yƎ��V.Z����Z�ԟ��ɟd&?ys��d�"%:gd�-f�lk�A�+c&�	cy��'G�'N��'����'���3m�E�Ju��	@%JH���Ӟ�y��'���'r�Ow�'�?�֮��	 �!�G�.ʔq�A���?�����?���O�ʀ�y���}�FHD?^8Z��π��?���?rLJ�<I�	���џ|�I�h��aNkOB��b�2qt5y�Jz�I�0�Ɇ=���?Y�O��a�������a���Q�9��͓�?9&�i�2�'
��'/ʓ%9P�X�G��L(caD���Iy��'���\>�e��	��4"��-i��̪V��1aN���㟸�޴�?i��?y�C҉���$S9Z��-)�!
9f[Ъ�L��?����?	����|�A
��<��s�x+�(#!8�M�F���q1|ð�io2�'�2�'�O���<��-��
�>���I/X����d��<�IL�	��tS,?+�Dp	A%��U6L�A(�$�("���O����OP˓���$�	8u��s���:`,�=�D��B.x&����<x����?��|��'%��QSdIg�X[�@pÖy�����$�O���2�	��TΓg�N�[���X����!���F���	z�`@z��#?Q��?ͧ��|>�16�K
��ת0D�c��=��I~��?�/Or0��ņ�H���$jU$%�u�6h�|�f��'�'�Y�$�Or(�y�ˍ@����=XP��6-�<	���o����t<
}S�ą�~�z����\??��'�B�$�y��'�맖?����y��%}�r�[�!�O��������O@��.�9O[v*J"\Q���3.H#+���R5��O\�9�
�<y��?����?	���ĕ��
 �!�]�#n��b���ji���O�˓qTXFx�Ou��KA�R(zD�@�5'	f�*�fKZ�	̟D�	�T�	��Ĕ���ȉN�n!� �ħ#�աS�<�m`p�Gx�O��y�'�.�&T�ș	���cf��87�GJ�t6m�OP���Of�DDN�)
�'�R��F��@_D��BjZ#1�)z��?L>	�k�̓�?��?����+P\�`���h�G�?���?��xʟ�O��;�"ќn0,la �ؾ"�$C֧%�$�O�ٸ!��0��韼��<Qr�L�y!z��C�R�kجm �oן�'�R�'�O(��c�PX���#g7H]ڣF�t�5y3N�O&ŉ�lB���OH���OJ���]�+���b�6z�\r�Ĝ��d��?I������4�<�N�>�d[���dF���(�p�|��<O^��OB�8�i�y��'a~Q Y�cO��8�!�1��D{�'p|\��S̟��O�ؘ$L�`�V�xwLV!e�����?���8����?�\?A�	�x�;2��ы��J1?Fԝ �4b�ֵ$���'.��'���yBO�	)���aҏ2ך%YD��?DQrU��y��'I>7-�O����O�$g}r�J[�΄��N�48��ڗO��\H��'���>��d�<�-�n�r�DQ�8�Є3�/pV]�!�_R1P�$�O,�n����Iʟ���;���<�2)� 	���{v*Z�K4�؊f�:�?��
O�<�����$�|B��S�|�#�v(K�/^�°����6� ��ǽiQr�'���'
�����O2�P�� `�(�'�Ui��M3A��˓��d��2���ѿ	p�	�O����O�P�2��,�0��K�~9@{�-�O����OJ��'q�I�ؖ�~�ɯظJh�O���P啄��
}c�d�*(�����O����|Γ�� ��1���.}��4@��@6.j��s�'�����$�O���?Y��?���-ȸ�)��w���r*B�׆��>.�s���?����?�'���?)S�.S�Pl�s�L�>5�4�6,�O"˓�?!+O �$�O��d�y����#`�Eㄩ��52�p%@SM�T�	�'���'S"����~R��0-���� 	��h�IVg�*��Ĉ��?�(O���O���NL��*?q]����$�&mW��S�;E"�'z���y��'*�'�?!��?��FC�%�tqh6N�G1ڭ��A*���O��OHm#u��8�'�	H"r���@ C�J��)Yx,��'	H8��'���jӸ�$�Ob���OT�'	�x��Z .Y���&*ѵp	 x��'���'�訜'�2[���O6r�[+Z"];L��t�ӿC�4��\�"�'|<7m�O���O���Pg}P����:'E���%�D0�4�%�ܟ�Y�k��$���O�>݉�'J�o�f7��@-	+~��@,�u��6��O���OH�$�P}B]����<�!��=?0�)�K�w�e�0�����IXy�*(�y� P�����'���'����B*[�V��͢q�P��>���'���'������Ox˓�ywZYbB	H��F��ٱ@%���"��$�*��d�O
�$�O.�'f7�Jċƅp��\:�肦2cX-�����<Q�����O6�d�O>��a,W�S�j�iqm%�&�!�e����d�%i(�$�O���Oz�'�?�S�Orx�b�R�~4j�a��
�Gi�Y/O����O<�O����OA���O�	x1a.a��ZV@�M�`M�7�C?�y��')��'��O�b�'�?��e�(P%~X���T�|���y���?	����?��� X�����H�{��許`F1%�tI���x��';�m�(�y��'~��'�?I���?1D_$'�A���'�ⅸ g"�䓍?��(���Gx�O |	զ��1C�<����z�m��.��̓�?���i���'b�'K�ʓ)7��9�Kҟ%xR��3�ǔC�P�Iޟ���A�H��e�IX���2y^,-��w��/���Ip�:]B�'�7��O��$�O��du�	ן�jl���6���7E6�h�+�����t'���O �$3�'��ʂ�p`���$����R�^��*6��O��D�O
��E��?�'@���Q�>$��J��<%b������0'��͓>4����?������V 3�dP��g� ���+酦�?��?AV�xr�'��|b��,C(�B3�T:i R���"�>W��I�`����	5��Iџ���ǟ��OU�p;�;R��h� �[q�y8��ʉ'+b�'��ǟ�����Ђ J�}rh�p�솞/� �O�/5��ɴ5���ɟ���ٟ�$?Y)��*�J�F�"=�D�Z"*?T[�Y���Iџ�$���	�<ɵ��������@Tz6#Ɗq�����Zs����T��͟<&?����O	,i)�m��@,�i�#�Ux����O�O����O�<�7Ov��,<"�eόW��<S� &�^Y�I����i�g9O����A��'��'��(�[.}t(x����d��|�'�r*�&�yb�|<��,�Uyh÷�H�Ddj6�'��`�'-b d�B�D�O&���O���'E�Y2� ��(ui�"�����?1��X\F�̓���򩃮iN�*�)Y�h��e�%ςX[� �O����֦5�	��$���pˊ}��@�MWށ�p�*%�l�7㒂&�b�A���|bU>�H��`����~Mz�%ȗ8����%�v��Q�4�?���?���M	���4������J,���Ů,�B�%�O����d�On�
P;O4�$�Oh�$ي؞�S�.�1��Р��'~�����O���WH�i>aFxR�ƪY'f�sG��]��4���Y����?�%��<���?�����O^V��֠ۑK��3d�F�� ����?Q����O��On�$r�|�d�\X�$j�l�6B�k�OX\2r�I����O��$�OҒ�6q���>�h0 �:v��=1 �F�F���D�O����O(�$)�I�xn�m͓�q��!�@�D��U��Q8��w�c���ğ��I�?u�O/��`�n�qJ%���܇@U���%��ԟt�Iv�ԟp�'���ZI�XiĎ��XG��[_����4��O`���OL8���Ol�ġ|��?���%:�bZ>E�	��h��dA$�I>�����5�����4
�HzPlX��17&F;�?QwT�<!��`�v�'�2�'d�o�>Y�ȋT�
�"wFļo����"R%��U\�����O�-�/h�:���us�\4�1`Fj�=�?���?����?����?���?i.�(A��-�SQN���A�n���'�HĪ��4��[tV�,��/��;�r�I�&���lh�E�1�ڙX��T�
Ѓ��YH����o_�9�~�	YO�r���O����*k�(�Kp�	? J��ֆZ*Ry�6M�Ǧ ���?����H~����yw�ϝ( ��w!
�}�4	�c�|��V�
�����:l�T{q B9Oe�ܨ�!5s�ycwBM�	;XDSˆTR�� �IG�lU�1�աx���fB�n�tj�k�MJ���`:l-AOJ�@xQ�ޫ
P�	��@�^y��;᠇3R�>���nS1w������&%a��
N��s�n�#1$�r"$��S�L�v̬��GjT?_�0�gÀ�y�E�!g�%��B�?q$��:�Y�1���['o�H����mW��[0#{3��RvA�1e�iz6��(�T����9�E�`H(xH؂�.@4ք(# fX,��ʢ�t�����O����<qߴ�\K��~t�d�&�=��
bN�.0@���QKiR���e�3�)� �a)�JS�}�bE���L=��5�S2����1�$p���E"m����',UbA�K�H��᩠�.��1G�4?�cAğ��Ie����G')	�у�F�v|lQQ`�y�<�D���8T��I�	�`IL5Quf�v?Y��)�*O�a2���n�֑�H�.rq (�m�t�o��������'���'���F�:�2# ��d�P�:�F�^���bR6#m� �w؞�%� ,������S"��[0+�Ψ	�K��/���3ۓ6�xl� ?�`q���8=x�T��-:	`��hO#=�c���8��$�#�@�L<$�S`��d�<���_+o���)�I�*/�|�g*d��Le}�[��J�ϙ��d�O�7mĽ^�M{���b�ء�9sF��'+��'�r��'V����QD�#R� PI���O�B\��icO�%�&!R��[,Ǒ����j�L����ݺ!��=�'`��<
��Q���@��=.$YE~��Q0�?����'uYl�!¦ -{���N^S��O���Y$V:5q�M	�^T�\@`ǂ+=�~B���K �Ҵ<�Tpjq�H�z�<��W����T$Sb�m������Y�Sßl��{7RAV Q,~o���B�Gf�@���iW�M�������|rI�	���h���2V�
̓��
���0W���WjS�o;����S�s�X��uf�5#JiPv��6T#��2����I�����~�����Q��&*�N=jE������ğ���	&o)�|p��8Oei�eH�h�Z�I� :b���ٴ�?��$�ڣh�ࠣ���6�:]Rq�0J��D�O,�B��mZ����	ɟ �'՛��J�_/��H�� ���ï��x*t���S�����S����L?Q ��� �"���#$;����5��P���\�uo�$�Sb��3[�t:P����4n(�'-z�9܎R�J�ȡ��	H+Ԣߦ��I�8��	�MS�'�?i���?���M2��6��	;S��y��c�S�<1t�+<���eCD%B>�|;u�P?���i�J6�'��[��[�P�q�0jކũ@�(-(u��B��4�?���?1)O����O��Ӝ0MJ7�@"!����$,�nd��,>a�㌚�?ѡ(� .q�)S�j�}:�Ȃ��=�O�K�i�	���1[��JS��5x���H/9$�<�5��=Q5�h�E�'�ȩ�Pa7D�`��i a�4aR�&�ְ�Q"(}�K!�ɬ0@�Zش�?����M��JM�Bc|�[� A�K���	�����	П�ja)����<�;|�E���_%"����gG�"��dD~��_��H�8����.I �\`C���r���6�	m�~�d!��`�A8�+އ4�H�!�K�>q�C�	
�z�J�Q����I-R����d�N?i%8hD$���eɰC�.�hbLGx�$[�*�Y�'t2��d�'A�fj�&�
��r-FU>	:�D�=o����R��� �A�3^X�����ʧ��'k��D�g��'2�X�`ݎZ���'��A8���2�6��"�/j)Q?�0Cɿ&�L���Z�~WH��#�>�W*ߟ<�IR~J~«O���UO�8��J�n�){�DL��y��ܺyvYA�D�
m���yq����O2PD�����(���b���b�6���'��5�����OV��7y��o�ߟ��Iߟ��'t��)ȬI��AY��<hȪY��'S2��Z�Hņ�	�|vx1�3�1*�qZ�� �nТO�����'�� ǅ�N!�8 e
M� �.�K<I �۟t��I������<8�0d����B�n4�-�F�N���؉i�����HO>eB��qnYI`�U�b� J�
K8e�^$ߴ�?!���?�/O����OJ�S�jCZ7���1���'t���� �_�B�a"��M�C�P,��p80G5M3x�łA؟l`f�.4J$gY�M�>ܨ���J���0q�fH<�Ai_1`�LC���F3@T@a^s�<I@(5 �kuJ�\���;ԅ�z��k�D�0�k�i��'��&T^���ˆ���5?�"4��s2`��?y��?% �?I�yZw*ް�F�U4X���,�9�1���M�p̑>��W�E3T�2(9I�fC���!7�B,����ԟd�Iğ�;t��x�ʀ?~���Ə�3�����?�����E�u�Ju�1dF+�&Uq�/�&G��~R&��D�d�Jo(h:0źz"-�BW��D^�7��lZ���Ix��ßDn�gT0ͻ!��d �lr��̀^`py�����E'J6P�ɧ��9�	^7S�yrnS�6q�0ͺN��ɄG�vű�lZ�)�g�? �����,����C��S�=��]�l��h�O��d�O���"ҧ0*�\��לs+�x��T6��i�OL��$lOFu:ƪNHv�E�"� HՄ���������1hR�ߊ!�8�e��Y�"��vɛß$�Iߟ(�QlJ��M���?�����wL�����YA�#H qu�!L<) �ʌz�nt��	��xƎ����pf K���'� Bѧ�Ԥ���	4^XMa�"Ǉw�Xi�4��8��p`���?Y窕��?��S�Y���ݦ����p�����F����?D�8��ؤwl�\�&E�%��b��@���4���$�<lX� �xt��!ל&��1J��^�x��"�i���'�^���	ٟ�'$�4�l����kX�r^j<i�)�
2l���N6P��n�����QA]��������6ϰ?�	�զy�p�̭S��kAB��p yy!��7��x�,��6��A��gS�0qc��A5�yb���}�4|���
�$���L٫��I��p>)d�D[$�Xッ�hN�)`7�F�<q�D�!��D�ck��r�RE�ȑ8��c�MO.Z��Q2�ł�@���-C4gc�U� !�x�(Q��X
�!�¿\����G�
��Ȕ�,x�!�Ę�D�vP�,��,��4iV`��$�!�D	
,�����l�4m$`!�$H[K�ԙ�n�t����m*�!��5�V��k�KR�A4���!��
wT$R�Cʹ<����C�r�!���[�hqy1���  �p���<%�!��0k�����B-{4t�2ddܼu�!�D363��UAW�����Ƥ.q!�d��1-~�XA�_�O	tPC7A kO!�D��i&�xd�ק8���@��#H�!�E<�"`�D *_Zi�с�E�!�������H�kN��!6雕S�!���4!�	�.�pG~T�"���!�D <j#��]88�U���F.�!�#2�*2W���3�K��-�!�DG�\������9�wj�2�!�I���R���wx0�B��]�Y�!���I��1p�%X:(z,\T	�<QE!�$�	9[fd�`+T rVq"�ٗJ!���=��FD�1AZ��c�UO!����u�U�@�mIʽ�:2!�$�0g��P��+a&(�QKC!�D��~dl]
��I�!���*O"!��<A�\!��*baX3Ț�!��	.�ꥹ��͟V pCp���P!�%Z��r�nM7B�;va�!�$��U}C�/�9��{�F�]�!��Z�FT�p���U��%ɷΊ�1�!����t!ATgv�K-�\!�$�0M�H]J�N�2D�a�Mƾ0]!��G�z�n�B��+R$%� �-7!�$��@�|	�P�K�cs,Pd��!��� ~Y椃F;QT��&J�VW!�\7d�fq
ե�jS�Q�C�R!�_�4Gʅ�R�"SB޹臂�!�9�H�s��k?L�t�H@!�䒻?w���<����,-!���VpqɁcǜ(���g�,	!�d
��ʸ��E�`�el��;!�d&T�X!�PCZ+�j�q�&�![�!�>�� +&�S�~%�dI;N!�ę�.���-�
%�|9A�ā"!��`�r���7�.�`��Y6~ !�$�����E#^�b�=!,�c!�F�-��Y(3�À=�HKA���!�� �`�D`i��!�gX00V�2�"OUS�BE��I�,�1 �Q�p"O��1��f���V�����"O��`lʡ&���Ö�?(����B"O�]�7�,U��B���0Uʆ���"O��ہ�[E�5HюU/��c�"O�I��J׀cǨ�"�$0��3"O���Ä�h���c�L��;��b�"Od1БP&O�\��jJ"��Y�"O����ũ|k0!@�I�\��h6"O�Ai�̭m8�mR�#����"OX��CJS�n|�"DJ=<���Q"O���߃�	���K��A�1"O���3K�"��X���<.��2�"O�l�"�.(<�Q�D ��!�"O��T@˘G�j��&���Q�"OX%��+L4Q�^��Ԧ� �:1�!"O 	s"@sH�9���$*�6�	�"O��A�Q>��SD��~��d�"O�� ����O)���q��w�~���"O\��0/ѡ`�l��C�����d"O ���Hۊ:[T`k�G�MCE�3D���ꆰCEH�*�`ϝM7(��.D�Ș���.2���$F�6i���-D�<�dI�-TcRm���'=� G?D��x�.
!G>��6$�O���kv�=O� )��7��'�8�f�0vf���P�@�(�}�	�'
������Nnbu�7�L�/1�))O:���垽0���OQ>��%
���W%#fNx����$,O�-ۧ�ʾ��}0dR`��s�0)���6)xU�wA�&4J�0�L�~���X�"�E���E � rf 7r��!�4˅�X�n�l%k�����S�$��Z\tQ@�-_��1�E���1�l�CKs8�(�X�pi��'����"�s���@�bք'�� Z�^q��E,I��q� ^�a�R�B��=�V܊�d�E��."P���l�G�f�:+3!�d#X�4�E��C�@��!MR+�l�©̡_H��p�ME�<�Za`�(��<څ$���O��rgBP�I8�ԫ`훸%��/OVX��&_m��9qH���'��!�V�yKZ�z��a�`MzHbi��R�����%E��H.�⟜s&�G	uI��;�	Y H���a�G%?9'���F�9;�`/}��;c�N�u���X6�("�pR/ίt�$�pD��`���ڀb�!���Zߓ6�||�a��S�$�Z��c��\S���<��*ٓE*��*�M=`p�4 �$��9d�X.0���N����qߺv�`�1�C]�?��~©O��Z�b�*��h�z5(��X�d���Tb_1C�rH�֫ցW���a�Ϗ M-�=c����j�~�?�)�{�@ZeD6��/Q�ވO6R^�K��P��h���	=>Q~� �n 6��'Iǖ!a�P�S%G���H�f�C�x�~d	2��%?S|�����'j����hN2J,H���<b���'��<�0�E�`_��&���o�B$@�'<`��9���*xB���Ȟ.qh�Ұ�N�zR a���l���:�Ʈ�0>A�K�x�I�����P�06IV��~� ��<dH�j0K�����e�<A
���3L�f�koީ�D��D��Qi2P�\n�G*+�Of�5ń'$e��₃�c�H��Q$	B�A�1/��d	'E�0 q��5��O,��r`�+h�����7���q�'��]ipN�s�~l�'Z�E��e��iflĉ��,��	{�.�;�lm�f�\�� R&[5* �3G�ߴ&��њ.u�\���;v�UK�X���&���G�����$�Z�T�����m��1
�y�`ͼV,�8��,��^�Х�&�������dy��2W.�7��Ӻs6��.u�ܔh+O�+g�Ϫ?���y���E.X���'���h&��4��t�rb�,C��0P7 �4��]Hc���A�n��b����ɹc]~	RD	���1j B�&"?��X�#H��''��W.>�p�'�9 e��9����W9�)ѲCJg��,�p���t��d`��l��;��vz:��O�O�* (ܫ@ࠨիP��z�'�B\�R
9j"X�5 I�Mz�)�OF$��+�����<��!�`���b�F閹�"O�����X�	�ri\�m�X�ps"OhI!�/S�5?��B���2^è�Y"O� �)�eK�F����"I _.p I�"OZ(!�	Ӽ\Ȉ�΅1z>NP���ɧ/��)A�O���wj��ɖqBG��ft���'Q�Ѩƨ3�PZ�.�"-�d��EQ8�`��aÍ%��)��x2�$W>w�p�@���OH��!�=D��ˡ��s0� m J����|���a���
ո���Zx���fd��b(&�����_��AQ 8�O�x�RO���@h���F��@��w�����gB
�B㉚�\uP�omZ���N9��Dj�v�8,'�,81镙�DE ��t�S�����~� ��gҤ��m����R�<I䣇�F��컃a�aXݓ�b�E:p(tN�=<�� .O���:3��h��?�	�i���;p$�cz\XT��=a)<���byZx$��`*8%�޴9�4����K�r���	w�/A���zڶHWi�vݐUx��(��4J`m��� HZD� /��� ���*b$A *��f�?��E��$�hqG�P-(i���%t�	Y��ތ	��,�Ɠ=�DЋ�hH�U�B�#��=:���ïļK��Ty��O�ы��i|b�iST�s��s@3�&M�兏7��)yd(�2u�b�w
O$ћb	"�l�
R���v$�x1��b�0
`m+&�<HI���~��Q�i�R%�
�w��C���YiE�O&Jf!ۄ[�i�`�?OJ0��Y�hza6�B�}DMJь� l�T%(a�5`�<�u$���	
��	K��"�2�B!Pv�)�ʇ?'m��b��_�8Hv��>�����>�1 ��x�Tݰ�d�4Y.�?+1!�*\�u��xm��gP�a�n#r�E��O`���\��CfV�dj�q����CS&�����>lj�h��+�T�q��)>����%�c���9�aC�A�5���U� w�v�Gtx�|z��=cV@"Fe0cVv<��C̱ ʶ����dZ�0k�e�o:��=�b�I5m�-i�M�O©� ���e!�E�-dǪ<	��'�6Mȅ,��)�rK���:��yBF�5Ɏ���i�HP�F�jeqO �h�Ƕ4��X��)3���Q�H	e�ؘ0��Ͼa��ɞΤ�q�d�{͎����л?���RU��s���e���t��$ܮV�\0�gK����8�H����'�����A(��P��F��3
h%J,��bM�*o�z3�7�SE�tdBMa�bƽ<��	���8k27�L�*$N�����<9���%�<`��[�m��j6���QP^�h��B�(��i�@f�e��{�O�3 
n���bӟ�v��;H�	�4���e�x�B�#O$a�w�-J_���A
�Ǡ����(g9�-�ׯțt���"FFG<��'�����*�(Q�?�ju�J�R>�!I�'<����5}2lR�M	t�
�T��Aic��q�O�<����͵u��刅�^Z�^I!�ә<��X�=E��'��+�Kͨ3���y�c��2�a(9�ؘ#��ܟqP�S��;��h��'tT�ݰ7�&�*��!	Q��3S��8g]6B≪H��p��~^�ӱ��D��`	��~�|��%F"[��U�rb�7�Ӽ":.��d�Qv��pB�<<O,���Sr��hr� �M�M7�������;�jr"T�<)A�J2�tt���Z ��<i ͇5[���
�
[9P�(m�ׯEqܓf�����i<��Q�$M�w�ĳ�pH;w���d�0��-a�T���G���x��z��)c��ќP0x"w�Vn����>��,�Z�oڿfI���]�^����l���L��D��( Y&B�S3�C�c�1w�@"v�V�L�0E��34�(#�A�dy��9O���eǼ�L���%�"��V"O.Ż�e�,)����$��N}j��%8OR٪��μH���ل�&<O(�ʠ ��}�,�:w�ă/w�9Z��'&d���P�9D}p`Q3����Us���,[o����#�>��� R��"s"�oa����팦u@�a��QH��#XAi�Nߜ%�t��!�D9�E��&wT��#����7�r�1l	&vP��GBЅ!����O?��D��E�o�&���NԚG!�F;:Xph��K��$�M�6�	�O]�m�G`�L��İe���i�T�S��Æ7�v8���0D��B�2��c5 B1L�F`3�:D��J`f�p`��YF)T{�`4�5E;D����#l� ���QX^ 7�8D�0��DEDsr���+�a d(p&-D�� �
,;`x��7�0���*�
%D��(��ȰVM�`g�ߩXnf�3�o"D����AaَH�KP
U�.�p�<D��+g��$o1O�m1^���;D�� ���n�;Fzt��eX�I�x+�"OP$�'I���1*	X��|��"O�����QG�r�1d���[�U��"O��9q� `3�a��6՘�"O�`�aA��&����
V!KZ�8X"OH��7�6{؄ 𤔴H@H�0�"ODZ`�D����*�cʞWX|�@�"OnmR!*T72���H���7Zx:�"O��C5-_+���pM�!7H�h"O�LŇA�Glm�,Z�m;Xy�"OJ��(A�la��q�!��
 ��H�"O��:��W��x�NȓT�
\�"O|a� g[��6\���D����k"O�q��e��5Iiҧ,��	�s�<���̪l�x���'�*{��@#�w�<�!��M6q+� %f�Y��JJ�<�$��<�5�Kr,�`��C�K�<idmP���0��w���NB�<��cI�I�(�2��L�GyPh����A�<'gG�Xxmce�c3l��tj�D�<Yv(�vW�� A��]DW"96�x����� ������� ��֓4"�쨆bF<,4�����7#
��ȓla��Dd��P�,-��k��EbD��$�Bt0 �C�Q �jS�Ư^�m�ȓ��(IRng~�|T!�b� �ȓ;��6�вT�ҵ�T<P�J��
�' �(x�!�>n>�h��U5L�P�
�'p��CU`^�DK��V
�$N�,�
�'���)r��&L3��ф��Jy���
�'�n<�G�^�'Nɢ�b��.��
�'(D �������u��q����'�y���G�/�d�"
�%��m��'Y$	���ͼ8ÂgY,�ftc�'��AX0.�TcH�Z%臩m����'�:� �fQ���3�*��v30�)�'P���%��!s��dE���'{��B��܃J��-��ϹS�Ȉ��'�z�ˑ�)RN<`�C��]�Ҭ��'��Y"���CS,u�"$�M�s�'+�#�h7pŲ�Z��ͶK�8e;�'Lu�����V� PK��1)8P��'���R"j!&�6��'y`h��'-���ա&5�m��e�#2��'g�0&- �9�~@��V�a
�'=R��qf�C*�	G�+�d1
�'Dl�q�ɖ�&�ҙ���*v�P�Z�'�9h@��*!u	ߐw}
��'*���0	O�	�"К�.O�D��	��'��8��J�dYXa�cc�A��`�'�=A��?s���c^�Cd$��'��IҔJի5;����l;2���'��Q���w�18U ȋl��!�'VBx��cQ�tU���)�_f@�b�'�>|�T���V���� �nYH�'D��TǕ
>4��o����'���$��La6	P@������'ިD���݅���`�SLlA�'�|��唆%q����=}���Y�'��J�مH�L�zCG�)A�D�'� `A�ǜ�#GvE��'I�'���'5^M�r-��s%�����8J$aP�':�REj�>|q@����!�'Ax�E#�ax�K⨓�}E^�1
�'�^E��D�V�����ѹp�(�y��� l�+TMս9���UHX$O�,d3"O
��A��&�X[�E�~%����"O��%B�-��b�c�����	3"O���h��`8�͙5?��I7"OB�7�l��ګm��}�b�(D�\��͌�(��(��d�Y�H�b�+D���!,��fi��#.س�X8�R�,D�D��N�7� ��ԝ}�@�i�e/D��c�ƚ��a��.�#Ej9*�+D� Z���GRR���L3r��U��O)D���ɘ3X���Rk��X����b(D�z�BGx���S#	�k����$O���e�h�(U�Ӄѩ=���H�A��n�V��ȓ��dbpLπ�hr �u�N��'��!yQ�B�S�O�
(���B�:�@
��J͚�h�'�
�Z�萰=�&��ΜA�-+�y�ΝE���㉦D����aȴ�.�b�+�y'fB���L��D�֥�Q[᤼i�!%�`H�'�FdA&�D2��|B�A�򅎇�p<iL�65�qOt3�%�jC@0�vLF�Y��`�q"O0(	t�^�<O|H
���M�h+"OR@�g��c`�uZ�+Ι����"O�-w��W��)K_�r��u"On�� �\�@������=(� �"O��إ*�R������C �z@K$"O� ��.7�-b !��!�<(��"O�Y@΄�h��C���\�bx*t"ODI	��W%r�Ҧ�7���"O�d��(ןZ_�����5[\@p�"O�`S�^�=4&];�D�C�0`"OL�2����	��"r�bs�"O���?Xa��*�JF�P�^0���O��Js�6�O�y �$�
��qUJ$�=���O��=�O�lDZrT�Tá��7,��3�/.��Y��%D� Z�m��A�����#^�ଋ�(�<aH�d#� /��� T�x}�8 oM���	ǈ�
�y1�0V��6a��p>YaFˤQ��l�5�T�,;q턶x d�B�S�kW�$x�!��WWNi��Rh�<T�r�Z�S��g̓���Y'm�)�qSG�?\_�)�?��%x$�F�T�9᪟��$���� $f4%��<z`I`Ǜ<{�!�oV�B���d,n���0��
+��0��,�",����N�該�B�KL�V��z��`���f����/K6y�k6�rB�x޴0�k�d��TkB-�b��Cߪ4	%���<1t�a�nO�A�.�`^�1ؠ}�f)�E�ayќp�@��B
��6�ɺ_����LsV�`�g�3c3�c��b�o�#�����	ͯ`ذ�0o%�	?p7H��ы ��hAm�BOn ;Ԋ,nZ�����1�z§�DK�T?�� A�G�*�X�)֘*���H�K-P�|��V��%hazr�"-��9 o�?Ha�a��T/4�� Ц�#0p����'3\����k�vp*ӎH�E����1���p?�]S�>]B�&�>m��5
�d^�Df���A�gs�%X4���
(�B�^'}ۖ��A�v1�	˓z�,3U!�:P�`��S!eѨ�Rg葔O�5�DM�A��0�2�I=4��X���i���iP��>�'�F�CǉQ�e;"
weƹvRn��O�D(�ڬ3m��b��?h80�d7�	�`afu�)�"o%����N+�pnF7P�-�R�Y�+i�A��'k�-��K�c�V<�U)�:��J��h?$�;�e��{Ra�&`-��,,U�.,�V�������d�B3r�Ɇj'���1)�[@����u �Yg��t�f�(��G<�$�`�-� %
>�)�"Ca��x��ŗx�)�����L�x��O\���*�l�H`�k��]��֝�<i��M�B^֜�a �rI6I���X̓/Jଐ���2E>Js?{���O�}
��#?v,���M�U���V��I�CG�հ� �d�d�KE�4~7�u:p�L-[���CRF��az�n�b}v�Pb�?t�I�EO(Uh�#�oǚ@���A3��5vkU�Z�:Y3!��u��Q�&d��Px��K�t��Q�` �]���$��F����'�����F���� ��.?��Jç�A�ůC�}�JgBA�1"� ��	�N"�{"�)EƉB�� 'P� "U��8���A�A"4�F	[5�>	W�� ����bR�J�P\Z/Rt�b/*��$�D.2θ�q�V:����Od�s�뜍B�p)C�U%Wd�ʡ�|��T'S�"ԁI�-=�hC��!�|`!R=H���7��0>��S�v�|�R��8Ԥ1�(�+�8j���
u�N�������2El�/O��?��̠�̓��倻~�p�j
Of� �ǥ{��0��	)�Ε����%L`x]���'���ra]���iry�)/g��k���|jvnS�-��g.��8I&)�~8�p�fL��DZ=� E��z���PJ�L8t�a� R�,g�8I��K�T`�Dw��vΟ�Th�KN��t�=��kN�E�`�f OHސ�S���u�I�V� q���+�t�u��=lX����
�n�¹�A�µ7�.���'�K�����!���p?Q`dËa�j!b ���&�BL2���	E�6���F�xjV%�D}����'c���λF�t��͵;�u�l�8�6q�Ɠ �N�1�b/u�D+A�L(y�*���L#j�I)r�B��Q�V ��R���AǢ�ljri�3�l9p�!�x�"%{� #<Ol8r�)�8+"$y�ӆf֜)"e�$.�0�T�dG�p����b�l��[o�ZTKr�>��ڵ ֆ��<��I9*ak�Ɂ#��1QP��W�ɡcw�0ST���
����� �6P;t#e��|��e^p�$�� P��Hc�K�1q-O�`"�#^az�����̡0&�6ʞ��Ƃ��Z.�aHu!�<J�la���Kl�ب���tW�T?Y!E�_SW ��sb�#�ص1`"^�)T�g��r�<��:������_T��
�[����a��=0��H�On�p���~�� ������ND�������,�@�$�h���"ONx��J_?P�����oð8�� @�7Old�@�@,82���@�<��LQ����<Q���I�<�(�$ǊGIT�KC �R8�(�įD�|�$R�#1@˔�{t��B P u��,����Z�C!,˓C �@�^b���Y���9�2 ��c7{�]j��<�l��}��rp��j���)�J�Ϧ�?Y�` ʮb�0؁Ίbچ5�w)?D���ӷ�<�����٪7	�@��|�W�C�Yox�v%��S ��x�&���B�	&�������fz1��/<�O�D��t!v}	ӣ��I`R]�gH�0KnϧP��I�ڴk����D�GG䝹$��&��9��`S�Rџ�qꊠ'@�x��β-m���j��4cB�Fn��	��. �oZB�I�~���֫�";j8C��\D���%�T%s�&�bH|����#�:�T��5{��`C�΢s�C�I�T
��� ��ĉ� �<K�H�K}�,V�H�������{�Ɯ�<�t[p̞�eb����dS���?	�΄�\�Z0`R&d��HU��>Ge8ёƧ]0c� �y��P��'��u��K5 �3C$�2�n��`�"���)b)�II�!۔�
&��B_/
�A���'�&�y�'W��`k�O-u:��J�O�����M�:jt�'8LA��8��Q��� !�Y�\��d�\"s˔B�Y�@pÅM�*�$��'�"�~��O���V0%���}��+9?1�&�r���cQ=Z� sp@EI(<Y�:�+c�߱Ү� �a� D�����d�L�xR�C��	K�W
eX�xeE���<I�	'���?�H�3�
:�\e�1kҦi�
C�ɳ,�Ɣu#ˆG��Cf�5eВO��A����']�B�ខ�<��aŲ>X!�<}ܞi�V�# ��$ɀ�U� K!��\�5Q8%Xł#�
�0�lL!��j!\�֋�z&��9���U>��-�	F�j����%��s�dȁ+ІM9� ��W��u"O�]j�N����/P;T��AQ���E�?y������'Rd=h�@� ��%���!��0�@KZ�!�F��%�)�P/R� �~h��*��u۶�;4�����S���\�@��%pP���j'ғR3��!w��]P>�?	ڱiM�F:!�ƢԿ!�.4Q4b&D�scl�0��IK�fR��#l�O6�@s��`d�Q$�"~���Poe.�#F�+#��0c֢�y�j��n�Lk�G�d)������y£� 1��1�@�c�����b� �y�mѫmW�1�X*XX+q���yb/.+�� 6	K��|P���ū�yBiW�/�J��&�M	H��B�y⣎�l�&4I�Ꞝ���y�����y
� h�T�(�$Z3�P�#~H�@"O�ѵ�М[����_!��'"O¬8��2LU���B&`��5"O��� L�bln����ϥT���*�"O@����ZIj���A8t���"Oh�Z�hJ<ed��&F�V/��c�"O��覢ćt�Ɯ`tKܣy���"O��[�#�yqۄ�X.���{"Oެ���.k1�шE��4��dX�"O�H���ѥ�|��F	/>�n���"O ��֤zI�	�א$�� �W"O)[��Զ�:�ɧ�ψD���*"O@��#�
��~�c@b�)�^=c�"O�(B��8B�lX5�Z8-H8��'
��A��_�P,|y2��>z��A�	�'S� I6���*�T-��j��j(ٳ�'@ԍ`�CŶb²�r�-́fh�Z�'�vͩBFǋ1S����� �ĸ��'����o��BnYAG�
I�T��'��Pv���#��E_���'g*���i�da�f�ŐN����'%�{�h��e��u�5�@�=8����'��a�A�N2wަ�c��3 *���'G���f��XU��@���%?�����'��}0�A�?������3�6�8�'�Hb��[����W�Y�?&J��'&�a�f��K����F5A�(��' ��[���D#<����p���'h%�e��UV��y&�W`"PК�'}��s�̨"�-a��Yv���'���6��7Tϊa"��U�I*��p�'�JLkc�]�/ɶ�[ g�L��'J<YAU�� E��Z�ҀK�
�'�X`ud]%��y��/�2o����'��#@��:=�pB�)��a\�I�'+:���#�$W\����
Հ.0���'�ج���>9�f � ܢ%S���'��Afp�['�ޣ펱+�'Rѓ�+��0<Z x��}��
�'B:a1��V�F*��7�/xԆak
�'����Ѹ>�5��g�j���'�=+fC�
.�럸`�IX�'6f= ����:H�HB�	�R�"Ś�'�|�#D9E�j�0���$ �
��'	����KN{ �`�(�!%1	�'�치d�M�_��5�� \�M��'1�a��H�|L��(V�~�:��'��z�$��Z�����IY�u
 )��'Œh�D�M�d���eE�ov	3�'���p�(ޝX�@H���n��41�'*F|���9_2�(!�C��a��}��'���p%�������`�] �'U����n�𨳑���lyNM;�'=Hi���9�
+t���nɦ	:	�'(<Aq)^�qڀ*$��r�
���' �� ��#sb4i�ޗ�İS�'vLy �̖;<Z����X��6={�'~�kw/��i����$gR�ʓ?'.�f��x$�8	���5H��ȓF�|	a�M�3�L(�3�/j����A�6@��-\
Ku�D�o^�B�z܄ȓtL8��� �|���abS�/�,Ԅ��b�c�哜qr�#D���6������J�s��0åw�J��S�? ��ࡨ�05o�4;w��΃?~E���]*�D�B��H1+K?4��ȅȓ=�����ș)7��@3��Ta��h����Bm�'x��p	?Iq�,�ȓ[�t���әT�z�*@��#_�!��>Vp
P���Gpn����+TPE��\�,�h�!�T�,�E�܁��X��#��!�G.�����6{�L\��V��yyP(=���q,b�ɇȓ!|Rt!%���5���c�/��C䰇ȓg�r���$h�0�3A�F�>虇ȓp4���K`Ơ3���+���ȓQ~vt*��˪o��K�_˪͆ȓ%p̣��A��\tPᇋ�P�ȓLU�Y!0N�&Q���R�\_!����o``%3��ē ���G�v���Y�`�
EA٢2���j�l�9���ȓ茰Sw�۞2k����!�p$��'�줛�/�
%�P�D�	VT�[�'��p���j�$<u��0N�����'�l{�]�Lt��t�����
�'��3�N��FP:y�dmW��*	�'��5�Ć���T�D�Ǳ;�	�']����&ы|4�9���-~��X��':0M��]$T��C��v�8�@�'O��BWL�S~�zck_�qg�

�'sjŊ�A��*!+2���n�X\
�'M����̈́�(����P��И
�'*kG��r�T #���
�`h��'Ȱ8��͌`����dg��6���'JH�l^9(l�I!��?(���v"O��:6aU��F]͏�r	�4A�"O@DZ�I�n2Đ�:CL���"ON% �kF�d�T �I*>UT���"O��z��8O�ua�T�snҬ�""OU:�f�9Ede���_�ݠ�"O�Q�#A5�D��U��#�p��"O|�!OH�*�T�d��$#��)#"O�0����<7N�`�]��Mҵ"OJ�aV�T�7Q�1Sf�'&ܹ#�"O���-�|�E*���If}ST"O�9rt�+0�x���oC39��"Oh���Է^lj��D�|F��"O�P��� 3�V�I����`�4"O��U� �1�j��t�ˈ`3ܸ�5"O޸��LL;d3���tLW h F sB"Oh��*9k&��W����)"ON��K"B
]�dKK.b7����"OJ�MG>6�Z��2j�J$E�"OH�Q����r��(ȃ#��Ļ�"O��{�瞤�P��(�W�L=�"O��X�A��p���N ��Upr"O4���CC)g��쓣�4,����"OTq0��4����F끄.���"O�Ģ�E؉{#|�9C�	�<ta�"O�IC��7� K��[EJi�"Or�H���<>MA�B�U`Z ��"O��!�g�.��[oûNFM�"O��K�HI�i_d�6n��Bk���"OH�@A[��l���K�q>Z\`�"O4�Q�'2Qi~R��!O}��"O��F5F���M+[3���R"OH���K�@�mStB]�U b�ʧ"O��{EOʢy�bt3AC�8Hf.UYE"O� �82�
��
�0d2$��7`53�"O�$�cI�;G�	$�Q4} �"O����K-ÄQ#��4��䰔"O����C8]n�|�竞7�$)xF"Oܐ�.D(@����J�23��ɚ�"O�Jg� �D��A�JL1ϲ�a�"Oz�B��	�OR0@�$ȀR��9��"Oha��b]�x$h(c��u��Y�e"O��#���y
� cg�\X�dD0�"O y�AiP�Wy6�	�!]�0���#"O�!`�� GIjsAH03�����"O��{T��Y}���� ��+s���A"O�A��& .ш�n h`p���"O�8�#&�c���cm$I$șq"O��B@(H4�â��D�"�C4"OF�8���P�pp1�,V��jP"Oƅ+Tʋ3d����M���MQf"O�L���_uKne�������"O*�R�j�8Hs|�SPE��Q}�U"O�TJ�g��(�rA���ڷG� �"OL�xa�'�LL:5┒/���4"O��`�`!h׊��a�E�6i� ��"O��,�1!aްa���6
9��"OB\#�/��o:tK��?#X� P"O5:�@�7l�V���@�#H��"O�,�&c�"H���*�/,��	ʀ"O*y)s.ƪrqg�E�Z��"O�EʃX=񾽁��]9<���"Oh���S2^7�(���Ha�ĵ�"O��B�D� �P�y�Fۯ-�����"O��fP�p��@���N��:�"O2�����DM��10�ѽz��5ۑ"Of�Ȕ
ϊG3J!�V&��"�4�P�"Opmޑ'�f�*s p���q�'��_� �P�EG��tat���wj��!�|!6�H�9�I��K6�0���LG�h"R�ۛr�����H�]�X��Wc��W��	.��h���&J~ч�gn`���Dl>��x"�GS�ЇȓNb�%P�K��>V\ȣ쑑����xۂ%�!��{�MX&�\�����fd+�o�p ��Rt
ڄC�.���)�N�ȕ�_�L�*agȕlBt9�ȓ�8,�r�2���T��&чȓ�Ը��GC *�y�"��s�j��ȓ}���B6OɅk3|��P�,4�\Y��^-�a��d (�Dc�+�6���6�� J�'Q���x�k��`�`�ȓY��US@�F�
i�T����wװ!�ȓ~�$�xĦA7vݺT�P��q?.`���(��g���]�=e h�V�E�<�Q@�9�2��`MW�MD�x�HC�<���rD�*d�	;_��ՋfgVA�<��]1;/�5A���S>��2�� Y�<��E�K֊�0a΁'��]{r��j�<Iu�
{N��'�zt�ʣD�{�<��"Y�eb��53����'�\�<	SÓ�KvI	���{�h�	��UQ�<a2�T;wu�mS�*�;LVA�\r�<w��<c����ɮ<�4����X�<���� ���F-�vk�����ZV�<��͔v���ӡI��C�be�B�NI�<q��˼��1��n���(�@_�<y��]�:1��KX�3�\�R&ED�<� �A*�ܞ�B�QS���3P5��"O> P���8���)�{Xq�C"O��+CC��torl�)�-�M�F�8D��x�	�<�I#��́m�`�!�6D�ܣ�F�;/6r�Y�͊s��j#*4D��6�J�=����@�!	�)%h3D��ʆEY�^���8��J�(:��&D�H��
\ BL:���&>�i'c&D��v��V�L9Ǥ�>M,�4C&&D��)�j,e��ؘ L��5f/D�T#q��!�,r�;D��ȃ�%;D��5��W*4E+�b��e�|�+R�:D�����=_�rY��M(#>�=�3�4D�`[0NT�u����R�F�*�K'	?D�t�VE�1ẐE)rR�0Pf�c�0D�T16=v8�%���q�l,QU�+D��3�Ƒ�1���}Fd$YC*D�H�vKֹ�8�éS8'�((���(D�(�` ���١BS6[�@�T� D��JU�I�j�4�Y���h���J�J?D��0r�8y������'1%> ���=D��cw�E-d� uNT�r�
 @<D��QZ�a�x�JS�=��  �)?D��8���#cx�D����J����;D�d��΍�hP��(�/�4 ��,��h4D�D�3�WA1�*�*O00j3D��5@��#/��ѓ��R��q�#D��Tƞ;^���C�,��mr�t���6D�@0��5+a֡;ѣ�s7���2D� ���A rp�N�9n�愢�0D�AS��H3 ��&�\�A�t�1D���4�̰O���1�O��*�[�,.D��;�(]�vY �,�vI�p{r+D�����"7T�C# �7PL�2Ũ,D�x� ��$��p*Pc�4Uv>d�`'.D��2��ǭtv0��!G�owK�8B!�䅴v�j�cpL#ZԪ�Yv'!�D��Z��[0��)x��f�D,YE!�T:��`�2�X�m�K�#S��c�'ˌ9���P	�6�x�o�p�0	�'�Hp�Á�8|��i���G1���'P�͒�O}2�l9c�9��ܓ�'|bx�b���\O�۲+׳2�0��'.��
Ä�=t���B��Z����'�d�8�"\qu,9+���<)�D3�'��TQa�4exX��U7���'#`��O�8l��ᣐ�B�N�(��'���#W�|h���	�N�J!��'�RPr�X��-�e\�vP�H�'{�-�)U�6^�soO>�0y��'\r R��Er��"���O^���'|0ATg�'sz8ac" 5p�}�'��g/�@��Y��Ԓf�uy�'�Bm+����W�P]ۗ���3=����'���-�g���@Q��b�M�<Q���7u�^���aV�H����N�`�<�H�I����Ҷ ak���Z�<!ւI�<F�=JU*=`�����Z�<4��5�`�� u���C3g�[�<�4����� _�Q�лql�\�<�pɃ.XR�k�jF�,�v8���Ab�<�+#4�<� @�=>^�*s��_�<�6� 0G�	jm�� �e
�Ϙb�<����1j��*��R��$�G	c�<� �����6� �!�"MD�&"O��d�޴=���:�nS7@��]z�"O�Q)3�ʓ]�Ƙ[� �md8���"O L�rn���d�$㕭_O�]��"O|��aB�H6%8��N�k(FB"O���mڢ*	��Y�K��U�<��"O����*:���KɅ!ⲽ��"O<��N��x��sJH8��,�"O��SF

R^����H��H|�!+c"O`1�P���BD�O�wCj��7"O���ԭR�l�h!�Qw8�]a"O�,��U ? HD� �7Uӈ<��"O���B��tjlc����.nr�@�"O6��W(��W�l��ԣO�m���"O ԢpfRD���C�(g�@A�"O>�H2��1|���O+�zK�"O��k� �^8��٥���B"O�(c�җ.ʂ����<]��0Z�"O��!B��8]�u"�{lT�z�"O6�i5j3(�il]9Yd�<'�'�O�Y��I��
�R���$SON%�"O*��Q�F^9g��D)� �s"O�D�l���T��^\	�"O�q�G,1�� �mQ���9
�"O���&)�/Y*(�H�AȺ���"O�� 2�ҁ=>"�б�:]��R@"O��h�Iܽ/��KBm�,x�U��"O�eCD2o�M�5��Pi�p!"OjH���?p���h��L<YsPIX�"O<;��� }�`X�b�T8�b"Ot�`��^</}v�r���bbn=�!"ON`+s͒)�h�(�g]�;2Q��"O��`#'�{6xxy'�%;؄���"O^�)�cR���!�pe�g����"O�ۆbΫ��y�vc�h�8�s"Oj��nF}���6 |�Y�"O^M�W���x�nXc��
5���b�"O�"� N�[���o�" XJP�"O�l1�#��c��1(�O=���"O慈�.<H~��G_.I�D,�3"O"���k�3.��Xf�XI���Z'"O����MB�� �?FZ��"O��e�L!l�ܽ�Q��;U�F��"O��&Ē��A��L'ho>-��"O}�rN�u�: �%!Ƶ0��9ƅ04��+�@�,�EukB� ��Q� M7D�Kv�ɒxr�+���օ�R 1D��7-1u\��	��_��]L.D�p�B�B>�d�t��E��!�� D�2 �<I)��S�K�>2����o D��`vm�arx0���4&�D���<D�����W�Q�\d�j��b��;D�
�#��_��XAE�C8g:�$8D� �b���
D cnܷCc�pq��#D�(z�O�53�dp!B���R0;@B"D���gަ|��#BI�I�d� $D�4�%�=�@=��g
�gT���&}B�'��z�-�V�AP����T��'�`9A���)Jh@WCɄ�vX��':,2T�WXܑ�N�
z���	ϓ��d>?A�S�( ♢Ь������a��O�<1p��izN<Z���\��+4�g���':�в*Q�Y�h�r�G�f挵@f"Or9I��Us �=���S�"O� �]��)̾)Rׇ̎f�.�ɡ"OrHk�LZH�Q
�'Y��${B"O��A!A��\��9�Ɲ����� "O��A�I*�@5���k}6"b"OT�$ۅ8��Y�%��H�Q�#"O"Y91NK�/ym��C�<i�.���"O�E�/@h�D�Jw���O(Ҡ��"O�"B�
}���r3��nr��"O�@zKЋ4<� �7U�n��`"O@pr���j�ڐ��B�.��0q"OF���M�CZ�X�r�_1�DD�"O]ǁ�|���QF�CА8�ĺi�ў"~n�7p�ZH���Ȫj����afX�_3rC�8/�bɋ�]�t(� V��dC�II���h��r`Xড�0l;����"}�B�J�)�0��YdO�y��Ф_��p��Q?�������y�ڠ1ʮ�C/�����ӆ!�y�@�Lv�9qNN v8�R�E��Py��[9<����Nʻc4�`C�i�<q�#
�&d���m�`���`�<��N�TH�/��t�6�H`�<�7c^7�(����&�fI3��^�<�R�[[^�X�#��W2|#W �Y�<�1��r��#���r���K�<9�n@,n8� I!E֛`a,�
$EF�<��M?M�*HZ��0xZ�i&A�A�<�*܃aRF�nX�r���`���yBj�Sp�hhG*�q	Ĕh��֛�y�ʕ�	�z�y`��6-V!;�B1�yb���9����(X&PA��J
�y� V�]� j��-�։�o%�y��W�E��}�����
$�[�F(�yR4/���W"V!�4�2
ֺ�y�Փ2�|����61�0�+�ǖ��y�Q�Dhtmb�;�2EK��yr�\����%��a���I��yb�Y�k��"��F�M��	T��y��Cz^-�ReҵI�`��aT�y��I@\�Sg&ݨ=�p��a��HOz�=�O]���ƌ
/k�|;�M�� �$��'u��7)�lՂ����N�(��mЍ�d$�'%�@��@FԣK&�Q��?�昆ȓ �D��Mտ���"�(8�Gz��~B���5\��X��W���8��X���O�"���ui{��Z��� %>4���R���dHi�j�3;�p��&D�Ш���&{�8��!���$(-��
*D�DaL�^���㐡���ٲ�(D��0W*�4}ȡ�G�PM������&D����
�.����F��9FJX� �0D���@�� ���F�R&g�
@&$D���'��7{���c�N	;4&D��`������i�2b$��/D���g�5TR�l@���:}�,�#n.D�P�b�M89�h�pRɌ�3�խ*D�,1 �˦o�y@���	%~r�eA*D�D�'�����7��&n4Pƣ2D�hg/���dIuj'�,Z�'-D�H��U&4P��
`AǷ�ѐ�,D�����ݨf[
�Q�C�%�Р(g 5D�t��	B�Tq��k��J��8(W�7D�ȱ����`x�X�I,J�v(��4D�:w��0AR�Q�c�.	�JR'0D�� �Is�ʨD^2����%����Q"O�R@�)���d�S ���ʑ"O�:R
W+0f���c��1X��LH"O~�"�.[�W��I���	%�6�c"O�2��MNw&d01���G�x��"O��i�20�J�
����>��"O��zaG�4��"A8[��U{b"On��rj��[�4��B�C&v:l�U"O���ր�)6g�u� ��>~lI$"O�R�N�F�%˥i�+lO�k�"Oj�1�o�Hz̙� )F�"F��x�"O�U!��םc�"�$ �"�4,�!��O�\�P�,I��QY S�!� �x��P��莴k":(ĈZ�=�!�QF����H�2 �c�<l!�$]�5�D�{�D'��QZ$�PyRLL���9g�M [96+ "_&�yBS�{a���K����M�y*MZy��[�cЖ������Ҹ�yB�J�^�d��"�3'�ڬ�y2��3�<�b�բ#{�����yꟵY;`��i��xDyK$�yBI��Z�\mC�g�	�a`�M
�yr��zU���sE�zr�g���yr�S�l^>���j!�$�� �9�yb@�3��Q���Q0hn(��8�y2a�P���UDBR5��d[>�y"���i�`0P���*JZU��m��yr�\Έa��2+
� �a���yb�6�X85.�5Kf2����ɰ�yR�D��v♢N8�}���Ҋ�y�g�'oC�Kv�<x��5�j��yR�ǌ����##��{��e��ܵ�y��Tr�Y�T�ݾt��h'�ވ�y"��6'�=X ց}��@E�σ�yR��iU�$h4A��u@� �,��y"lR�{G�X�ETrpnM�b�9�yb�W�2��ignr-�׎ã�yr)�����A�X48�Ҝ���"�y,��V�@��f��3�2M���#�y�(��	��Qۀ+���P/��t!��M*q��5A��)C'�!0%��v!�� f��������1�Y-$�!�d�,{��y�w*����ۦɧo�!�$��,��}�)�|�:	�k�!�$��s� ��p/�"wJ��t�L�
�!�dÃ_��k��37��kTdF�f#!�C1p� AA�B�(�z�u]	7C!�d�nM�Ap`��;�n I �~<!��upԡ*�`�5#���3!�$�d���H�BI \b���?!�Č���n^I�`�J/�6�!�DL!NX|5� M����T��S+e�!�d^��LdS��I1S�x�K7���!���hۊ9�ݦG�����#�B!򤒫BN��#큸~l��+R�+�!�$@'IC���j��xAe�J-#�!�$i�0K'��#���1d�!� ��R�pb]=�:���*�2�!�D�L*���q�'9~z�I��d�!���2��qʁ惜"oP؂#��G�!�/2��e��i�pTĵ �̆!A�!�d@�����T2=n��Q��<�!�[9��"J@YPV��ծ��|�!�� �a�%eB%BMd��gAީ���+�"O,9q@	#d&P�i1�uź	:�"O��Q�$ڙ$�<يc�a��ib�"OV��B�{耚�G��gJ���"O�� ��=dK�2I�.k��=K"O���$ Q�!���i�h��)� ��B"OT9��$� `��EF/<.��"O�8�%.ݨt	��r�#W�(ӘPC"O>��F̓?f�^�`�..���"O`�c�+H(xܚ����'"P��@"O�x�/.�20����6'����#"O\]F-�05f�H`��KPԼ�z"O��pdF<�D�#fݽf�j5(u"O�m���	�|��U��Dަ��"O�b��	K�\}�E�w�XM��"Ox,��/��S���V��Y�V�Т"O��S�H�&^|-�ǃ��gg� �R"O�ԛ"%�R�F����$Sf�@�"O�)�*�?�,���{PE�G"O�%�	�r:���B\�FO^���"Oh��	t>&�
S�I�7*Fu+�"Ot� Q��p��do*X�x��"O�=x�=��e����1� {U"OjI���~��8��R.v�n1�S"OtUaULX�@X�0�@��|B���"O֥�Ş�zێ�����aB��"O~096�F�n�P���n dyv"O�MXp��J,ۆ$��VS,���"OD�ʖ㊈n��u�u1'Ƞ�E"OL�JaB�+��L{���Q2�P"O�u��.�/W��4ZPLJ5u��b1"O"(R�]��`��I*+ �"O�U0s�T>�h�w�D>Y�,`��"O�]ˁK5{�lys�埐Z���"O�P�(��^��$jCFd�ac"O��0�	$b��2���)�{�"O���φ�S!��0P�}(��B"O2�c�BS;`.x!kC&_�n#�qp"OVSEdƺ��d���T�
�P�6"O=X�H<kb�*B �h�40V"O8 *�Á"Vf���o��T ��aE"O���D[���BT탧)�f}R5"OJ��ac�$��8R�Kȏb��s�"O2��0�H�k| �@�V"�����"O*����"3S�0ȅ)9M�\�D"O���b�)-��Rԧ�,E�T]� "O�9uM�:@JF��!郊
��-�R"O0`*Q��%;虢@�P�{cpS"O,�`N�	$�ɘ�E��_�y�b"OB��U&I�y�z1�`#��,v�ġ�"OFU�1�=YT@���N���g"O�aI7���^���aV=���F"O�M �b��pBɀ0Qh]�@�6"Oj0�!�dl���s̓�[.�$["Ot� Go3�^!jхT%n
ԭ�#"O*��C�ʋ$w0��6B+'�e�6"O
�!P�@X���F��P�A"O��+��6[(��%[)�
�і"Ote��3U� ������2� �P"O�e�e��/^��
ѫ/e��G"O��q���f�,J�ѱw����'"O%��(|��A�˽So�x��"O9��"�/0�� �v�
'^Z�Y W"OpqƆ���(<#���OP�5�"O� ���?W�re�L�2�(���"O&��Ȋ	ɪ	�*�4E|���F"O����bEo|.!G�ی@���"Of���!�n�*YT��@�<��&"O� j��^	F���G`&
]sc"O,H�%̈́�ajM!�摧+$�h�"O@�3F6d��p�f�>""`+�"O��:�Z�>���@V��2Is\TY�"O:��$+ˆr!H���'V��˥"O������:��t�CgҁB�x� "O���C0<6��� ���C#Nl��"O$\IQW.	��Ϝ<"ड�"O�L2���<U�V���c/}0&$��"O�t�4��`���Q�Ct��	!"Oe�ՏǜF!
����(-���q�"O$`y�O݋���8v$�$��y"O���āьL���8'*πN�i"OX��` ��ѹ�銕 ��	Z�"O�pp�-��2���(��YCB"O,x�bP������o�C�:4�"O2�(��2f��mAE$U�\��"OЭ���u���
u�I�)����"O������S=J��Cd�"A6pX�"O|}`���!���a"Ր�^���"O8	1�MǿKe���0L�)�Ei�"O�L-Y�bYq�]$RD�ц&���y���'��L@�/`�X�k�A�ՈO��7�' ���ڀ-O-1�<A���/iyм��E�P��e��=x�|cb��{����ȓU��0��M)�l s�f�]I��ȓ~���F�b,�9�$H�QT�ȓU�@�S K=�x��cB:J�b��ȓ��Z2@�"�j�X�g�I�N���ӊ@���2��7���U�.-Q�"Oްhp(C�$��:�$k�'^ў �	��9� �2#��q���;D�py���?Ƙd��� F��X@�8D�<(r`�3ޒ��W��ͪp9f�6D�̛GGޱnA
�8d�GzRl�{�H4D�@d��'t�	�����~�x�V/1D�<r&�Y���=�0l8� ip��-D�����`�DX�$a�1(( ���(O�=yFh�/w�΄`��]�&`Z����K~"�|��i>z6�Ñq=yXg%S;R��r��!D��X��	#1�($���U;(�T2�>D��2J�>�։�B��/�
D�4�7D��&CF.(�$��RB� ��e�7D��)q��O��#6d�+0��y�!�(D�T���\d!V��u�Ȕ��=c �%ⓒ?����S*w֤�&�#�f����OK���_y�|��)Z� 8���H�3���Ȕ�P-U !�D�(b��Ȋs/^*z��{E�5u!�D�%Q����L���ʕ��!�!�$�UK�tJ��7e鸥��l�!R�!�D�?8����A�D�h�]7~�!�$�%h�>����\�O�Q� D,vaz��C�@�Lũ��]Ό�KS��=w1O�=�|p�-$��q���Փ׎��eV�<�����PH�.�� 2>����[N�<!dpy�צ˒\�A�b��R�<yGc��bˮ\�k��jɎHr�'��<ɍ��?�&��ǜ�7�z������ ��Ӏ9D����P4e~�SbÙz���-7D�dʄ�[*�%�	;
�=�r핛)�!�� ��+�T�*����gO��A�����"O��QV �vQ�ܑDN��1�R1��"O�%p��R�^M8���
�I���C"O��r`(�)pD8�嗎 #Ba�"Ot���k��H���(@�D$2}XMP�"O0]�CRz� UAf�!"O��TKJA���a��{d��	#O���
���|����{fJ��D�3h�!��]����������O�D.|��ȓ$xFг҄P	�,�+!��	Ro�E��B��-y2móX��Z��J�XD|r��Wژ�q 	\�w�	�1�^8nvJC��=a��Y3d͇��i��!��=����<��Ο]�|��"�ߜ��q�K�y<���d� �B6+С,�d乃e�:�p�+�'[�8�p͞�U�dqP#"�)=�B��'NZ	 ���l3��86O� 9�@q�'"�5 �H
HǸm��+	,v��dK�'�vyi��@0���1!�8A�'�FpeE�����f�G�X㓅�*���`T=&��� �W~ԅȓ�z�	�M��=W��"B�x��	
�'�fq�п3#~��ud�����	�'���c� �G���A��䄫�'�x 1�7R�xPH�8q�r-��',�� ���27�jeͅ{���'�r\�jIo��� *"��ӓ�?YI>�����\�b'��B��A�Fb�<�� Ǥ&��Ibe��S���o�I�<�Qn��A�|ӖM:�0�B�a��<9S�K�H��AO��t�b�aJs�<�!Рh�0����JBH��3+�x�<)��9)jnhd��=#���![]�<	�ԴJ���P�!jD�c�L�W�<��*�W��Hb#��L��ICa�[�<i2d��FQny���<C�,I�F@�~�'��y®��W�*���L0:v 
��y2�"�b�B3��!�h��_��y
CL�P'��h`�3J�9�0?),O6��d��P<��x���*l�,As�'b�	�B���T:?S�4p��ǛbC�	{�X<��?5�z��!�oRC䉓-;\���	_�TB�'��HC�I�}�XP`��s`�(�!mMB�%C����iE��J��oD%�C�	;ik\��P�S�%A(T�oh����<I��z�Y{D�Z%�������T���?� M�?~U��)��5��ap�-�1��x�i 29��xj�o�?=�`�sQ���y��1z��Q0�゜_�Rp�3�E �yB)�*BɄ�{���#QӢ8�B��<�yR�F$n͒��tA��z� ��2���y�m��Lt�UR�N�m��8��[��y`�"m"��;!3\'��pg%���y����S�-!�˾Leb��W��8�OL�=�O��\p�9Q]�@���X�^Q̒�'>D�±�H� u|����%cN���'��r�D�)C��<Q���$gZ�A��'�����,��rw'ߊ	���	�'ӾU��m =V��BJ�K�i��'��h!�NV;��ti&-��*�����'n�H� ��k9���o����,C�'@VH
#`��N�$10fL�nQ����O�=E��` tFD�p'�]RŖ,��P<�y
� �5��P$\x@��׋P%f�Z� d"O�,����i"�=��sb�񷏗}�<�c��dX08�s�ڭcq�d;�BZU�<1� Xf�0X1��<��àHPJ��P�?Q��@�jք�*�ǋd��c�! a��hO1�F� �#��P8�� �˲CȠ��"O$�p(Q�x�N	sa@�1'�7"O�I�#��Y��I��&xp�"O,�g+U(jv��!���⬩�"O��F���g> ��!
Ж0�Uk�"OV�i�솀io�!D�H1�d�)��'�ў�J0BЀ���Ԫ��p���� D�t�4�K����y�B�q��=D��[���p ܔ��Q���@�<D��ځ%��*�t�����Ό�T�:D�,�`)��}18	8�B�<-��UK;D��AZX�!�"!i�A�6(J�NC�Ir����`�!҈["
]C"C䉋D�#�*7���J�.�B��hI�i���0�[* hB�C�I�6�xi��& a
���M��4��hO>u�T#�� 0�僧����f�(D�����8��@)3O*g��8uO%D�|�bhK/>��%&jE�'���:��6D��s�B�*G$P�_�}����*3D��B�		�j����^�Z�����1D�`1��<!���� ]�]�����0D�8Q��56��}�JY_x���]y��|��9OX�dP�Rsj+�J��v�8�d"O��"`�_�x]��(�"/u��r@"O����P$p��uK���&lr�9s�"O"�2�!��2��l���P`�B�34�h�E����&�IA�V��F�,D�0�C��?�����2E�n�&c0D��ԉ�<6gH��B�BY� U2D�0���6 Lv��G��.e�
�)`�.D�C���#3�®�J�YCdN-D��StB�i!��Ҵa��4��A���j�����$@5"���b���&�ƈ�b�;g?!�D�p9�5q�F� Uߜ;V��N�!򤆛o�|xǦ ���ar��
{�!��]i��X@4�����15&�C�!�D��YL>�cb*ЪN��]����w�!򄋊T�Yu��H�X�#�!�
i5&qzD�@)��Ƞ�W�7("�=ͧ�?���Í7.?.�� `H�R��,:'8�y���2'��6�����
�yr`ăN���U�*��L�0!��0<9���� �,��2�D3��G�^?n�!��r�V���\�%�@���ˊ^�!�E:��ix���#n�93B��u!�dJ�p� ��I4a�����GZ1O�|�?���ȃ�d�T*� ��I	q��l�<)C��%�R�x$�� 6.�TL�m�<� ��:=�f�pw鏇?QMC�nUh�' ў�-� ���_ڈ��[3�)�ȓhӈ�X��_ 8τq�2	�1|���4d䀆V6��V�\
%Ų݅�t��[ �G.0"��aM���-��
u��``�^�z��A��ƽa���ȓ2��{�kٗ�R(���3 Dr!��a��&̙SJU�#��{N"�E|R���R@e1� ��  I���=�B�I�Hv���
�u���s:C�C�)� �La�Iτ@�����
�dl�@!"O�Trso�0��1��m��1"O�{G�6m�`��` 35B��"O�PY���1�"usfOH"k\�T{"O^i!gc��jQ�d�S�H`�e�$"O����hF?RF�|ۂ�W+��24!�D�nzb�s ܌(<�%�P�EAb!�Ĝ��6��-G4���c\�,.!�D����K �C t
N��"�Yr!򤏨��A��خ8�x��`�[9n!�d��E��x�bNW�N�Bd���BBO!�d�&Q	M���Èr�" U�E� �!�?g`B�6��*I��W'�!-o!������KRd�)�@a!�d��	<"�z��
ss�����=D!�d�t�p��i �n@Sæ�$�!�,x;pt
c�<R�`���_�4�!��{�n���C
�5�YX]�n�"�'
R�q�/1�B�j�+Ѕ	�4A#�'�fY���
~2M�������'�R!q�Y�Y�1����,Gʘ�
�'��(�����E`� � k�	��a�'v�A�ʞ�� ���0�`I��'4����$�3%6��#������b	�')��q�:*��2C�� ��m��'2���"�.v9���5vZ\�'�4�H�V^a��G̣ry8���'��`��~°��J�hl�p�'ܘ��/[h�XsѢ�\��,z�'�� A�X3F.:saG<쀑�'U�T��O�?1Ը��ʊ)!Z�ay�'����^�R�(u gm�E�R��'�p���P85�e�㧆<@r�h���ğA-z�u#�* �0��_4n�!�䆘i�У��Q��j��F-!!���3z~�	`�&G��رK�*�!�%3��9Xv��4��CƇZ�p�!�ā?*M�i��h�8�i��o}!�S.8�	��%ޞ>�Uy�f�R!��(Vr�Տ�)j�D���ȤG>a|��|2�E"-� XbF�@�9`X��M��yg��I�pER��$h�(ڱ�y�J6z������Aи�r
��yB�\Hn:�9�k^6T�	ө���yR��chF�Tb�;�^��""��y�ꚭz�B��!n�7	P��%P�yRG�m�`u�R�_�n퐑���0?�,OT��v-S�|��Q4
I�~��XE"O����ҥ�q��a�`Ba"Oh�E�ظ	R&1 ��Q/,��"O2�x�*�/'W|Xj'H߿
8�h��"O�H��$��l�݋F'-J(X��"O�h��B�Fn�A�R�g�>�J7"O���߻(��Y�B����X����,G{��	�V��,�7 ���
4�F\!���G�F��ǝ(�D0�� �W!�䞪!��*���u@���n�8!��Xb�R�
�S �(F�c�!� ?F2���Ë
+�ʈ�$�Z��!�䟥 mj<��1Y������՟�!���_��b��;���F��9�!�D��U�}�g̗6�4`���/!�$N?�vJ�-F�7Q2Mp k�q4!�t�Vay��A3^XI%jNO�!�� �5)$ԍ"��Ԓg d��5�D"Oʥr�Ew��Q���/@>�I"Oa��]4�`P4oI$�x:�"OpX[&捜Y�U� �rz=-Yj�<�'��
L�RV���Z|5R�^!�$
Q� �j�p�-r�Jۭ&�!�d˥;��G�п[Ƕ�A���\�!�d��m��a��
!���u�w|!��}�Px�)�G|�:��I�Ux!�$��m����L.v�u(�F��!�Y�^��xs/ӗ9wZUh�eD8!���ah�K��?c�D]1��#�!�d*ipv�BV�+X�T=�$�O>o�!�W�0}��`Q;l������B�!��2�tM�Fȕ1f�L�
�#Ҿ~�!��>4:���AZ�/]�U�T�"�!��%[؞IZ���^C<��B�Q�4`!�ă�PO )xSH̫m)ҒN@�[!�K.o3��1��#q~�IB���!�?V��1�h�pY,�Qs�޿g}!�D�/\O�@��D�>a� �B�0;�!��,$N�*�b� �N�J5''3{!����}l<3E о\���Ɠ#�!򤐜<��P���G"D��Lc���#0!��ơc��#�+P1M�&�s��1b#!�d�#S@�ҀNR,=�(��KX�!�R1*	J�xj\�(8F�ɰg��j!!��ޯQ�^肤aߠy��ة�F��N4!��6'UH � ��V��Ԩ$��_!�D�M�A����+AT�1��ϛ	_�!��7:�6����N74h�Y0�C�[�!�¦W"J��&���3�%� ��(\!�W'�L�Ҷ�<�RDaF=+��0�O����D[+P`��T�A�'ݼ �"O�
�(R�u�~a��� Ɉ���"O(���*H��� ��tÔ�z�"O�(VL�7h���]�R�0��q"OJ��rI�6��+��H�0�j��"O`��.V52�p�G	y��L�U"O�`���4P�^ـ���vɤ���"O!���\;$؀��
�v�>b�"OX���{'�C3L��^*�#"OX����,�Kg��8c\v��"O0|��L��@��ۣHޟG�(�"O���I	�3Y�|q%��� �|��"O�pJrE�MP�U�E���,�"OPI��ƕ��Da���r��p�"O\��Y��Z� ����Ńs"O$�P%�M�8�2��� �4k=�T P"Ođ2"B� �fD�����g2Zt�7"OR4�qN�Sn�U�@��R�
Mi�"Op`C�W�H�`�h�K�3s�H��"Od�B&�?X�XIq��H�%�,y�"O�L�S�V�U�5�#�ôa���[�"O���Be�[E�U�B'F�+f@e�3"O�$y%��Ey7�^>JG�	2�"Oi�qÖ�{n�pCO0�T�""O�ŢR�E��4aÎܞ7�2EA�"O~4R#˘�"�����&��j 
M��"O� S�ɩXsݻ���f�X�"O��X`Ô�(D>%k�F�'�v�Y"Oj� �%�$ �(,���8�4���"O� ��i����9��*O$vz�ub5"O�1�N_�p�С8�j;]���"O� R%��)QOT~ٳu茦���"O�KЈ�.b���Č�5���"O:�sg��="���[�2�l��"O�,��)�j E�F+.c��t�"O�u������H��W٢p�"O(��A���*��ybTI�]g�U�G"O�T��
��P1B�^b��"O��4�X�D|L5�aF�
����c"O6d#��\A�E:7�3Y��г"O�[���R°�򠓯{F4��"O�t��+���3P�\�8Q"!"O���Uc�o����u�J1>�f�"�"O��H��=Y"�a#Â5q�\�3�"O|jgA�7N/�1t��*1��l#�"OrQ+`N3e�=Ih޻i+�R�"OL�����:�tAr�@VG��+�"Om��n��*Ql��FوH��9�"O����g9����$4��=��"O�i��S�L`�l�g������"�"O��PgoR�x�r��bU�@L�"Oܕ
G-�w�2	 ��^�.m�"O���] ((y0$�N��9X�"OJİ�-R�&�x���U9�>q
�"O�H	��_=R�
���"33�Z}ҡ"O�AQ�"j<���A� f��"O,IPd�r+X����,RL8�f"OjA�)'U�xtI\�f���"O��9gˏ=�]1 h]�|��D�C"O�`Q�!�
B��cfԙL��I:0"O�C�CJ���B��L�|���"OXݐp��$��!�A�v�ְ8"O�x㑪V�Z&��lV2r�>@{"O��t��uڹ�t�]�N�v0jb"OJ���J ���K�_���ya"O�Y��'
Kv�y%��=�j�с"O|����� ���J�
d�'"O��Q�f�Z��k$ ΈLM���"O�����2�	��>F���c"O�D�29nQ|d�"͕�s���8'"O��7�1��Pj�EF�H����"O�� �D��)A�DZ��\H�"OL���%�B�BH���Zl6���"O�Q�P�YV����"ɲ���3"O:�8�$S=|��ᕤG�d�� ِ"OPcti��"v�h�����-�E"OȐ %�~�@��L��\zՀD4On�O��S�g~�A�� a��+���_8���&�K�y��X!F����ɍ�]�	�F'�y�-B�f˖�k@k
�ҕ�ƒ�y"�˟|��+��Y*aE�P3�yR�Y�P��q��Cz��d%��yb��i �q8��X!xx<�T�G��yR쏷	뀵
g�6wRز��Ŷ�y�i^Zc��j!G� GB*�C��Z,�y��d�ċЉζ.�=[�����y�a�h���dE�*.^!ڱN��y�??D"4:���+x6��a2k�%�y®�� �d�Ɔpr�D�H�y"�,�bT�g�ٱh���@/��y��	�|�4��aZ��)��\��y�F�-f՜ s�D��Y��H�"�yb�A33�<��BIK#2=���yBh�n���#�*�<N?v�I���+�y�� *�Y[��#F�֕-1�T���S�? <tÃM@?v��uL�.ܺ�;�"O<l��ˊ�R�>ݨD��(D��t�"O�ը1kBn"@dcA��a�f"OB�Ӏ!@�(nj%1㋋��+�"O�Q��C�8�0���DN,{l8�,�yiyx@-��̉8��Q�U��y��9 <�#�	�6ɞ]u�۴�yr���E(M�D��c* D��*��yr'��f�����UD׎:��U�y�-[����/Nw��b�m߸�y��̖ry��X���Ro��F�L��yR�̿=!�=	�O�QG>��$F�/�y�EI�����+�Kj��4�ʗ�y¡U40�4���0�JPړ���yRkN6D%L`'O̴~�>�9���0<!���Lm�tJw�C�
���2���|~!��S�t;2k%��$R���i2��%1!�$Q%{.$Af�%jaӁ�<!��&=�J���*޹7T�hF�UP�!��	;s��(�fē@FΨ�g��:�!�d@�@���*D� �ni�C5Uk!�䓻/� �0���]����8��^����ۡG���v�ӑ�Ծ2l����d3�S�' R��'��E���cW����ȓN�Z�sh�����Hu�ˑl�:D�ȓc����&
S
r5h�e�1a[Ƞ�ȓA#,PgG�q ���`��'aN���l�:y�ࣈ�6A�F�F�@ ZH��;�.yx��G�Ly��a��Lr!Gx��)�ǀ[w�Qq3lԐ3���ٗ#S̓��=��a�`%A0,�{|ƀ1dE�N�<ـ�ϰ;�\9�!ʓ?nO ��S'�J�<IR E,@ �g'
  �E�R{�<��n��<�5���H��J3��r�<��n]�4�&	��@�BO�* ���ȓSd��p�Y�{Z�%�� &��'sў��?�5S=%z�  h6@<�+�#I��'��𙟈AF,H
z6��4��eQ�ec��"D� �ö=��p�M U�q�*=D�4�'!�A�p��*>|aSU/%D�XR(��L�n�A傍�G��u���#D� h@�[ZiN�i���~�l�as@<D��cE� <�X�xc�s,�(��%D� �Tl�	hr��B���\`�̖w�����d�ye(�@Q�m�>�)��T�!��C�\b�H���Q�r���ŜJ�!�dN�x��|ؒ ��hs�K*8�!�gs.)��ĝ0+A�q��Q�k!�^�VM��0W*ǿ<�!t�_-
[!�d�
)l02A�_��9p��7T!��onh�H�(ّ 3�T����|6�	b�'h��͟���]6'6H�D�h��E�G�'D���u�ҏKgR��/h�p�a e9D�� "�uaq
^*.��q*е0�B��s�9BEÙz���@��c�B�Ʌ iTyH6�?
Y��q�3�^C��*aI��0C$!)�=���J�3T">����h�q���e݆ZS����	Yx�Dr��:kz\[%�Y\rB�) �0D�(�P�Q�m�d0����f�P�:D��0W&ԟ]����Ͱ5ќ%j�f=D��ڔ��-:����X�_gD)��a(D�x��&T$UR��[D�2de�z��0�hO�Ӝ+5�蚧M�;o�n���	��[��D��)� ��5�F!8:����M|(!��"O�ͻa/�"t�nɀ�P_Q8iB��d=|O�|��aݑM�J���P�$O@��"O*�""��	��E!��A�"5K�"O}
�˖-;Y�P�^�#тij�"O��ɣ$�#5i�1
R�Y�V�:9���i���I$>w(�9PO��.�^%óh�gn!�$Ix����\% 6lL�h\Hm��&�S�O߶,��F�+'\a�7Nؓ)�>9i�'=��:3*Q��N�
'���4��T��'��h��+:YX����)&��Q���O�h@bdŰZx��8
���ȓ
��ϣ}t��2B�D�+��Gx��)ZF�A�4q��i�aJ�6f6-�D��t�<�t
%wS��Ib���Y�����x�$��K��9�^9r�lI1Vk��X	��|�ȓ'�p��gX�Q���؀
U4��ȓz�����ϺU�\Ȁ��u�n5���?y���4B����a�yi�̹��g�<Iq
ΘI	��AP��'Mp�ge�f�<)2���FJD`!�!#o�PS��e�<QqF[("8�г��^�s+2���e�e���D(�'.X]9��α9�왂#�7K2���ȓX2 �Xv�ءg�����^:i"�%�ȓKk��3D����:KK48v���؟��.��i6)wjYՌ x��B�	Qs�1�K�m�\Śq���)��"<a	�
�h�Q𬋿+��Db���?\��d��!��x�۱0��X@�ӹ[&���'�'R�?x�o<\�̓��u��Ysm:D�܈A�
�Y�Z�3���S.�1:D� Y���>y�\)�ȋjg)�Cg-D�rǃ� 7v�;ҭ�$NB�"GK)D��f�
=��#p.½+H>�a�E)Oʢ=��G/5�h���>P�`�XAGMu�<����<p3ᓁ(�$J 9�fQ2�hO?牯1���1�%��=Ӱ�j��y��_���:� 0	P�:�y2����lz��7{����ݏ�yb̙J�*IxSgq�,�S�KA�y���<�tBWoG>m�
U���[(�0>J>�}i6q��ѧ'��R�ݴ��x��&[C�Dk�B�B�|�%���y�U�`�4,��
q���t-Y�y�%N�b)N�#0�J�Zz��pD(Ȃ�y�E��$��&�8W�y�tA���PyRf����9'���0��u�Gg�<)���s.LTy�J$:o�TկV_�<R���(ʷ�%V(d���^̓�?�/O�ʓ��ʎaYF��c:	�hP�19���'j�}b�P�aD e@��7�
QBP�T�y��6<�����f��}�����y�+Kn;��c� �/K�؜gO��y���(���	C��0	D*���y����0�Z�Xg͎
ތ�3�J��y��ʝ(5a��vI���0����0=�҅^+@~�$`ذ ���p�U(�y;Av!(�%Lyx\�s�
�y熉%�iX R�A����Ћ�y�!@50����i��HUJd��3�yҡv{6�0��_->C<T�f��y��K��@��A���P�`���yr��f�d���O}�0���oH�y"��	J�~�J�Ämk�(�R'�;�y
� ���ЈPo,�ؠ�\(M5(5"Ote�e]� G��Y�O�5����"ON Z�����m�3/��t�J���"OP1��ܚl�I�P�$�F 2�"O�8[Fɻy�)�
�c��%�V"OJ�1d"�1\�����&��(,ؤ�E"O��uSG.�	QAH��/#<�"O�<곋ݖ~u@Ѣ��X?{��b"O��y2e�s�(�� !^.}B���!"O�jP @_#�00��� �䍓�"O�tztj{�����Q�A�4�ɢ"O����N�q�nP�N�'(2j�"O��r��.~�8��Q��1:ƈ� �"O��D���PQp�8��߰vY��!"OP��֤oY ]�p��D �L�	�'���0�#s�h�c�Z���	�'�0�j�؎kΜ�����pR�'P��tAU�:�D� �im�֬͹fў"~Γm>L;c�M!#L���=X��ȓH�Ĥȗ���q�5O_5RgR������O6�'E�Ai� 6{#�@RgK�i��Q��'�Й�Ϥ���k�� {�'�J�:Ĩ�Ct��C�[%�$�H�'�����V�L8�t�?Ԅ���'��!q1��,6R\�� �^�i�'��! ���3��}��F�
r>��'Ĝ �&,.�X��6�YYF6� �'�ў"~��O�E��8����'6h� OF�<)s#�)b�@P�QhK���rĤ\X�<�+�L�b��A�J�^�tmQ�ˋP�<�'�ې*?4�q��$m�ݢr�Yd�<I7AE�.���p�SP���b�<ɰN��&U�y��O֢[x�\�a�\�<� D��֘��J��t��N\~�'��O��?u�珊�8�1�L�Rw^L�.D�\ҍ�,M�I9DI�&h�D#*D�:�#"JjJ-�����Ip�'D�X����Y�СQu�P�BR9}�VB��v�,���h:
��@H��<'HfC�|$8�mS�	���F���Hk~C�I�_������ uR���Pb��Y�BC�4����c5g��,�"v'�C䉗4Q>9ۡF��YREe�_�bC�	�,~���k�l9����(C�I�7�6������S�h$��;�JB�&%�~���L4�x;2�̀sM�C�	�L7����Nܥ�,!��ǿ4i�C�	DdlR�H��?�L�����/
8B��%�D�1�HM%_��5��(EB�E����hÿN� @z!K±3�B�I�(k�#���KD���D!@�J1�C䉱6����VJV -e�1r�K��~B�b#��0��,Qd�pjݧ�dB�ɿl� 5
�k�# �er��(L�8B�I�y�z��qۼ��E (ّa(B�ɇ��r��[!w~�x��[(q��C�ɤ1��uB�eձ=LA�P�1m	�C䉙kM�$����;�*-���W<ZC�	����[!�f{�p�C� U�hB䉆E�`<�����t*U#$&��C䉷d�������d����B�QY��C�I ,=����=������:�C�	�>��E�I�&u?@y��]�C��4Xۀ3�*�U"�i#�잍*vC�)� Vy����\�`�,�1i⾽2�"OV�2rO��j`,��*�>[;(D��"O��)��``qɄoֵV%���D"O�����	,Ä�0��d���"Op-�P��)7OF@�F��R�1!"O�i悇,)�����Ƿ5'~w"O$����� ?�:	��JA&,D�`z�"O"mI��D'4%D��Q'��A9.��"O���2�\1Ǎk��ņ`�$�k�"Oh9) ��u��[R�1K����y2d�7�^`!CM4�`��4�y�j�&n:\����8Z�@���Ɣ�y��/-�B��냴PD��C,Q �y2��r���2}r��'M�=�y�E��{y8%�w��#lאL��&���y�d©Q��⒏gqr�����yb.��
�Di��Պ]X;f�ܛ�yBe]>��=*I��W�2��R/��y���;z��X���4'�$asc
�y"LXiQ�L�E"S rs��w�N�y�GFz�"UK�g�Uq��C��yb�ѭY�~ �1BE�c�`,*��W1�y��1E�����XL�ui��4�yBK\bԦ�5	ݔS�~DHukњ�y� �=�~����ۛG��|pD���yc^ ػ��۴1�T�ʑ��y*P,F�6�� �ё�$�f��-�y��z(T	�������c��5�yRa�(�Zmj�jє
f�Z�)G��yr˃�I�ֈ�B�{����'��y2�`��@%�m��L�w'�
�y�/��N����Z�g��8�w	@�ybE��"����֚KLH�'�W��yrƃ�s0��M��S� ��yrj�;a䆸���O24,�`����yR�1tA���ߘN�M �%�y�aH-���S H�@2y;wAG��yrF�qN4�� 	"<P�鍰�yjW+�8��׎��OR$,��@)�y�#es��a�L$�1ïК�yr�!8
dZb��B�� �,�y"jPnHh�j�#��
Q�5f�!�y�fS4Uuؐ�dm�
0Ѥ<�yR�I)a9��q1��;O�*�zF�7�y� <2�h�Xs�ɟ�F�'���yBM�2讥��(T�P -�7�yO�44O�M���Y"��1�,_��y�`��fT(�2��N>{3Vѡ�@���y���
B>���T�H��=8���y��O�5�\)��)�: UZ5�é�yB�A���uEN@��S`J
��y�卫A� ���)�<��8p#A�y�����X6H�m��1�C�)�!�$�c��=ɓ��:C��I3Q�3d�!�Ĉ�E�@{0�&��"A�/s�!�DÙX������1��u�E�ǀD�!�D��BL���*QG�p���R�Y�!�F�{ޱA�;0���+�Y�8�!��Oq��RC��}�D3u�\L}!�ռW.�d9a�=�NՑs��7}!�QI�z5K��+E��P����^!�d��I�6Hx�d
3Z�\����[�!�$K~�D�HvEI�SXB$�=I�!�ŷyP���b��*NYr�q�m��Z,!�� ���(*o�@:EbX�*-Zt+�"Op�B�B�*f���c�	8���"O�m�"V-Xؼ<��kQ$f�5Qd"O��R��G�F0PQ��	v� ��"O��4"T�5~F}z�'~ptܡa"O8��/��P~i���?4z�a"O:��c��+v�T�J�>#ܸ�"O,���lS�r�������5t����"O�1@C��O��8A4��.��1��"Or�,]*ڈ�;�kR!#���"O<8��"�T��$��kU=n��D"O
��(ŷX�d�p�����e�V"OV�2���"�(�����@��ub�"O�� 0���{�����EB��Hc
�'��ċa�E��������@�.�{�'e�H�ჿca�8xb�A�8*	�'8���
��E�P�c�L�@{n��'@�h� �N�ZL�5�A�F�}�
�'���bR�^,|´m)!7����'��{!��d/�����]�W�dD[	�'і�w��F�(�A�?R��x��'
4�Jd�̗fFpݨ�Z6D{���'s��[��ֳmM@���O�+԰Q��'��4�q�_tN�p��˒2�J�1�'V���E�B>��Jv�Ӳ-�fPk�'>,� '�%�D���d�����	�'�F��4,I v���T�ό*�~HX	�'��a#����T���$)�����'%|	��_�^���BҢY�9y�'�PH�!���b!E�?�PC�'S�	j�b��W	�`���*A*
�'��4��iÃ
��i�^?j�k	�'k��s%�FW�e�AL�Rit=��'g`���-͗w�Vh3I+5��)�'��yR��b�!���4��q�'@P, J�%H�!Z@́1;�T��'3�U�"��
��p�P�9��z
�'�QR0M��[\��:ʲ���'��%���_#Pr1��C ]����'36ܹ4FŞw�^8�%ŖɌ�3�'�d���.�b5l|�E��A���'� �w�6N�͙%K�6!�
�'^&*�A.� =�7���I� �'�2=R#�R4�5�Џ5ShX�'�*|ˢ�׹l�H����b����'�t��D4>�yp7eΆY8nٱ�'��Q��!��c��!��� �y�'j(���M'B��[���f�xE��'h��d����ӈ�]����'�~u�Ђץ<�j� �G�'A���'7@�DGܱm���3�g�%o��'�����޾S,T��S�4a ���'v���&vu�T�S䔫+k�e��'sfѺb��hq��F8!�pq
�'d��2W�*`�,�B
E!cC�1
�'��!ٗ �Rz�b��N�����'b��������Pgװ^༜ 	�'��3��9Zn�J�Ŝ#Pd���'�F�wS L��+@JKj
��'���C��p�xl`'́�F�6$:�')�XÆ�* 6 �SPI�m�b�'�JEK���ޤ�"�I�l�:��' 酊U,ɬ�s�ݍk��]h�'�"����ˁw���u��^Ό�+��� ��pe��a����"��.��d��"O�mˑF�p��Dm	�-eVqJp"O��:1`Ș`�:8h�k�('b�a�d"O���,�������ޏbK��"O�5�0A.�ye�̴?�L��"OL��j�6S���i�0����"O�Hp��]�n1�p׈��M�b"O4�� "ՒtJŧ�	W��Xa�"O�A�(�7�����%ǲ'ͮ�S"O �W.A<D�t����٣N�b� u"O��Q�J�p�s��S�f�<�3�"O��߰1����T��m�Ra*2D�8���VK���_~sȹ��.D��3���j�i��S�,<�y�>D�,�Q�,t~����f�|���&>D�H�D�0GZ�t3�(M'̔\��>D�d�6	ױU��=����{�<�*0-:D�;�gȒMa\��aP���o6D��	2F�"�AlG+gP�%��8D�$d�G v�@ 9���"����F�6D�8cC�̶|�D�)TC�>^�-��7D���՗T�:�赃��`��9��2D��s�D�Y�T o��h7��I0D���!ř�j^��Ŭ�C^����,D���Ê�
��u��(�T�"D��$D�����ޘ"�P��1���x���q��$D���O�N�� _ȵ��&D���O>\�Jp�o�
Ĭ��J#D�(����L�V�;Я��k�uPL!D� 3%�71��XQDQ�!�jr�- D�ԣ�Ĺ	��}�a����U"��>D�x�҇)S�"1Z#!N�8���� 1D�ܲ�oX.W�Ȁ�#/�� �M.D� �c`=:��i��(�>��tS� 7D���c)�/e)�G*���	4D�@��	ū~�r�I�ع=�b���1D�|ؠ�]�B�(�V���(J� ��.D��Q&��A�H	0��ds�uC�'2D��0  �g�P��7��*���խ4D��  m+7C�����7��P)1D��"@<ܐU�� H44ˆ}���2D��E(��)�p\bUeC.3TY#O;D�tB!�0A��
DĂ�X���+S�;D���w�C-\#� 	�ʂ0x������:D���˜�@"t����Vxr�F.D�B�T�_v�P����X��P�!�+D���%�\�rA�2�
��6�)D������r9�����px�-P"&D������V{��/�u�|yQ�+%D�h�����SCF�$�<`�D!�p!(D�샷��H�h�"��f�D�0ed(D���R�ʸH����#�˶\X
%�/%D�TӔ�R:'ς�
��D@:�5�%D���p,Q���ʃD�;��1 �?D�xhF+�:`�Ƞӥ<�Ȕ��G>D���o�I���jB�@_�pAѨ1D� Y�L�,М�����H\��q#0D�`6@�3Y{rl2�.�J;^��A,D� ��u�ѻF�/f�T$�6 *D���3�^6Irī�A�q�8���2D�@�"e'���������l�T�1D����ʢ(Jx!�k�:r�~�[q�0D�,YѬ�6[�VA`��(���-D����)��n��sJC�H$F�!�� } F�Va�x�B%ف-'B�(��i���ܣ��� �I,C��a�a����z�����I߬D;�KΩK�p5ba�'!��_�l��c
N�m�V�1�n�$!�=4�\���0Ϊ��k��	!�I�A�lP/��
Vf���K�	p�!�ן)��cq.ή/p~$���0~i!���,m�8����#V�c6�E�6o!�D�x"��B�94M���h'G9!�D/�J�m�% �r�!*K3!��#2;����-N� Vl�TBH*P'!򄂜x�N)��<��DҀ��,$!��<u ��o�j����4i�$(��I\x�L�w��?�~X���Yfĸ�`�<�O��'���2�IۺQ	���qC��/� Y�O���$ˊ>~p������@�%Շ:lQ�\Dx��~�J���<0���V�n�:�bQk�<��K�=b(�Q`iJ�3ҕa�&Uo���MK�����dO7f�8�p���>|{8X�IA�<���	�%f�z���#GGI�c{򹨥�	{��~�!û��0�� ����6�0>!�8}"._<A&=���"*$@.9R�d̓��?)����wMf�kDc��[ �)�dM�~�<9���7R|��/�_JAjd-�O�<)�%����db
�}��a�dLpy��)ʧ+3� ��72����H�<r�a��([�gK�$^�X����x��ȓclTXwC�!X��Ԁ��ɍkc�̈́ȓ{gB�E]�(������'�1����=H��8��- G�j5�ȓm�ě�Gq"!j�7{Ht��c+ �C I9 �M2�A�7M<���ȓ�i$�S�ab�y���3x	�9�ȓU2�"�� 1��pFӷ���ȓe7�,�B$�%n�4dO0.>L��ɷ`��I=QIF�YW�H�B���D�=��B�	*d,�'�|���2N��B��B�I	�B��0 n�eF�(��\a��*D����F�"�J��5�}��DR4�g�G{��i-���C�y��|���!/!�� ��c�O�]YT���6"�O���$Ǯ.�8E3T��/����WF�+�!��8�v}*v+�d����(#!�D�7h$(��r�'4Ll���tW!�הj����D}&��c7�
_D!�CU�L'�	�(�Z��֧Y*!�d�	�r�BҬ�`|��Ͼ�!�d�;h�Ԉ���11���4D*�!�$[92}�:�n�-1���"���!�$À�ʼ��T#|��Q�@�l!�d�����4˚ykPt�vB��w!��Oz��X�3/,>a���� �Js!�DUBѨ���91i�mڷl�f�!�M��;cʁ$��$aӭ�!�䙐j��sFc
�%�h@��&�\����)��)A�hߙ&�|4򠃐���s�+D�@�A�Ah� �q�ˣ:�@��L,D�l�ԥ�� ��ib���!h��p���&�OpO�L���g|���b�ՠg�Q�"O��
� +��qd��v�ԓR�I)�a��FI$1�� ��#�����j��y"ňT����פ�)U��y�n޹�y��8x(��#��N�`������yBf_9b���`FX�Me��%+�3�y
� 8�P�8���%���<����"O�������G"�#�lD��� �d"Ox�S$�FpZb�7F��Q�V��e"O��C㚬`"�Rdj�<LҘj�"O8�!�
LKlC���8�Ҍ��"O�a���W�P��h��dG�2�B٪W"O�e��֋n���f&{�|aӐ"O��§nU�0}�����5���jE"O��p� �o���� H��rB"O��T�T 
V�{@����2v"O)3A� 	G֪�
���L=!�"Oh1
ԍM #)�11�E�+�:��"O1�Q��#�@�:Ѓޯ��	'"O�˧�׿�Tmx�ɲ{��!Q"OT�Q����N���H��g���"OlT��eD�T ��7E��ڠ"OX��C���ߙP���H�"O�	t�QH�ԌZ�,2.lq�f"Ot�qP㛥[�~up�%Y�fz��"O�]"a'�|yXP�F6N�"x�0"Or�sS-�����v�#����"OI`���@"�n�}��b"O�]�Ǻ7*D�F�YL4�m%D�0 C3"~^UbQ�7g��=���7D�db��<q�aT;v�m�B0D��ɏ:L�,ڔRἑbU,+D�L��� B<@I(H�#eV����*D�<b����7���a�F*}�t���>D�"�����`�4�W R'� �6D*D����Jގp T �@�%ib���J(D�؂�+8
�&״{�hhC�<D��AcG^%.���)��S�|�<lȑF:D�Hq m�v�z`��4yd X��5D���ŏ$B���)���V�/D�p@s��o�+���1���*�Q�y�gH�a�Ġ��q��%)��$�y�Évv�5��C�g�Q �R��yBEK��9��OH;^��#N/�yR��9:
��!QB�B�`D���M$�y2�	;c�u'9Mx�:��yb.N�w\�� g�B��Y�!
��yb�B5k�P��$#��$�a�+�ya�f|�\Q���*$�(�!,�yB͗�T����#���?"h�Q����y��ژH�2	҃SFk�X��cſ�y��P� �vE�?)���[g�_��yB	ӟRK��cf�:!�h��y2��>(d�h2fJ�&X�꓆(�y��p�"3쓛V����:�y���jR����R�`CPpK`����yr*,p��CE�*�5k`�y�=i{Pa��'��6��هg*�y��ԍ/y� �MJ�+�j�d�V��yb��yv�Q�'�=��91Tl���yr�=��8怅rL�+.�1�yBΚ�}��e�U��z��Q�@��y�₥�h�dj_�tOU����yR(�(aC�!��lgT���>�y	�*����]�Z���"	�-�yRf�{���֯O8D�Ɲ���y���<7V]�Ո�1A�1ڶ�0�y�aåD�и��g��6�|Q`��	�y�/I��h[2��2s���I��y��ʇ)�x���l_�)ώ�8 ծ�y
� ��i6A��:����*7��K�"OԜ��� t��Xf���� [�"O����P�B��,����)k"HI"O]7@��T`�)�'�ImS��D"OR�� \��!���z���"OL9��
� $X<��G[	7�d���"O6����T@l]���^�y{B"OHU@�K�*�:��稖>hɦ,��"Of��JԡC������a���"O(aj"��W��0;�2U,5�"O1����<x(����8Lh�"Ou����Ot���C//����"Oơ�P�� �����;���S"O��`��!,� 1S� =�:�ɥ"Of�`�o#�x�%A/N�n���"Of�`���t
���W+"�t��"O��ї�^�F�$!���\oQ�X��"O6]�eS�t|���_@Cf<�"O(����ФV��Zu�Di�`�a"O��*��G�u�����	64l	D"O�lA��^;���!�l��Mk�8
0"OT}�s˔�QS�yр�Ԅn(��T�|��	3!����VkF��T�$iND�B�*s Z$æa��K7����g�P"=��	��6����C��?G B��ȓ)ݑ�S�<K'��.u�(�qش�Px��E�+-t附�|t��(�E���yB��S�V�����z���������y"���|}!:MXp���2�Y5�yĎ�Q<`�34m�/kw�q��!��y�Ɔ5o(�K��.*�Ѱ6�C��y��a�:(�j�'���@f��y��V Q�8}� m�0"T��Jf�>�M+'
?�OH�P$�,��$� �L�J,{6�'i1O����$<WN!��D��Q��!w"O�ɣ��
�F욠�Փj�����|B�'�����#<��u����D��X�˓�(O���QK�s� Iɥ�)M|L���T8� ��D�9m�Z�Q5O@j���b/D��`��&�Bv�а�^9x�.D���摆�P������*�A����O�C�ɘ;9�� ઑ9��CuA���"B�$%�a�� 3���2	żq��|�'�:H�棎+"ŪȓB��j�@���'S �T��/AFt'�>3㚬�'��a�E�r�^e)�lT%\��*�'[��׭W��-�S��X%����'�&5iZ7R�AS(�J���P�'&m�@gHM��ĮB{��	�'i��9Х�9���u��n�@�H)O��=E�gŸC-v1�w�#���J�O���y"��J��y�/_�DKШ�� �yr�5l1x<8 ��8�|�;F�E��Pxb�iT(e�O#.��Po�"H��|���� �DYJ'CK�TT `,ݢF�m��IS�'�|�����8��5����?*�^����:�S���H�C:�q���V�Є���P!�yR�׿{���d�e�p��X��y2��:IyD�a�� N�Fl�����yr�,[TȣA�{�	�TΎ1�y�įV��l�P��y|&u���&�yR��-)۪遄�ʩb�t��3���y���������dL����sdS�y��ɫ:G�!��m�YL��gC����hO��� ��i���>�l�u�C�9���"OV	����A�F-�f@:I� �)"O4�#P�J"G��H�%UN�!�"O��[��[�zl�2�� �&=�"O����
���r�l� ��""OJ�u&I���bw�T�2��,I�"O~�k�V���"���@�*t*֞|��)�
 ~ѥ�N�Y��r7��$��C��09f�E����W2��` I1��C�I�[�-3pGƨ)ɪi�ѬT0+�z�0me���Iz�t	���v	��вG�D�DP��<	�x����7���:,����+&�Ȇ���Z�͘>��j��ZK�j��<�e�)� VG�S�S�fd^钤��&M6c�\G{��$&E�`�Ћ�ƝK+��Ch����'?�i��	*�D)�͘:y�`������#}�B䉍I�}����u�L�k�r- 6�2�dx��k�+Ր�������'���e�"D���QoZ36 (��m��7~���g�`�'ў�'6��44N� �
�
����G�ഄmy��9��K!i
���L�@5�gjO��hO?�䙶A�D��@Dه�0�9�n��t�y�ቛ	%��qA�^��@1�tL�&ȶB��h1D�:%(�#u:%��G�+3�~��(O�	���d�H0U�d��!����M�.X�x�>1�Ot}�)����Bc� 0��i���d1�S�	V�3�H9R� M���B���i�!�dV�4)!S@ׁQ����2��1�!�d�Y��е�&/�4��diG'>�!�d�4(�D���홆�!���wЮذ��܃Ij¹�b�M'�!�$��',��!A��ze,sr@O2
�!���n��p��/C�|9!%� Lt!�d�\ҨmiU��0@"y�tF٥wp!�Ę�2 �k )
�
߂��'8!�$X�`�(K+��	��Mz�qO��=iI<1a�U�X�X@�7�U�.��`���q�<�`�Ҭ$P��6��"A�Y��\r�<����"-rP*0��!&2"$����n~��'m�I�0�NxȰ��I_(9�11�'�p)��&`�tq(u'�&k�^!�'#4���F�+XW���� _�<��'����VύF���3a)&�
�'��� 1J�=#��=q���
���
�'�>`������b�A ��3�'������L�4H�w@�"��8
�'%F(Z���>�
���Gݖ-����'���Dy��I�-"@���c��M�p���H�k\!�ՂI�fi���L�O��U�#��Z��T��H�N�ˠ	� U��T�0;�a#�"O�J�*�;*8�3/#ĬL���xb�'ОX�B27��5�agT�)>��(�'��q�H�/Y�X�ʊLa��K�'S
�"c�sqX�4���9��@�M�H���)�Sy�6(��g^&�I+�'M1V�C�ɑw[�(���"p[�T�0[�v#=q��T?)��Np.PB��F1���B�n D�hʗo$%}]�dI&}wVL��g"D�
"�,��]�&�,��f�B�I]t��BΊ������2B�	�o-���O�#����1/���	m�Id��x�C�8E:\Hփ+U�4�S�A0�	J�'ډOg$��gÓ<X����I�f�9�!�d�OT��I؆	��AR�/U�1������Q�d�=1�y
� �����B�铒��dU���t"OZ��v���I�0@�Ɠ�VT|�	��??���iZ�c�04��o��?�h=;���u�!�L:	�\,�U#B�>9PM*$d��ax�	Ԇm�eE�8dT�uB61����$5� ����aO�YƄ��̙��|��hOQ>���e�7V�J��% �2=�r�(�:�d �S�'taP����J�%u�]Rb�[+�\�<Q�&к����\Jn���*�[B���ȓoC����g:Y��GƄa th�������j0s�y"Ҏ̼#?��6i;�!��1I�ZG�uB<Gxr�)R5���zMx�c�J�}��I)�d�<�U��`��I�#L���99v,�a�<!�T	��dAq{�J�萉w�<	� ��u�d(qE��@�83��s�'$�?I ��D�ʩ��,�0�0X236D��c���z�<�A�^�nֽ;'G���*�)�'�9��dM�B,)�˲bA�ȓ!�^��amH��J3�)^�W��m�ȓ���� �[���
�٣�Ή��8/�@��C(R>��B ,�5�@�����2'ѫ'^��0o�~cD����
PujZ�7{�yr��\���ȓ,��ݪ�&�B�����
O�,�ȓg��,��B��c�YS��m)�a��x����F�o��(�eG)���ȓ2��#��؋5>(�Z6��I=�y�ȓeo�L�#E��+��\3bu��8"O$k�"ɳi5��f�8,�D��$"O� ����m�b�*����9s"On�1e��2wj5xR	�"w��%"O���a��d�]a��Cu���"O>u���>I�`���N�<^
�r"O���`HBu�\���R�A�e@"O��9���@�Ĺ�r,<����"O�ؠ�H�@vjlJP	];FX�1v"O�Hţ�.*g�Q��� �+��~�<iéF*���$��!L"� �-�y�<��	ܿm���`LLgB�E��,�|�<*��2�k����2� 1f�z�<��k�P\�Y0�*���b��]�<A�AW[�,�@f@;`�Xu��.�^�<�E"� ���@/�2�;d�Y�<�XX-���V�a*�K"N3|o!���Ub M�'dd���c��&�!��O�VȠ�h���.p�Ij�"�M�!�=:��H�U�^if��1�+��p�!򤄔w2��;}Cb勃��:W�!�$�S"e·�]v	�ҏN�b�!�ÞsZH�4e�eK���'d<!���-(� ��n�j��8!�������Jj*�2���!�đ"�5i5���#L(�b��s!�DG	��e���[T�p��=�!�ĝ$>���toT�~R	s��
�!�d�,��kB03�~�s$T�;n�x"�/�Ґ��/P�W~���6��9~gnuK&Η������ڑ ��a��q�l;�ņ�u�޴Y3�^�I�dt�ȓ辡C��c=���qe_�5��ȓl\��E ��fPc�$[���u�ȓc�����N�Lޔ��&e���X��s.D#7j͟i��0�Ñ��B���4/jш��:�4H(逭:��D��S�? �% ��N8��A!����K�"O�\�0���r��ݠ��<���@�"O�d�'��,��}��V�:�|, q"O��S�hJ`������#̐�b"O^%�2���'ip��W˃�{Є�J`"O�d�b�%&y�Sej[�að$��"O�,*�4z���c@�B�h�"Oe��JR,k�6���K�(�p��"O�	��'Z?t \�T�VU���C�"O�X����� �|��m[a"ON��E�
"6�=*�e��Y�xÑ"O(��tbT�Cz���w.A�����"O��ӅnL�@v8�z#�Sh�$��"O�<� �/9���Q�Q�z@�L�"O�=��g�	p�6�$`�-0�蔳"O�MӅ� K"	�����#�"OhP5N�r�uZ�M�kF��5"O�(��B�I�&P	��٠PL8h@�"O�
�מ=�I�k@50 �E"O2E1�'�(	�����L**=z1"O&�yV�(o?b��#I�?.ve�"O�Eap�PU�l��ai���)�"O��ó � r�ޭ��I��d��,�"Ob���C)0��0�Ƙ"7�]""OV��R��9?%&1q��_ ߎ�@"O�1��Q�N���Y�č��"OH���&���%���Ҁ;�"O
�f$�7���YOΣt���P"O�����	M̭��Oӧ#(���Q"O<0���ٴv ��x��Ѩ9��"O����#C ���6��!��]`�"O�]�F�[N�=b���tm��"O�D8ċS?Q�HֆqkD�D�Bf�<�1@�v�l@���	7�CFO�b�<�c��]�l�(KG�[W��BP)X]�<�eC�I�����BH�c��`�<	�%D2*��5J��V�r
ӃAF�<�S+OV)|!Qg%��<\��'�Je�<!�@�<gD8� {*Z�d�g�<�4A܉���Nji
9Z ��y�<	�*1�F!R1[F�D���!�_�<� EM�_��J��Qsn4��n�<����7]L� ��B�`���3��d�<�q����.Hۥ�%�����]e�<�p$H�"����B�Y�-is��}�<�r�؋#��%
M�nQ�p1�#`�<���Z�jRz��B@�3zTP�2"�{�<�3��Y�� �&�*��hBt.t�<acoߏT����B�=%��,�I�<���� �W��4&��1�	F�<��Y�'l�۷i����q��Sj�<��n�tI��P�8Y�ywH�g�<�2c��I��\���
:Z� �\�<i��[P M�Æ)	� ч@^�<9�ʍ4dO>�#B��Y�Yj���X�<����ؒ�g��>�\�C��R�<!�耇Wz*�HA�y`=S� �M�<�ѥڟO[ep�'	+�,Q�N�J�<���H�z�0L�\|��(#�^�<Q�`�<4#�U��J�I�l[�<��<԰Q�Ǡ ��)��^o�<��N�
�l�Ԭ}DҨ�фf�<�5��WUެ97��c�0��ܔ�y�&H/}�P�T� *�N��"�Z��y
� �J�%J���\#�$,B2��"O���h��"r<����*jA���'BH�Ӡ�d�D�V�'"1p��D0��Y�����	����Ϳ#� 8h�&#*PB��'��$�� I�M�ɧ(��9�N@%^�\���9w~t��A�'����g��c�	�	**�HH(ڵI�FX����R�J0������7�f�`�%0Fx�ɔ:#U
�Ї�-�@Qq.����?,P���v�~ZQ��W�\�c�OO�k�j�֥E�
k� ����O��,��(ƑkXR��@��{∏7{"����۫q>��!Ԫ!}Rm�T�r��C(ՂpHT,�1&�V�Z|s5�?9�W�EZ��5�4�R*GA�583��xrg�^�zlÒ�X��D���II!+
z�rd��4*ْ���)9��� �.B�~\��-�N��hP��bE
9Y�8�&?�~�3��')XԙGH5r�O\�`�ߜ ��2"��//����e
@7	���!�L*%^�Ԓ��
:Y��� f��Op@�w`�b��:���coY����)�ƺ#��4��>�O��4`r�M��B*͞D�ᡐn�2Jx�ȉEh�$�����|$��I"��VlX�H�^��E��cFX�	rP�xk��֌#F�!��Iv��	#&��6k|�X�X�Q�_�=�L�`��.
PD��t�S�p?��Y�~/�8�W��|.�١��!{��~]����Z-;�g��9��E �~�8��?/�����+l50p��UU�'��ї%��<^��C��ByB��<H�D ��F��p���튨16�ѣ���3Kl�عpG�/Sݪ�
sZ<I����]�k�4�3B'X�B�(d�৞�wbH��"p��yt�C�{K_��~"�i�� Jg��V�3"ʹKĵzs��3`�J�a�=~xrEԃ�O�4#6(c$��ŉ&?�d���|�i%�ۨO�R�	f���K0')�Lu���ēk6�p&n�?uʌR����y�e͕y�Аd@ �xt���I��0?�t�O�*d���R4RI�m!�iВ%3�Ƀ!!(*˓@O��8�O��w8��?Ɇ-�yvP�F]�t���2��S�'ۺ�RV��O�"��'ޖx�֋Y�+��� ��(�䉅
C�@���H��+T�6-�P�bH�9�tj��}�h����I+����_�\��ʲ�&�0���d$�2S� H)P$A�7��9����yr&Kw�:�E<���p����Đ0-"���U�E�#���Ӻ�"�Y�T�**O�q�'�H��}��=!��5�'�v�j�ş�:`Uy��޲%O*��s���ht�%�S��\����z���kt�I-jdL[����?��mP3 �y~�#?� #Z�d���'���框�p�]�f���t��!�%��c���8 �U����d��%L,�rЁ�jt}�t�4��T�$�K����Od�T(�D�z,�@c�W4�0+�'"<��G��b`�E#� ȤJ<��O�f��ɸ���IX�^�,|ly�B��BbD�Ñ"Oֈ��/T:sG��H�_"o΄��"O��� �*|����W�,Q@���"O�y�"�nvbq�ҏPw���qF"O^p��JՕ*�aJA��+Ap�sS�ɛS-<�q��
U�OV��˳M�9o.�zC���م�-�L<)� ��>��c��@��-�r�� j��� |���O��@�+�.�
���7CU��:"O&A�֯P,�>�9�ԱreT={B8O͚`Sp�Fwf5<Oh�@-�:J�@hy����Wj@�R��'����B0*>U��N�1U])2U �-k�f� �JS�H��ի�ڈ�j�=��"�	Q�Z��׍�x≥�Ё5ZtEVe%>��;�8%��Q�2�����х
�$хȓ����D��w�H($��Gؘ`h�/K�H8& �,�����?//:����1�s�����>T�p��P�|��I0$<Or���P�~��Q OD��M�&�TRf���g�%Yo0݊�KK�<15&~j8h�U擬��<Y��A:��e���ۧX�`�a�Or�ɷN���vc�f.0-P��_q��3�Q)A;^��ٌQ��*$K]�^``(�O�=s�h�4L�J'q2 W#�D'���6�$�?q"��㦡��ۦU���M����̼�e�Q+ �ېm��^�\���K(<9���3�2�D��Ek(��䊝-Q�-#�OӒNY�B�R�M���I�}��`���6�hdr��(�~B�)G��8R���}�5�\��p<Iӈ�UsL0�Vŗ�vz���E��I���a�	��(k�OҩsԢ�;rLExE�+|�J��FE��P�ɧ�ӭ!_i���3Q[��G�^��f��X��G#-��Y��J n8�i��t��I�L))�L_�7 .���$����r�R4PO,�O)E��OEc��b�Б$
�g Z K�P7@��Y��KkC�lZVb2 �1���O��x�E�08\D��!܇Y���x�i�����F�54���	��� �<K����f��( !�ɑ=]���2Iϱ!0,�LL *���e*�	�L�̑���Kx2��5a�lȑaOو;�Z�Z�#���0<yU�΍x�R��7�W���"�cZ�[ٶ��G�Į��P�ǂ�d�ȳ�{b��3E �����O��`�Ӭǿ;6񻣫��t���Ot`�'�W�2;d�R�c�Iy��؇A'��
���*�K�5G��|�ьǷ/�v�@�*ϯW��Q�O��D��OV�J4�A.|f�4�T�.r� ���B_̊��2[@yȂ�׍&r1�B�Ol�`M���Ĝ�`X%Q�iNШi���#:�����i�ԤM5zT�Ã�˃[�T=q��ݯ�L�ǅ�9��U�����=Q��IV�r���@�O\%[�WB�,�rOH7�Lm"#�'5���ȿ%Gȴz5i�U����K�,?�0����?I� @q��C  �E�و�Z��bD8f�4A���TP�9a�>�6��61����S)_\Ƒ�=§Yؚ-(���e4t0�i]�'�TX���Y�c���"~Γ-�4�B��$�V������tܸaڠ�.��Ha�K�O�dj��/�<�b��|Γl���]�VJ&���L
<d�ԏL�*d!�1�|�%NL�%�"�a��O:$Y �	��K?�wa�#}��>+N�;�ǉ�
r1O^=�rB�y{�\����h����'z�T��G�
j���ŕ�a9�CѮSV���Y8r���r��a��Lw��zx����܃g�1(Ӆ���m�40�	�B�0x�5���.������E��K�Y�q�W�=7�YJ�LG�.~�Q��`�Gh<y��%D<�Ȑ��3*K�,3���0w?B]JԓxBN��d�d��D�F2�O�������2�")R�F�f!�:wȩ)ъ�6e����J��n`,��]���Ek��<E��'�  ��K[ Y�RU�`�Ђ|��'!�U��i�$ko�(
�
үx�0��'�lT�6Ə�6�4��'���r�!�J�b��L���z��a>�UHvC�|�|�cc,��C���R�����ȪO�B㉊b�.F1���MI�ȸqxG�>���k!l�c�h A��%��^�$Q*��8�6�С�y��q���ŮΆ�)6ʍ�b�9yAgK
P�2I�"~�	,x�H5R�ڋU�<ж&H�W�JC��!S
I[�H�R<��a�#e�4�G������p=!2哯�4|�2� 3��WE�cP!�܁��l��ǊH	�4:@oZ?!��(kd`��E"&G���FnO�!�@�B�	JŁiu���C�έq!�D�7+,`	CD��k����2�!��+3�B��� T�F�8���	!�$��(�z��VK
M����Ӡe�!�Ē�lB���p��".��	Ö��'4�!�;bAb�A&�@��2�9�C�+<�!��4Sm8�QE�=q(2d� 5C!�D��%!���c�[lTI k��7!���� ��&B���o����	�'� i�`3z+��uhN�t��=y	�'D�1��i8O7����aA�>1���'�|HqUB�=rr�`�
X���*
�'-H|�6"YkYX��P&� );��
�'�I�s�A�]Ю=y�IƧ&�$=J�'�4�SL!H���ዟ.U���'q��#� Ccv�J�DO�xQ��'_~Uhv`�$Xm"�:P@�O�t��'@`��T<ʩ�����y�	�'p�TÓKE���M�7h�/p$��	�'*�����&@��+�dI�}hܥI	�'�2�Y��71V%�a+Fr��p��'t�	r�gKB���*l�R�h�'��#���@�V�rk~= �'�έ���4;�X	��Ʋh�,͡�'�؍��
�Q`@���
+k�H�'�Bĉ$�7/�.���_${�����'�J��AȌ�Y|z}�R)��
�'eT����h�̑�ШZ8-��x��'��x�塟�n�t���FH�.���	�'�8��L��c}��p�D� n�
��� d	���O
����"2�8�"O2Qx2m�~��L�G`�:#��H�"O���J�XwLp��OB�(xF"OL�2ѣ�ILHAr���:�
���"O Գ ��!�����-!w8��$"O��i_�jD:�GP�1\ʹ`����y���&м���}^��Al�
�y"�C|L��>#������ybo 6�DĢ̼9�a���yr*C��\������ �I�
�y�k�}�\l a�ώj��P�AlO��y�D��,��D�]�*O���1C׶�y� �D�"�2�'
_¾��P�ڒ�yr���uft�M�����GM�7�y�
Z�cj@�T톋+@�E��.��y�h�/��X��%ǃ9�J���y�gH�f~��wĀ.���`�ٰ�yb�**n]��d�ܫ&����yr�~�K�3�:�8�hǬ�y��&�z�v���Fz���F�"�y�0+QnXу@N�zŌU�*��y2B�:�����B(&�� Z�y���#�Ҹ�7,Z�E1:x ����yB�تR�f�����(==���Gf]��y2o�|�b� ���)87�J<�yB�U�uY"$�JҔz��p�ӂ�yra�4��S��E�t�x`���X��y"�����9���j�.��m��y�!�pTh ��kR<|#Zm��N��y"�*L�����#�VP�b���y2���+D�|������|�"�U�y�Ξ.��x�ˉ+�8��1�\"�y�!Gǈ���%��~��9��͋J�<��$�qx4��k�5d�pE�$�e�<��ғ^�D��L8�8�HviH�<!Vʆ�'�n�a�m�\�fm��$K�<��&�*���3�����O�]�<���F,I�IXP��m. [��F�<�s��H�4٘� |֐�FCj�<�0 �#PzN�a�Xf�9��k�a�<��'H�@�H�2G�?��qئB䉭En��fG�q7���G��G̺B�IU%;��r����?i~�C�	�,[�,�i��LA�C�6qܔC��[��YV���t�z��ќ|\BC�I���3bX S���p`��z C�I�r.��QE�u~M���0�C�Ii��bEU�
�Z�Bso�&��C�I�F����_,@�Q�2���C䉇5p�8p.ťn* D��c̫M��C䉣9n�@����N�H�Qt	�yOlC���|C�ĝ�!BxyA��8'&jB�ɳm�j����'�^�ʴV�HB�ɚXtM��NA�|ę1
��XB�I�xp��"ԋ)���4�f�C�	1tp�q��:���t* rGC��"ɂ�y69:vIk6��.ZW�B�	j6��@ю��$F�,��:զB�	Y=	�l�\G<m9gʃ�P �B�I�m U�V�C"�&a�t�e�B�Ʌ:{���(�;2�H|0��m)�B�	<S\��x���.P�R��aj���B�I�)
f$�ЪФ�Ϭ�x0	&D�H°�ѱ<��`�	ɒ0v�1��`%D�� ��p$!�lq�Ã̮/��$�4"OxM�q�)���Z���}]��A�"O�(Cs인}xȶ  D�D�&"O|�э_�G0�W	B�}�����"O~}s��)QI�5S�bP�S�j�J""O�9�&n��|Q�� �«��p �'��B�@ܓePDQ�z�p��������Q�ȓe{>9�K�p�F�8�nZ�D��'���3!CȺh ɧ(�  s�� � �6�"+ڸ�b�'A I*�-Dx�I�4� �U�B�7�N�s ��PF�a�g#�Zt(�j󭄡9 ,�;5D=Fx�a����e	� ���@���I� (���i�~�`ET�P� ��h��.�$&�=X�ma�"T�v���n�Cg*P���m�AG�
n�JH	��I椡Z�1}ђ=�Qc���#.<�X3홈+�1A��4V'l�A�����
�H�|Պw����x얎E�T�j�cYp���y'�<|JXC1ĩ`>�%QgI�p�D��ǄdYȆbT0φ�?�*֫�JV�B�m��]٤��i� ��d�11]3U�'��ɹ^=B�JM&gP� 2��ѭN�2��`� 1��p"�!&b���~B��3�I^�������3��@��,D��\b<e��"��Z�"ҧ��C�Z�>�b��B��Y��'Sk��1���-:�R,{�L�;w*�V����=yG�3i
�"$�S�^`��O.t�h�#PH�C!I�8��9����Re=�l��c��C�b�;G9��!�� 3��l��'��T"��U,�,l5:�[d����&#)�<\��8'Dh&���b�J�St�?q�A�o�BM�g؄S@������O�(����)
�"��Ș���F�FD�,���k�"�rR��+���Q��;��]��ς�$�r�IϞGF���^���'Ƅ�e[& �g*<z,Jၚ'Y�} @�~�xՃ炴��l����z.B��2�!d� �f�@eʹ[����Q`��'k"  ��$�a|2�%/ Ȉ0B�g�d 
&�K]b�d�1�	�#P2BX��Ӄ�fDq�\�}<%;��wi�?�\!2��;Z�u�"LBR��`9VaH?LOܼ��3&g��1d�E��
�`�撊|�	�Zlz��I(џ��ċ� �D����s�"��3�_G�P���
4X�a�t!1"EL�/m�`�GЏX8�m�������,�O��ɣ%U���R��E�]c6�s�<O�AbeoM,P�PD�-O�<;��T�6�Z=cI~2�`�F��SW�:t8ȌI�i[e�<9A��?�� �@��-^�a��n}�	V�xE�"�4�i�m0�
V�,��$�'�tؐi�)���Bbɂ (O����6�$��1��Gn�X�Γ6
S��y2� k��y�O�L�s$E��%�����/'p�B�1UX���ĕ`ۑ�<��C��`���J������"���ÊT�"���(<�O�̓�K_5� �2�(���I/|)��Zt�|̧@���&	yd1�чA�y�J��VE<ȱ�哿 G�@"2�F�r��'@���d$\M�S�O�(@�1���������+	���	�'�viy4J��Jt,�CǮH.W^���'x�{U�c��Eb�kɥb��p�'V ��A	��M�S��5��Tj�'h�蒄[1lU�TGD�$���!��d�15�|Y�8ʧ{�*T��@
�1&rq�Ajx�ȓ6�~)��')߀�[�˅�n�j� �e��M�z���O��Ct/�[ ��NI0x�T"O<�%�.�Fd��-LN?�YJv:O �
��i��L�ԣ?<O�=q0'аc�����
&E:����'�\(ira��S͎ �˟�_TA�c.�27F ,b�O�}���d��0�L��e�7I<��#n��Ay��Gh�5mЩ"�Jt�'3[Dy��U�2����7l�;9_Z���xt�h�l͜A��Y�q*[�S��ِ��Ȃ��G��M�)O?�# ��s#!\"�HKF*(T�B䉪&X��X�ORp�q�ӒY���I'�����`6%��I�#?�irU�ԾR|R��ы�<7Ƥ���V�]|�a�eϓ�t`��b�Q) ��2f�u*'4��[Q��#*R�D�Pᒍ/��h��@(m�	�B�(DR�\����	����ٹ9B�)�o��yRm��kf�Sj��#LLQ�F�;�Ě6&�G���0J���
������~RaұHP\����	�H0�0�0�yL��,���rӽ6M�d6��D͕z��%��I�>!�-"扙E�)�� �1���>V�d�X��ݞ��+"O��!倒T��%�E�r}�EH\�U 0aE�/}b�0�g}�d[M@��@�^l�$�{E���yR+N�@	�PzeI�b��-���5�MR�O�� yL2|Ox (��?�X��L��e���K��'Д�AuQ;y������2��EiS��T�zU)�2u|C�ɰjH����3�8y�$�vb� S�B� Ͼ=����9zA�=���
�i�L�2$��R�2B䉎)�H��l�%A�:�9G-�U����իoǌP�Of�G��O�����L�cw@`��&~t!�"O�5[�G8|�vi;�I�Uh�8��i	��A'�W,i�<��5G6<��+�J4��TH�5U�|����R�Ջƪ��?���[$}�ݚ�X�"���S��R�<���S \��A3�ÁB
�3��H��4t2A�O'������ �x�������BB���%"O�@��N+������j1�	�0N 	c<��{��9ODy#��HEM:Q��ò [NA#0�I�x���`G��b�O�a0�mF�p�%�@Y,4�a�'a&����˦}�̔�Ơ�&i`��F��i�x�wJ�9��)���P���3悁�4�YIwB(�g�=D��@esRtᲇUS��)�!�g��(�ᅖ-|V	u,�Bx���s�΄z&���׏բz��e*�N'�O�Svo�#q0��	6�\9*���0���h�H��E'��C�	(C4<ñ�(M�0x�3�G�:&#<Yg@& \�X&�G>��O�Q[Ӫ�$8o���Ӣ��gJ�r�'����fTqD��(S� ��a���>�:���JЗDQ��S��y��̔]28��E�&��]�����yb��(�Jْ���5[�Ո�y��(t���,�2W+�yr!Y8>}xAk����| ���L��0>���Jl>e��g��$������uؖ`R�1.�-b�'��3�=Z���P䗖0k����Dʹ3{ P�y�8�?-�V@�>8����!�8�x��F�,D��B!�Z�	0���Q&1�AM�)��XpE��ҧ��a4 ��ԏOi���tEK��yB�� <+\���</��3dN?����	V�i��?\Oz\���E�U2��`f�;&�{"O���"��/�*��U��s��Lc�"O �r �<�`�JR��_�V!�"O!��ʙ:��غ��T:b(�eH�"Op���JtD�3ퟢ�؂�"O�|QH[�/]�)��L�W,h$"O&i)�B��#~f�������"O&��󀅑Q�l=�� ��V��c"O�x��]� �(s4/���(Yp"O\�[`�Q�>�z��2�Թn���"O8�C�M])l��`e#�Wڦ�YU"O�� ���
WGl4crZ=g�:�@q"O6��b���W%(]!��D�t�0��"O&��0�S|�h��Z�qӳ�^�<�S$u �``�̚7$X�2r�_q�<��LC��|� {~�p�`�<q�D�3Z�e�WN��� ,LD�<Q`o�� �n��c��4m¼1��L�<	��B!s�^!C�^>^HD�P��v�<��Ā$$�U_^�Q*S'Z�ȓ �.�"�#P�6p�	�K��q�ȓ^��]ɵ��+pA�		��^^�Ʌȓ*д�x2��/j:J��L�:u���ku"�c���(�ܜ0W.�ne�݇�J�ce�ۘC�^	5h՟s�9��#�M8f�A&�z�2���(� ���
Rf�!v���j\:6�A�F��I�ȓ/kZ<p��1s�B5:v�E�M�ȓaG4l8�
�#Ol��񀎓�u��S�? v	9c��q����Q~�����'��=����Cf�mkd��ZMФJs�]�7�,F@I�w2~���'Z�<��FJ�06d�I���29��c��Q�<��CP���q�Å�R����҈�T�<�"K�a|P�X6��VĄ����F�<��jG$�@u���͐s���@�<A��[�wS�A� "�yI�M�@�<�RÐU��QvDJj�4Y�viGa�<9ǆ�˄�C��#E@�`��B�"��ʧqhp��S��{����@�cVұ0バ�?�gJ�-��f�
1: ��~jO?���f��1BrL
$L�
�84A�:n����7O�P�$.��Aꧽ(���"�A(�5Bs͑��A���>aq,�i��m(ЎZ$��%�'+6��M�|�M@�"�8Ǹ�͓�-��'�+j��,O?m	g*�a�V�P�^�ZU���8n��UC�1l/�BQk�>Qç�"�1ffI9YxReҩ��tIA��ab��s�'�F� $'+�ST⓺+����L#q�!E�^w�`���-�џPRG�S`�Q׊6��pS���2J�U���I��ၤ�iӔ�z�É�(�V-�B��9>�Tםk�O����7��hi��@I2s��b��Ϗ,���N�S�4o�Y(a�DG2,���j'��O��|(���8p|0��߫t&6�m��~�Q�Y��
J2,�u�<pf!�XApа�dC�S3�4�谅��b;��[��ݹ%8��1�d��c���q��f���}��W�����Ot�J���ǿg�X��'�v�Xs��Sbf<�q$.�N��ҁ �>4���"s%��<�{�'~������-A��e9$J�$�,J�'ƥ2ѮJ�s�uQ6$W�Fu�
�'�J 8�O�?q��X�$�_�Z�
�'~��	���
�δ��+M!.r�P	�'����W�c�`ٺc�F�,w�	��'`H��`Cč�^�H�o�m^��'����fcÿyq���B.��4��d��'I��@d�!`W��X�c��^�J� 
�'�Nᄍ�B@��$ŗ)�4��	�')J8�(�(�	��`�p]���'o�՛�Z�dJ r��CfH�	�'pH��ܖ6Y -㦐9c���
�'���
Al�<fp8�eO�>p��	�'|��dIL��	-�jF��
�'ᘱ��K%�,���fþ�(
�'aC���] �0� ��T-Z�:�'JT��A�g�L��O3lVYy�'�tPZC�
�]<��d�ޏ,e��'��Y[e��3�:��``0#�'
0 �B��	��ÁQJfi�'v�$�%��� _�-s� ����Y�'� ��v�ֳj#�1�aͮG����'�F%c�F��X�,���O *ph�'���a�E��2��U���2����'ז�9�d&=6�(�5`�Ͼ���'����F�	���`�
H�i�'{�a��!IC��"��#G��M��'�{�Jp�H����.CuA��'��$j�)ՌM���.��$��'���k2b�P`�$bfn�"<uf���'����g#Y1��u�C581�9S�'�B$��J�.a��ьDT(l�
�'�� uJ�,H`x�'ݔM��'�����ȬC�t�B��(g���'�U���O9��рr��KP��
�'�vd�GAM�3�:I
�O��W����'�.�2�/��&�h	�����X{x8�'e��������p�ֈ��9����'��b�K�	��$��[!(��D�	�'���ɔ_6�X`�������'����EӮZ3������L������ Mjc"��T\t�D5%�4�s&"OT,;��A,l38����X����6"O�0����5�Ȉ�`:t�T�z�"O*��4�E"!|���@�
W�*�0"O�5��=Rh�e!sO���"O���7=n���!& �+D�R�"O�D�5#>Wr�e�w�S�K����!"OX91A�H2S����=_��͚"O^ȉF�Rc���ڒ�����ȓVo�9��''T�li"4��S����}،*��H1=����8)��T�ȓ2>u갯Ģ}�]�F̘19P�ȓa�vaXj?j��(2D�(�bф�o�^�%�O5��Рq�:@����E ��#aW�h�U�4mG�o��̇�z���g�>|�t�������ȓ9���ڔF�v�H!Z�h�_�x���v8�b�i��RՃ�!����}ǌD;D&�e#������9���ȓL�:u$ء
��E9
��r��m�ȓa�T���>n��(7��4 �LP��s�&�0�H5-Fh�2B#
4y����ȓ>�,�	�K��<]BM�G�1[#����|�d�a�GѾ��#�	:�����4YܱcM `gL�	�/�=i3���diJ�04!Q�dD��!B�F�E�D�ȓ3��q�"Գ����	�+ʲ��ȓ}�Aږ���a d��g�Z"R����ȓTW~s^�Z��t���ܸ@p���ȓ'%P�� �A�5!�T�S�Q	�6�ȓg>m�S�7F�`A9r�M,����n������|�28)T\w��m��+|� pB�F)58����Ҕu����X��&'F9T��4��	�l���ȓ1�䈻"BY=��*w�FR�E��+���2O�"P��4�`���<�|m�ȓ0�t#u/\j��!e��(a�P�����w�Մ,U����&ei�5��5r�I�2b^�d`�{��P7kL<�ȓ)�! �%~x���6j�+iX5�ȓnD��W��}��yRԃBm�@مȓ#��8�f���L����G�����ȓ$x5XG%��7Ƃ�)�͚�rlm�ȓj�z�D�A"+���bY#����A.N�Hb�C'`�<�x �Zu>L������ֈ�t�r�hcC�	0�z���b�t�%mK�U�¥"!�`�@��Z�t��-U�C����!�*�l���
6t��CI p�-� ��v��ȓ-P��C������n�9�NT��P������?%��a``I!b6�����*�����q`�[C%L�ȓ ���橄�n�]� .I{�ܠ�ȓ�x��ģ��a1�9�'�Q;��e��
ƀjiN��)tb�Ic�Ce�<�"�{$L�&�i_��ʥA�b�<YJ��tۚ��N�,�D�^�<AA�<1�Y��E� >F@��h�R�<9�(�A�����H�*���	��Q�<g��9�����?.��<�
�N�<1ƠU<X�T1�H�a��H2kLG�<��M�il4H���!�jEbb� }�<�3�+:$@(���={�V�Zcc�{�<� �����dNJ�z.��ŕr�<� 
����j�4��t�B�)nd���"Ob���M�<b�BH;�K�Q�V� "O�� !S7*)4HʢDH�a.db�"OT�B�!R2��pq#MdQԝ��"O(x�6Ȋ?���bud52�0�"O� X�� .F��� j�
��`"O�Th�`�+3k��	�	�/�h) �"O ���H�ejH���/�6-ж���"O�a;T�S�l�^DA�#�85Uٛ�"O�r��\8� 8�߅t9��"O�LX���<7ZD0r��P0ZĐ�'�>�[��5A�X"6�I��n�H�'?r|�JKij���AY�^�*\h�'����D�<!-�Ŋ5d ��'^5@p���/}"P�t�R1xHJ]�'��� �j*>m�t�E��qx����'���+1dF6`[E����"�I
�'.���pJ[7!�@C��'<�D٣	�'������?J�P6M��:���
�'����P�G�X�|K񌇼�b�+
�'8�ػSLN�7��Z`K�#.�
�'���	�
���A!`cɆ*� �'d�	aO�!]��	`��T	"���'��I�%�ы�&���G	�`�0	�'\����##�`��t�P
^��R�'Lȼ�7�,_Ā�����N$��'�.)�ī���(�SI������'�&,� ���y~ԩ+ïÓN=a[	�'n��P���{UjD��I^�<*�'1J��UcǢjp�,���ʥBrƘ�
�'2�6��A[`rw)	�7]�QH
�'�� I�gT[d��sց��:�B��' ���l�!E�$&�+@�1P�'7�T`3d�=x�8k�ٚ�	
�'	��3�5���ۄ&ЏKJ(a�'�TH��"� ��%p�І>	���'}�8[��\&9�(���+��z�'8�ق�7I �rãP�
�^P��'����`Fܸ�$����ܿ|;P�8�'?�H�̀kڠ p�o����'����c	Q�H`�v�̷9#$@{�'O����@4F6�� �+(�,�3	�'_�;w���c}j$`WDJ�w����	�'c|I���A��b�(�q|�a	�'�^�ŇN�D�J�Z��6nX])	�'�*}H��߻*�|�`1���y�z��'�f|{�+\o�@h�1H�w!�e��'�쀻3�&e���a����T<

�'�B���`��-!��K�l�
�'�5REM�89Ik��T�װ0�	�'i����N�*ۅlJ~�FA
�'� }� �g
��b���HI.�I	�'�-�g�BEL� 1�9�Ɯ��'������2x�4���ڽH��i�
�'���@D���F�r�l�����	�'V0���4ێ�����S��0	�'.ܽ��W4t6}�'�U�=zh��'o�!#ե�C���	���,�
�'�XӥJI^vt�q���
TSĘ*�'�6�B�L�@�#��w�b0��"O�q7ƈ-�T��ôk�X��"OfX;e�؄s��h�ꖺ�z4"O���v��nF[��U	W��N�!�ք!a��S�-$�le�#�1n�!�� �X�&�9f��z"�A��Z�"OP�1F$��0� �#���\�N��D"O�b�6�$X�
Ãy��X�"O�a�2<_$�ɤ�ʗX|4��"OR��$jEax��jȒ~va��"O(� #_�xв��go�;��11"O�D�c�њ��" �
	F�$�S"Op�x�E��t����Ȅi|���"O�a��íN��C��տlA�=�#"O�}h!�T�Kh�\چ��;"t��p"Onl@�9ީ�P��t�[!"OR��ǣG!;�=�̞�
h���"Od��4(�Q)�\��kR&W����"OT�:Û1YH�����/v���"OLi&��	d�Q�@��6-�x�"OB1oK'#׊��׮5VX:<ɷ"O�qiW�ڌ��GL׋?��"O�,
���2�p�׉�;2���$"OrQ�Ӎ�5\d}�FـX#��q"O�u8b��)s��bEeQ�����y"c��
����'-r.�2�4�yB�I4]$�=�WD�%���s��	�yb�O�ڔ�TE�%Q� �������yR%�|WDYdbO�N4�Bm��y2$̉uAv��H�M�D�)`M��yBND%�@U��o��Y�`���y���D� �&�@:{�b� ^�y��+6��(�T�uE`MS���y�kˠ:[����Ѷnv@-٦D�1�yre�D�\0�c���j���VG��0=���g�,5S�	q��6͐j[�X��_ޠX���L����P$����������I*b�譀T�Ζl]�ԢÑ-g����m:�����,g�RQ+uU�u���X�g�T)H��/eA5��A8�=�T"�Ɵ �I�GM؜�Q�ϙ1��!0��[R�����ɟ��'=2]��E�$�Ҕy�z䱆.9A��s�Q�Px"�i��'���:(� ��<��ش�M�T�i}R�}Ӫ5Y�DP��u��Gy�W?M�Pnσ~��H�!��0��,�麟��	ʟ��%cf�Iʟ�%>�X���< Ԙ�l�5iI�%:���kAR�=�Q?�x�kT�Z� 0�%�}�����#�	#(����O�����'5 0"D�?u��1��Ǔ9��P�|R�'5��Y�$
t$�!?wJ��@ -Tj��p� \O�o�ßh�'�E�C�C�8<�V�͂d�z�A�*_F��'[�)���?a��M��%��|)4�X�3%.��"W :hA�OH�$D?���K���K�,F�'� T����-�֡�'�@����C�LL���;�n[��0�?�Ҟw� A���t��{@&�N����k�O��P��a�I;X��>�FD�ԛ�l�>cZ��w(^�:J> hD�'��Ia؞�Eg�K5�3v\�ެ��)<}2<O�7��On��ͦ�O�r�iB԰�t�!6��e�$옒.�$�*�'����.jӂ�d�O�� �4��6�͟RNK�MN�r����QĊ�4����2��i؟;��T�J���A��VL1��p�V+o���t{��.\O�!�c'�:F}��(��'eq4"��ix����?J>���?aJ<i�/B_���7��hQ�<�'�M�D<�O��Cw��63)�9��!#����T��Οd'�b�4�?i/O������oZ3z'�}�%�kT��I�+Bx�4���?9N>ͧ�?�v���ē�d5�¢�<	:�����!����ɑ �A�dP�a@qs��*k��yK�@�%S����G�fO�zB����?��B��u�cGP�NL�"cұO�΄K�+}��'��	W����'Be��s���8��=�WL�9[l����j���ēF���Qc��:S!���EО�M�iX�IY��yش�?q��Ԣ3P
��s$�'q��Q���~B�'8�-ǒ ��'9�d��Y��m��GS���إ���'~��C� '����S�|c
����_8��m =Nhc�p���O��$YW�S^�diݓVꮠQ"5{b�<�vb���\��{���+0ޥ�ܣ6�;O��d�1��B��0��4M|�Y�� �͚���
rك��"D������Oh���Ox�O#=��G   �