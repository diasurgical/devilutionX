MPQ    ��    h�  h                                                                                 �gI=��	�#�V���u�xl-?b�_1i/\_�y��
���ί"��~n}��h�2�j�)R��K`�hp��RZ�ҥ�1E/9���.���p\[�\��1��%w�%x̝!P�? ��
 �͉}N���r�O��5��Hr��D�⧳�F��7�;���Y�I~vaT:c��i�(�X桿�
�o�4K��ι��k�|�x5�u=>���jP��z�hU��ms�ҩ��]�i �iu���q8i<%�an&b��� Vl�	�5A]��ߞړ��Iy�7�C:P���Nw�fՁ�Mas��D��B���~/�;-��KE����*���a6��`�cC��AIUZ9X�[�D.j���R�1�\��}oI>XQ1���B"�`���ONw����%��|��$�L�@V�WQ>^a#��[A^+�&��� ̼?�;@H^���4R3Byp�6��K�DHG{ł)� U�J=�8�	�'mJ��C��	������.�p�ݝ����.!3�f����'�q-����W��<�z�b�}T���2�}�Y�V������g�g'��N��Z#Wʱ2���m]������wQ���g�~�����U@���m�$�Җ|�5h���Sɟ�\�=O/�Ⓐ�A�r'�C�܄�?
̕����ُ18lrl��x�@�`5���@�Ob��T�Rp�u������z�E�J,X���T�|���"���)y��ػr	j��@�J zy��Sy�U�@1I��D�����嫯��&M��n)'���z�oö/�(e�u�3�v�H���0E@�,l����'y\�q�5��=�6f�,�"��Q�O���q���ꉡ*���ܘ�d�4���^`%]����-�RM똎x�=m�A[���������T�9�/��s�	�Q>�BI�Q�k3�>�z�Ɂ�)��Z�n�<�pa6:��xpE�_�;���^t5<�:�|�*���f���C�31n�k��;�C�&�*��]�7K��)�~�!��#C�e;,4Һְܶ���=QWNV�9�˗�!OfHxV'7H.���f�Yu�[9��m�>�G{�O���|C�T��f�`����h#�TPО��tҲ�̆�xo5�������w���/�4�xw�ao� �~��]{m9�p��ÇB3��z�Q�V}�>�N�>аN}�v��$QB�Ә�����$���dg����ƾ��z�Og(*�o�$��|��m����{b�E�]O�iu_1E��D�����/�����J����U>�h�d���-�`����\��˫���uZ�9É/z'�k�ߣ<���|QT� V�@c�!�"����!7(׊����"ud$_��\���G�-��@�s(<i.�WՉ�[��\2%��)Evbg�2�v�a[Y��`0l�%�,��9,Q�.��O��J1�[P�m��'9b�>0�@/ML�k7z��9���o�6J��vaS��Yd�S{�P@N�n
�i9��v�M֏�H�q[
��^��Wvo�^&���{E�1�-��:�iQv6�u%̶C�;{��݀��R*��k[Ò�9Ȗ�1t�rS��E&&#�������YgA�vI( ��.gXQDGC���E;���+�<]%��N[�^��� �9�S��K�Qq>�o��ąU3�E��	�]+Ǻ[����0Ң�!⇅�?��!��d����0��	��}�	��:�O�Sϼ��+&�;��S���gh+ң�*���c�d��|�O$��YT���-��	�˒awA�ZlU_L��}f[���A� &S/	���7uUOޥ���or�§ (��X#�#ys�2Il1�/e��x_�tk�"�jb�Vj9�����<��>�j�2#���n7��&mFѾ��d�~�qaϬ�t-�P����XG�C뚩�(���7�������^E�=��+PcDtL����yW��dБ\�/�|���Bۛ,q
 �������f���<���,��zy�[}>��u?r�7�>Qa]ہp{�h
��ޑ�\G(o$qs��\��q��i;l0�b��^���$K�In����qY���c|��ݐ��p���pAU�̩��]J� Ն�\p5��`S�z	��,s��rR ��u���'k�S
I-x�A{��c�r\61Ͽ�tذ!�ﰿ��XwTǥY�]��/�hJ��W^�(��L�-�>5�=�V"�^��}��+�X9cȞ��v�؞[�Ԗ�C8N{!��n�5�;��!��)���\�M^ݗ��O��1����Μ@��-/TQ̍s'��o���� �=6=��媹����;fHΝ� ��&�5"��q���S���+��t[��.��ɛ�o��'�-�	��Ĝw�,���R�le,���]�ӎ��*rw��\��7�ۛ��Eu�����o��a�3Vh�K���j+��}DO�"�z����M@yG��*������t'	T�2Q��W�;=�65�9nW*�]�\��ȕ�谳��W�X�M�`"�A\�Yw˽�G��á��t������� R������
v׫�q��y"L߾F���e������lZ/��!��*���cm�dƋ����%2��8^"�4B�O�O�&�ݷ�y2ڛ;_�n�O*�e�Ym����V���c��Z$�O���f��{C��^�e	�k�UVZ��� ۰E�C�c�jc���ZE����Q|{�y�Y�b�Q��s��F\p>�1	�\��4w��'�i2��fS�xc�Eg�X��_\=�\�^��2"�hn��w�M;׈zsc�ՋU?�����0�S�R�1�O�)��K��*��ڊ�	��	��y�_�TAg�O�6bP.��?�Z �@^��{��*e
t��F���!�����K�SF��{��A����ȅ+5�#	t*�>�#����x�����XH���7�:%�6F��(���wu)������Tu���( �e��Q#n�$9�#g�}�P���YM�m������`O��!����=�ݐϊ�ϸ�ϷW=\;�=��蚂�� � �A�"�/M���#g���/$��Cͳ��~�W������]Nj�p��lL��۠���U����6fӡ�����RbU�����/t)�瞱��5��\��\ؾ���`�P%w����?j�o��=��N�}�4���y�ӊ 5�bzHm��D3�
�b�I�Rw�I�8�4��~���:���i�!P��ݿ�.ء��W4��"���w���M��u8��j�����U�ls�K��( ��S ���"8��,EiW�7a�d���uV�F�>cAX���s=��L&y�i�q��t�w����JM\���OmB�L�~J m-a�K 
��Χ��XMh�\G�Pc�[�Ad�9�͍[r+�.����g',p�H!go��QLг��`�]VOJ�-�s%�,�Fj'��V`�i	#sL�[|4��o��pg��L;ػ�y�HA��3�
��3�($������EG6�3)��&����8��N'�6�F��������I�Z.�9��|��ͪ'32^W�2м�l�+����a�?+����ж�޸����n��z2g��p]�.���եG��3��]g�2����w�?�">��%[����0���\m�n� �|-�w룶Qɺ6��g��
z��d�r�!���b�?ei3����٪��l�����
�{N5�˙�;�Ok*:���T�m�ۍ�18�����E,�<X��TDp�Õ����_������M2Ŏ�@J�EHy�6������/&D�m�ҹ#����F	��xl'25uz^��J�eh|�^���y��U�0@,c஛��oyS�qP=��Xf�F"|�Q����J���Mw���15�'��v�o^����]�0� ��R'�/E�=��[���Yr�E�,�o���:s��qQY�0I(�k�]�>@$<�dϷ)�Ė��	���TaQ�a�d�rp ��_���:�57Xy��
*�n�fi9p�K3�Gk7*��������ܸ�K�8o)���!ECƑ�v��UeT�ƟP�W	#�9�/G̜6HS-@7��*�����^���tŞ>�n���&�m�CzȥiQ�[�S���#�7������O�����7ĪNQB��qw߬+/s����ɤ�7� �V1 m����Tʇ����5�3g�ŗQP�)0���}(�����.���?�?�-���$�-7����O+&���Ov
n�i�?�|$,&�����V"E-���zX_�����q�7�$���A� �U���h�p�du�����ޱ��E��>6ˆ�w�GEZX��*�b'�L�^���#�Tt���=��\�b��I��+�7�V���/��MXu��F�g���g�-�-@���<ĉ-��É�Ɓ�Rܣ�Y�v���2i	�aV?���Ձ������nM,�MШn*ї
����M�mzf���_b�1�4�KM��k ��\gS����22}�D~an�Yߙ{���N���
�=;9����js�j:Yqv3�,���3�o����g.E�+�L:��vQ�%GNlC��{u���z�~/��yB�[~�29�1�<S��K&a��⢿Ƽ��!Cg�~�IC
ܓ[�X,�_G~C��0�p���/Jw+eNv��u��vS(K���[,�j���R 3��`[�	!�+���Ϊf��'3�	*}���?�Li!���r0���DV�}a��5pu��"��h�&�����}�B��+Fv�����^L��O��
n������&���a��D�/���U�a_�L&8;*��M�{*
�c���U����6oͽ�b�q�ׯ������ӓl�He��xZ*t��a�[U��q�5�N�%���Q��`j5
Y��Y_7v:��������d�N��Q��犮-{�	��\vG����d���r�v�����ۙ+=�JP^�YLEt����hÑ~�j�
�<�H��Bv��qL�Mx Ǔ�i���<�;Ӹ�1�ŸP}�}9y[#LDrn٢�Y*�]V~{������Q�K(j��$�t��jq��6i��E�=�u^֦���IiE��+���M�����s������ݴ4
U�$��YoiJ�cl����5>��S�؋U�x�� ~���Zm�k�!�IH�wA���cx�k6l��sm!�� �D�w �Y��F쪍�h%f�W�3P�]R�-��$Ϙ�="���^��{.��+��:cS��y�ؙ����C�V!��>?�;���
3D�h���H�ݗOٛ�1��d�J#�@��/����nH�����e��*]6X���%Y|);��G�����������m�5��Zo�	���Ё��	���K�o�o�'��t	ʉ����Mcm��"�e�_�Xr}.i���'���%�-�vhn��uu�������7���T�f�^���j�XC�]s�z2��HQ3G�%'��>F�޺�t�T�7�ߒ!�=����4J�W�<ƪ�b�)���-J1�y;��T�M�:�`��\��F�x��+@��E��ó3���R�8��U�����f�ٹ��LZ����&��E�Q�r��/�w��Q}���Jm=�i��:(ú�i%�' 8Y*�4��6�
���Oy��i��n�'�*E�Yh���ʐ�Pe� ��$(�{N�&B�!�e'`K��Z�%����EUgjc��@�(
����u�b
\�M{��Y�m9Q��s�PKF�i����1���#茇BFdiM�f��x>�kg�\�����=�[�߹�2�fYn�e}u";�}s�[�&L6�����":gSF�31�.)��+K��"eU�%@�	�M��B��_<ОA���Ա�P	�?�ʝ�*���c�0�Y
/�_F-"R��p{�/sK��_���<(���R�+�4	��UoD#o�K�:����^��S>_i��7>�!��ά��y(ܣ�((�u�����J���U�C�Ȝ������#�v��Ȱ��垔Ȼr�=��{� ٜ�n��%���6�O��&gW���H?��ԃ�i]� �-6�]��M�D��5�g6������^���&��2�O�/2|]�#|p���l���[���p�G�,)v�|����R)b��J�Ü�/��g�YT��P��\Q�ؙ�Ǜg%�ٝ64?Ť4�TF��4^}D�	�m��Řg5:]�Hh5D��ͳ�n�mGˉĎn��~�}�:�^�i�:�7��sr��l4A
F��u���.�����u3��\X�j�lɦ�(�U�G�s��*�c���v ܧ}Ƙ�瞖ir'�ado����V��J��AS���T-Ǘ�1�yG9��wc�w/۩շ�nMW݆��3�B@�7~eg&-�\�K��m�	}\���e�W��s_mc�V�A�R9c�[Mpn.���9'K>��[�o�)�QgV�8��`rM|O���@�%���ǡ�'���V"��4��#N��[�*Q�\-������r@;�W������3������LM��ۏ�Y�G��)�� �@�8u��'�B���J1�� ��Pî�K6\.�"�ݓ���F�3mu��Ω�g���y�u9k�\�s������c��]���gY��+%"Iv��PH��uD�H.�]�G��\vw���ݐ�Ϯ���m�Z�+�mFFo��-|�:��^����ˏ�3���eR��	��r]̼��`;?�&1�lX���lhS���׶^�5+�$�6`�O��wt�ވ&ލk ��v���A�E�+eX���T����P B����ϼ�({Ў'�J61Iy�`T/%j϶$�Jg�D�YI���k�,l�\����'���zy�e�He�E�������P�0;
�,�tțJ�y7j�q�
���fM�"$�Q¯e�S��"���H����k��f�o�]ֻ��[�'R�6��J2=c��[d�����������E��sLk�Qt�I��kƨ�>{�q��<�)����$J5b�al���߶xp���_0~B���52D��2v�*uEzf7���3珬kr�x�y`��x����KV��)��N!�[C��4�����PҚ7����W��9	�^�>
H.$I7��R��2��ï�/=�>,��z�r�CXWP��ԸV�G�J(6#h:�3q�j���F������@b��f�w:�/.0���=�W � iN�T$�moZ���������y)�������F�n}�Ṑ#ˌ��&�����Z���ZD��n{C�4��[}��O��S���Z�}|��
���`��j_E�tֽug�_�F��G��-b;������r��; uUtӒh�J�d��ӣ-A����R�<�aJ���aZ����%�2'p���e��T�UI��6k���)�$���7�ſ�����:�5uZ�ړB���9�M--[|@���<$m�Ͱ��vV�R�_�\��v��2��aQE������W%���I,G�]�I%�E����k�mu7���bf��OpM
�Uk��?�)���7vMP��?a�P�YZ�{_�>N6'�
1�9�]��Ź
�%L�q�|��d��/�o�,��x8Eҁ��5:H��vl
%�1C�i�{M��ݶ�[�y,�����[99��!1j��Sj'b&�|�=������|Ȕg�1hI^����X�G���{Zo����!�2ihN��l���[isSc���f��e@�;p�3{��{;@	��+}@<�	Y��f���S�;_(?Q�n!3V��~%0r��|}����0d��	��#`�&��H�I�>�=�+�:��`6ܠY8���0��(��{��U����qg���L�P`�_��/������$m���L�
U���ԋ�o(�s� ���&��@��|��sueA��xU%%t!���`���ڹ�9Vۺ����Oj�G��D7ф�x)��7�dv?��_Q��"�<-�V��pGO��B�/(���6@������1#=*PY&;L���p�^�!����Hʳ�����B�q �Q�C�N���<�#���{� ��� �}4��~B	r)��t#�]њ�{����
�Z!(e�!$'�M��c�q��i1ǋ-$^�~ZQId�Y��!������E�%אm���P��OkU����J;�'���5���Sy�֋H����T y=����k<�Ic��AqHHcS�6�U �-!��,�mTwʘY�]��%!h i�Wԑ��w�-����"U�^h��s�+d��c�z��xBؔ�f�L.C�K�!m)�h�;�+8E���^�C�\P�O��1���ŗS@���/�/Y�����]�:ߏ�v�`6s�q��W�;�<���ְ�|��J�(���ā��.�@j��e��dFkѿ�oS?f'f�h	��m!>rv��)eb���S��c�Ҡ�ش���XJ�Q2|<u.�E��|Є�<��ףсx��`���3ڧ��)xz�t�C��GRv��?�L���YtV`��<b���=#���/F�W�ΪҼz�Dzɕ��ݳT� ��xMG�``s\A���3W��F頡�k�Î��N�FR>�����Y���!�%��QL��Vț�'��'��Ѝ%/?t?����Zm�	��_�C����%h��8TR�4��=���ځl�y(H�����n �*�DYc���g���;C$� z�VV���)E�te��0�0�ZNN��6;�EЪcr���c�������J���{_�tY蘖Q��s\��F҂j8 �1���~�B����ih���\�x�Ag�aŕN=�z���(2�0n�f��F;��Os�;���b�����}c�S܇1�)Z�K�Gm�J����K	����S_���A�Z�,��P�K?5Ũ�vK�_跋	n
�CFH��v���KW���
)�7s�L�+���	�PI���#J]��u��Q!��NT�ĉv7���F?�+�(���c��u_���+�
V��C 
�KE�G���ڄ�#�y�;a˘���#�]�7����w�̆��SiR�궖��RW��/ag�-̈́��G �9:�tfMP����v�g�8��]�y5����I��j�F]���p���l�;�◹����;�W\Ӧ9�b����t�/*�I���k��\�[a�t�����%I�s��$? �9��C�9�}�e9�H��� L#5�wHc{�D�
��p���7o�?����u~'<>:4��i�s~i�ֿ.���G�4�Hu�_�����I��u.�B��j�[*���lU��s��s���!.h� �v��t����i���a�CN��k�V�r��AN1�߯1�P6�y���8��Rr�wj�h�RMRB��U8KB�K�~��g-W�JK�]-�Dr�f��RA=�Ύ�ctqSA�KK9��[(�K.���	"FI����ozϬQ�j��â`M]�O�#�c�%~y��T�}�gV=�^��#)�c[�@��
���r*���o;NS�(?7�^3�J�!���^���IΏU5!G�9�)�C���{8P��'o#�|���'������".,Z������3���h��b����2�0�X�����Z��dU�.�֚'����Og����dUM��
�[�e��{�]�������wb.xʘSϙ��v�����fMm�(��j|��V�����������@�8�D%r�����~U?��'���_l��*�m����̄5���1I�O!�2��ޣ�����Qw��+��Eb̥X�a4T�������,��v	�䋎bm�J�<�y�߮���qN߱e�BD�p�����g�����}�'�'^z�-����e^�{�Ļu���g���06,)�UyR� qF%o��y�f��Q"�p�Q��s� 3o��쏉�0+X����y�/'7]�fV���R~��e?�=�4�[?|��]��{�d�;�@�sLQ�x�I�k��>����ʄ)�&���Taa���Z��p���_kO �p�5-PK׍/*0<�fR�bf��3�P�k��%��W��O%�ne�Kx)�I!���C|I~�ҋ��<��6WA9$X�̒e~H	;B7��n�����@��l����{>G����F�MѷC�T쥵��Q�״�_�##]^!����c_�R�)(~��P:��iiw�Q /��d�Fz��(� Df��7m
�V���k�S{_ګ�#D�ōؚ�ߕ���}^ǻ��	��a8�<�)�u:����)�I���o������EgO,��[0J�u�	|�����,�PEc0�p��_B;�u!r�Hs��-�@�z6��v_U��h�D"d+b�^���҉����<����qZ���� i~'�8��ԫ��*�Tj ���P0��sę���+�79U�GD�Uѻu��K�t�-�@�$�<z�쫈�m�73����7vI�2���aLkv�q�ͷV跙�.,ר$@���M��,��mp(�8�-b!2��j��M��k�k8�z>�����шÃ��a���Y��,{:CFNq��
�DQ9��^�  ŏ�}�q��"���K�o6��͝��E�#4�>O2:@Qv�cp%=�aC{0'{��G�Qv��tI�/�[�	9��1��tSE��&��p��H��l��ׯgrIy>q܉nX�
(G�o�f��c�M4T�ƯN�ǟ���}61�S�� �"���`�wĖ�f36i!�;�	�+X���D'@�3<�������$?�!NAt��s�0M���}��%�+x�d)>��^�&�]���!,��:+�����ҠT���Xp�a`�=��:�s)yֺ`s�2���K
�_]���Dt�*�v�qT�����CU CF�� Io����؟�����x��F�x�e�@�xPe�t|2@�ъ+���&�D�2ە��8tjk홟Ou7,��W.���d�O��:q��]�-�x|�{�EG��|��!��J���l������X�=��PT�L��(�+}(�<���t�5���m����B�Edq��/��	i\��5c<y�����u�;J��}/Ǜ�X�r�|.��<�]Lׁ{qlF�ETN���(`��$��ē��Dqٍhi������^L+���hI_�d��V��Ì����v	�%�H�!�D��dU�4"�~�J�H�܊�54�ST�����aj t�����k��I~gA찪c.zz6�Ȟ�Eo!�5���aw�1�Y����2hۋ�W�����-����N��"�^1�$r�+?b�c��ů(؏G�ԧ\�Ci��!+��4�[;q�K�;�ʞ�3�>�����qOO��1���@,!@v�=/�ݍD[!{���x��1�H6�=R��~2��;���um��5�F� �����>S��4�%�����Ѻo�.@'!^�	 ��薔���e��0�N�|�}��[CT��ӽ3�,�mGWu�่�˄�"�d�Wќ�����d�U|����zhS�>ӛG�������3t��x��b���=��x�*b�W;Sw���6�_X�#m��/��ʼ�M�q`Gf\�L&���ԩa���;X��i�����R�Վ�ʙN�~��ܮU�16�LP�v��*�����/��΂Ǭu��h"m3�T�:�o�0ߡ%qW8O�4Se����.��y����u�nG8�*RdKY^���ů����V�c$9��1~Ǐ,M��W��e����Z	�ޖQ��EK�cM�L��F�+�y���Jq{�Y��Q��s7,�F���`�1��>�ٮ�����i����4x���gJŬ�0�=���o��2S�nևak�w;h��s���\�,��͔�ج%S�P�1�T)��K�Ƨۤu�[c!	��2��v_��@A�Q�ԧ��P��?p*��$����樢
���Fc�]�������K�DJ����2�q��Ǥ+f�"	�0�#%�������\�I��|7��F�����l(�� �u�S���,��evQ��KU�����֘�Z=##�����]��~2Y�d᱙ْ)����Ύ"���Y��3zWN_J����9�^�_v me���M�AM���/g죤�`*���ʥ�������v]�-p���l]����9���|�"n:�2��t�b&_��l4/��K����Ɇ��\G�e�O%��%�Ɲ��?{�~��-�9^�}:.5�#�d�;35p�H^	�DDXt��i䑣G���������~b:ω�i}�����Y.��Bs47���:���W�7�䷽u)�
j<j/���U�zssfvl�ٜ5��b �e�3C�]�i��EaZ85�`�UVX�����AI�s�
 {�[y8h:/x\�-��w����oMM�G�\�B���~��1-�QIK�7�����)#)�M�"�)�kc/��A���9�[ZY.V�Y�81�a�Y0�o5��Q����.�$`(��O�:���E %y_c�W�H8N=VX8�*L�#}][-wG�����#��(�A;	�^�{��N�3��S\��������܏�0�Gg�)
Y��6�8+�'Y�;��<��n������.U"݉R�^�3�ҕ,��]��/���*����i��a���i`>��ܱg���TB�F�a6�����R]8�9�茩w��T�S���N��	�����'m|%���ݳ|>�&�ԯ��V��)q��B���r����ȼK?vM��'��q�l^���H)d�,[�5al#�,R�O|C���l޾\��a�K�,UU�fT:E���X�5�TU
C��]��8�>��bQ��l����Jlh�y�~E��,����IFD~���c�k������N�xV^'CѢz�Ҷ�w	e�s���U�4HC��%01T�,t�����`ym� q�_Z�� fÁ�"MݜQ���[2Y�~׹�sn�����D� o����W]�1��RR9j��l�=Y�[\��
9�����:�0�s�L�Q��jI���k|�P>�v9�5x_)��3��*.��-a��c��c�p��_�@R�$5(|���'*�R�fm�3�I�3�1�k辆ͯG���F���;vK̽")�"!y��CW՗'�g�&�O��.�a��W:I�9?���^H�q+74�~�TI�����*���p>bDy�pن(��C�q��PW��LJ� ��#ޟ <G��`��:@L�dP�����ی�w��z/����~�MQ- ���j�m�o������(X�fG2_Wr�L��xu��^}�̵�uD�?:�����ِ�Q�P���$wƪdp� t����O����0�-�|��X�am�g��E�>�k�9_�>�0��c�g��9A�U��oU�@�h�^�d�]�����~�H������]vZ)@9�NF'&��ߏ��E��T�
mЬ���_�����37�)���p��uP:��/x˯��-cJC@���<ո��C�(�R΁Htʣ��vNԼ2:�NaG��̅����g�,=P=��zޗ����ymk9���b�mL��L�M ��k�Qf���j$�@��%,�փur�a�l0YP^x{��N�_�
Sx09{�$�{�?���nq�n��P�Z��oq{<�8�UE��B� :��v��>%���CVc{�[ ����o�
�wR[�q�94S�1`�S +�&�y�s���t �2��g-��I������X�G�G/HB�����f9�D;N����w��]Sٔ:����[\���
�3�q��[X	x+�+3F��[�����7��O�?ǧ!iL4�t�0(T���}2���&�������}�&�S��?�E���+�"#��-�O���`6p;\�5g�>�N����oS�͑��Fԯ_�4iy��ERX��7�D#���pU���ʕ%o��Q_f�(u)�#=˞0k�ew�xK��tב��ն��2����p(��s?�jQK��z�7�ys��*27dl����9Ϙ�T-Lz�v��GYm�����e�����qv��J��=`�PO��LV�:��hv�W1͑ﵭ��ކ�wBG�Qq��n^:����K��A<�G��1 �vm��}*�4��r�~��ua]�3u{LX�����Q�[([ʫ$�8�H]�q��i'J��:Q^��M�q�IZ���<��~����/�� �#^\+�݅B�U����j5OJ��
���_5�,5S/nd���,�I�7 o#�k�fk�J"I�L�Ag9�c	z6\����!�g�#�w@�Y	���3h�ΟWJ�~�.#�-���ϩ��"�a$^L�����+P�c���J��؊+H��DC$��!F���R;L=����9
A�9ZG�M�O
I�1Ļ�:@Q�/@�6���v���1��x6�������?;R�l�S�|��z⬡�(�p,��/D����T�`�΢��ѵo	>:'�X�	 ��c,����>c�e�v-�I�?�d���ὖ����p�2�ud3�ڨ��H����oѷ���V��������z�)�9DJGw�����/�t#��8�C�2=Y�%��W���H��zVk��.��
����:M}�`N�\�26˩��|����d��D���Ę�Rt�f��k&�}ח�i�L
!L�\�Q��QL""���	 �/��]��t��'rm�.�����k\%�EW8J4�n��;M�I��y!���n�p�*�7YY*�!������qL$�q���)�g�G��H�e��f\��Z����lvEƑc(vz�ٔ�����]�m2�{ՈYOiQ���s��FH�n��1���4�sb�i�\G�R�x�F�g�)����=�V���2$�n��?��;C�esO�R���+���~�3USw��1�?)��K�e����$o	��8�S�_mϗA�h�"�MP�3�?�����Pa�ŷAh�
`y�F~����f�K�Գ�0��-i����+!��	�
����# }���%�����D�z��7o}o�ج���(m$�ٺ�u�����M���8⹗$���=�i�P3#S�ׅq�H��I<�ٝ��a5��Gk�����[����� U����W��$y��T?8��2 H�����M��3��Z�gGe����M�u������H�]�;p�0rl�q�ی�����b������@���%b�Α��s/��m��`ɡ9�\�v�*r��L�O%uѝ:?����Z�T��}�����)�v�5�HY�)D��W�N�5��wo�5ɘ���+~�t:jO�ixE��Ͽ�����]74�%�����X���u$R7mB�j��ئ��U�C#sAo���d- �t��1��l�iÚ�a�Lh�;��V�3��AD���e��Ɵ�ySDP��-���w���Ո�MHlb��)Bq�2~�\�-M��K�1݃��������H��Mc�jAЏ49}� [���.��K��x�����ʐo�z�Q����$s`��O6�����	%te�ǲ�i�vVs�E���#�w�[h��-&�����̃��;�����U-%N3�v��P�����a�L}G"'a)%������8^7'�'��Ŗ��թ�a6^�|�.8�2�nk�9�b3{������X燤��{����P_�䩃<�rޤ♚]Z��׮]gj5�\<~�s�������u�]����T-w�Q�IZ���lW�Ӝ���]~m�À�p|��6����&K���	���7��1
r.�G��?�k��R	�R�lٝ,�#|��g	�5�ᖭ'{�O׋֢�}��'��+��SO�tE�moX�)2T�}nÁ<#�Sx�l�ݻ����JJ��y�=@�������D�F��>I$��y�-ak�s�'���zJ�����eT�+�z�%�o"!�0,��,���{4�y�oiq<�ѓ���f�f�"�iQQ��c�Qc�9��(�}!��a
��[_;�e�0]���laGR�����=��N[�[��E4���h�؇��gs}mAQ���I;LkWIM>,}���E2)�`�5����~a����P��p�WH_�Q8��9�5#ȍ�Cx�*���f��,\�3x2�k#ۛ�J���]��$2�K��)
K!���C2��b�����S�ട���W��i9Z ̈�H��7o邕��i�zܯ"w�`di>}����/C	�`��;�G�̴[.\#��W1�ۅ��u������QwKv/_���pK�ș� ��X�\m@*~���}�	���!��z�3Ńߕ�{��G�}��N{��2����G٫���_��$��������mnO����-�髓�|��<w��gOE�ƽfT�_��e��4��~�i�#���0���=�UE��hט�d����Ի���a��|����a�3�nZ�C�S�'�a^�J�d�` |T`�Ї��H~,��E��>7�Ӎ��ZƋտuˏ���4��(�-��@�:�<0����!(�m������Xnv�2Փ�aBm�'����i	�O�,�;����m����b�Jmfj��b�b��]��M{�k~W$����j���Y�_��0Y�a�*�Y���{��eN�+�
��G9vR&��Lz�VA�q�@�5�o�RT��ShE�'�����:yv�ku%3�C1�{�=�݇���j�x��s�[j��9O҈1�u�S��&M���R^�����Jg�	�I��{�Q�X���Gj@��L�{�|5��^c�
N�Q^��� JS�ȵXFU�V��L�-3���̛�	�n+�U��#�7�%���L��?�[�!�w���p`0�e0� }���! &��_�T�*&jyպ�����+2GE�1�g�J8��40���P �c^)q��0��h���A�,_2N$�N�`>��g�v�����UV&_��J~o9O��N?��CL���ݍ�y:�X�te��xFE�t2��G@f�����:���K݇���Xj��a���{7�#~���|�Eߕd��&�����7�-��O�q�G`.��PYր�p�b�g�L��ۅ�=�@�PJi�L��̻�tH�r���j�1�v�ކ4��B�VWq�;'�e��vߩ2�G<oA�s�z�����x}%�����rZ�ʮ��]B��{'dԳ�B��E}(V�$8�S�
�q�:i�ԋ���^�/�+K IU��痏O�9�{�'q��g���^��� �U��)���Jl�2��5*�XS
{��5��䠽 j�F�ƶkm��I�Q�A���c���6X��{�!��ٿ~9�w�Y$�얛 h�1+W�lv�ɨ�-���<�"���^g���~+�]�c?vh����؅/��]C@C߷-!a_n*�t;'���ö��e��4)8�m��O���1)�r�6��@,�/{mc�z�Zq1�K.��}�6�UK��複;��������O���BY �����y�Ar����5�$ѰK�odmT'�s	6�$����@�yc�e3~��D�l�z��n�)l���h����=�u��*��nT��l���	�������d�Īu�I z����4��Gc'�pmx�J��t����y|�~��=�aɵ �/W�騪1��t������@�)MI�`	u \R9�dl������1���c�����R��]Zj�/�RHb�g�$LFԙ�,�˷�� ����w/P)�=\g�
Jm)�o����æY*%9:�8E��4	����w�dj�y�a����n��k*��YT}A�x���<������$�k��-܏��F��e����h�Z�Ö��+EA5�c��d�a^�F��:�{��!Y9��Q	{�s��F���	��1��aϏ�$�.�i��7��2x���g��_�f�=���%@�2�M�n*fat;��s���Ւf���A�䎟dS2��1�)�h�K`$�Q�fڑ5	�ầ���_(�A��ԝ�wPu�c?�T��G������Gl
D�F��	��F,A�>K�Q�����(K�]��+�P!	��q�#�<z�&ᖲ")j�?V��ɨ7*^�+��u�(H���u0OP�㎔���tx.�o͸CG�kf�#�� �뫘�U��4)��X���و,��]i���݊������}W��4���o�Y�Un #'�I��M!�r���g�F��#����7��Þ-?�;_]UJ�p蝞l~i�GI~��ѱ3/��A���Lb\�ԑ��N/;���E�ɼ��\=4s���Ǉ��%����_?1nɒ@=��oK}0��ٰ>ӱ%O5���HT�3D�R��	����ˉ��{^�~�6=:5�is�&zX��_�Q��4-�K��l����9Zu���%�j��%��Ux-�s�n�O�y�:0 ȣ�?���E�iޫ�aP��WQV�BQ��pA?�m��R����yn@�%Wk��^�wD^�#s�MC1��f�B,��~�C]-���KgK̓���_�L�C������c��+A�a%9��[��.�Cr�n��ҷ��o��fQ�A��$��`�L5Oq�í4��%o�����OV�h� �'#���[�C��cP���1���e; ����3d<U����//��N�f��G��F)@5��,�8��i'ϳ��M�(��\~�����7=.S������y3Y�9	ϨS9���#aly��0�_�Y��߄��C���g������Ĕ<0�|)�4#>]n5���<Mws�n�� �����J�w-	m�����#+|�Æ�JKD�A`W��}�ѱ����zrɶС���?,\��X;O�1R�lT�����zע׽5�w�"ċO2�}�c���9�Wz@��p����AE3n�X�=�T:�<;a�nN��u����ގ��J�~y�'�^�Ϣ�Z���%Dt+�����i)�7��n�!'���z2�ѯjeϲ��U�廪��]40'�,*0�6�y�Zq�4Փ_w�f9ly"��Q��E�����z�CW5�H��<U��o�� �]�'>���|R�M뎶&L=O�[�{ ��OJ�L��]�Q;�s8��Q� oI���k2�>g���k3�)���ǐ�'NWSa��7�ː
pg�S_���A��54Yמc�*a��f�N��3SS k^e�宁�����HKBa�)%5�!o3[CM;��y�\��▟��W��9u���cH�?�7�;{��\l�G2�}��\f>�)�f^.�փCD9��@ԸBZ1���S#T��r�k�V�!���� ��U?��2`w�8�/�16�C� �m3@1�m�����Їd�i��X{������u�p��2�}/8��G���Jn�m��ƫ<�F~���� W��V^˱�1O=,������|�[W��9���\E4#��a�_S����n��f���B&�Bx�'ݺU�-�h��jd<p�ӏ���#>��>\��͏��n�[Z_ŉxJ'�%#�;��{G�T�?��b^࿃3��O��ݛ�7J��x5@Ʀ>uF䓮Y��%��-���@��<��쫹�k��*f�>�e��(�v�J�2p�4a=��������Zș8WM,3Gͨ�Pm�1p���!ma��IӣbRE�SM�r�kY}r�+��Zs����݃�_�a�XYF��{�U}N"�
�?�9q9d�1u��Qq���	��_oo�I@�n2�E��s�O�h:46Vv�%�#}CE�{9@N�"��e`c�@��[%�}9jq�1V�cS֮\&������䶯�%g�<�I�|����Xs!�G�XF�����8�^+��N����m��H�SO�����{�Q��ħ%!3g�*��	n�j+��>��Q�ҳ���6J���?=/�!��̴j:0�/uk4 }hm��tؗu�`�J&*���5��� =+m��̤�EG��S�����k@!፧�Er�k߄�<�_n{H�B��{JT�⢲Q"��8u�U����So��0�	?�^Cݭ�j�TdK�H�e��xA�*t��~��9��������&�����j< 0��07=���!�`��dbA'�ː���-����l*�G�#o��(֛H4��d��'�x����=��SPEj�L�޻\����W�����Q�o�o:B}uq����:-�M�v<��N����&} ,?�[�r�>��G]�L@{�ӳ�����(Qn�$�[k��ֻq*Z�i����>^����D�IP�m��[���3z�B^:z/[��A�҅�ݻ��Uܼ� �J'�~�-�G5�(S姲�4�A�p� e�>�!�k(�I�v1A]��c��i6��r�X�!�cv�ن�w���Y?����hl�&W�J�dN�-�t��_�A"AIM^����-�+Ћ�cz_�ŀ�؀S�Ը��C��=!|E��N�;Ϧ1�U�o��/e��ɑO�\1D�*ı�R@�/�ld��{l�+��#�b�X6�d�V��ӿ;ȥ���
��d9�W]���0^%��}M�����f��x=ѫ��o���'R��	Q$0�Y�	��7��eΥO�?�~���Ҍ4�D�S���۽i�u�8'��T��E�Z���X��L�F럅���B�z9���/��G����+I��e�t	p
�T�O߹''=�ʕ�v�WL�1���C氲���I�����{A�M��`��\�_��^G��ͼ��ݐ��>&�:'�R�1��o�����>���L�k������X������/��|��c�%�m��ϋ��S���%�N8@2�4d����R�Ty>M�]�nn�@*#�8YO�-�ӥu���d���u$�B��µޏ�v��(�re�f*Z:1L��{�E���c޻&�O�8��f��O&#c�{KиYT�\Q��'s�e�F�'��B01���H[���i�hP�H�2x�8{g�Q��=;=�6�߀��2���n'���O;�߻s�8r�-�2�ϫg��HTS�n�11��)�WK;��s��,s	���	�e_�nRA	���-PP'�?!��	�۟��F
�.�F�,���F��KCU#�f��#�Ѽ��+�Ɔ	E�|AL#�N�a�沽k��:�G0�7�^�F����D(#�Og�u������v���/�OI�8�3�0�F��#�~���'��ܔ��cIo�����U�8J��?�ɊV���YW_��'���Ä� ��k���M��	��yg�G+��Pi�兊�kK��ydS�VM�]�p�*Gln�#�~���Ǳ�����#�%��b�ls���/�U� b���M�\�|��k�����%�����@?��Β�
�Ί��}�G����X[5A"@HOsDU ?����7�+�Q�VA�~uz:�:�in���0ɿ�)�,��4�������]W����u:�#)�jmV�7G�U�6s��w��9��k ��Dn���?�i���a�ղ��:�V	�CQ�A:�t����<�	y�\������wV��վ$-M>���B���~�J�-C��KB�̓0����C�>A{�:��c`AT�9s.�[���.���	h\rηj_&of�,Q�;�t`���O�|L�Ͻe%j�W�h��i V�0��NX#���[�ٟ�c������9�;:B�5�#2n3?"�sG���,�������YG���)[�\��G�8�_L'
`��������#����.n�+������1a3����ԧt�N�ޤ@8�I��7j��x��?P�G-��M���\g �f��z�R��Ti���o��]	����D	w΋�ʄ�;+�bRp�RJR��mMd?��� |O�����\������㬙w�0�?rd2��6W?����D��Lr�l����ف����c52-f�-fO�|��*�d���̫�����EΎ�X~q�Tfĥ��YC��D8�b/{�o�Z�N��J=��y�r�<?�]5a�ьD�/��P�Sx�c.��iT�'T��z�@���{�eJ��0����6�W��0"��,�:J��vy���q2�d�:axft�Y"�Q�O��l�ק�W�^��.	�&�џ��E]�R��"V�Rj#�ѳM=�6�[����������S���>s�Q���I
�k��>��K�A�)�j���k�	C�a�O��FWMpBc�_W����
e5�@��n�*W�f�]�Rh3.��k�s�̀��������~K�b�)@n�!�C�8��^A��\d�՟rG�Wk�"9�(��~C�Huև7�g�%�}4��o�sg>�M��P���C�%�!eP�=2�}k#(���N���c˦Y��c�����̵*w/�Ԩ5=���� �^{�mv���G ����ڗ��go�yfA�K��md.}ʝt�`݌P���(�u��f���������[ $��.����O�~2G�����|���(��E�^~�\��_����a�v��F��
����b��U{��h�l;d�)��Je��>�`��[�˨~w��\<Z�����'7
����#���TV�=�=�忾�0�T�ث(7�ҷ�30���Ydu��ԓ����`�_-4��@���<�m�t�gށ��壣v�5�2la8C���U�Bk�S�,�r����ܗlf_����m\,��c�b���%�Mq�k4�P�f�����}#=�у���a(Y�Bc{�FEN]$�
$�9l@�׌�/�̄iq�b����o"a �	1�E論���:�ruv��%){^C狷{tb�ݽ\��`���� [�h�9�0v1њvS���&ÿ�Dۛ�L��C�g^�;I�&'�u�XN��G����Xr|�����i�}vN\=������S��ൎ{z�L����t3"L�|I	�U�+ľ��0�d�m�����͇�?�"G!�-����0�����}����ж�ʙ&E��հǛ�di�+�淚g�ݠ@�d�q��l��醁j���8֦]쒞5o�7�:_��"�׹��vn�]R,�S�s�U��Xͻ�o�W���^��yZ������/���̓eH3wx<�2t�o~�u1���0U_��î$�j׷����r7��S�CE	�{��d����0e�IN�-Ã�g�6G9���d\ֶ ��X@ɣ�z��0=1�P@�hLgq��x�� �`�]�,�����yB�q���o���h.�<eH�)�?�'B�2}��E�#r�Cw���V]8	{�ۢ�1�8"��(L�$�c�yëqEޭi� ��_��^8�*a^xIK3i�MH���|�]͋��ڐ��!cC�Vp9U�ԡ�{VJ��H3�5 ��S����o��`� `l��|7k��I�{Aؒ-c��Y6��a򱲓!��4�Zwq��YZ���hGW�W�Hµ��-��qϺL)"��'^����+��c�h,�+3�{�m��CU��!�K� >;��zl̨�
}��*'Η#�O;�1_�*�,�P@�_/�9����g�ŧ����6�����g�"�;�&�$|z��	���`w�H�K%��o(a(���0ѢkU�Ѧ�o,�'	I	l��Ԭ3�j��Òei�t�:�LP'e�G�_���[�ۘgDY�u5����ZN�Y��P�����[j�z�/����z��~�*W>G���D*ဍ�t�FS�/:����=*Sz��W� [�y�����3ҳ�@�붭$MN4`�"�\����o���8�'Ju��:��u�tRE������ �4��a���FeL<#���>�s��~����/B���i�@%�mֻ��E��T%o��8;��4�dC�l���^�y���8�n3��*�"MYJ���.�0���}��$��^��]1�B��e�z*m��Z��8��[OE7�c����?����"xS~��{$�YoP�Q��fs�c�F��x?#�1���E�1����i�����x`��g6�Ŝ��=�����\�2?nBL�W��;�3�s ��ȳ:��5f�D$S�c�1L��)wg�K��M(��))	�k3�d�*_��A$n�ԓ;pP+�n?\�-�}�wֿ��Rf�
�9XFώV�~q�LEK~E)������1�+R\0	1���1�#�r�����X���5����U7�Ba�ke(����m�uf����p���7���:�d�	ͮ0&�!�u#�n�B<��z�֔꟧����~�;�K+�z�i�񨗹��qW�x5����u�K( �T���oMW����JgXi�L��� jE����T�W���]�3p��kl���۽؁��F�xTӞ%]�`��b�Q�����/�̔��h���\31ػJ��8r%PC����?����{Υ2�}&���@Y�'��5�ܪHJ��D��B�����<��#�1D�~N�+:;`�iip.0)��ը��Go�4#a�����C�4�P:Wu�x~Lj(嬦R�@Un`;s�1�ŭ�5� �au���IYi.JaFJʃ�>�VD!
�lEA5��v%d��-#y���*���xw�8q�Y�!M9��.xB��R~r�-���K�݃k��U��9���[�c�A!f�9�&[o�p.Bd[��	���Y�o!�6Q	���&`���O�')�j��%e7���$�{V��:u#p(�[����>�н'�̔B�;���65�h3(�H4Q�e�n���/�^�GS{�)v�G�"�8��'E,���`����۟r��� }.�9�us��ʍ3Ϡd�ofr�I=���	�EY�R��U���F��U)e�.w��eg{�K�s��g�2�.������y]�>?��law)��?!�Vlo���A�-���m�c����|�H���f��w�����㇡��k�Xr�kk����?�6��l�g�nlJ�4R��}5�­�<O�$M�����*I��Mwe����R��Ei�RXyŁT���ò�ɡ�Z�����JІ���5J�V�y�:�Q;���+��%DjT���.�����D҅d>U'��vz{�"�hle�qރV6� q;�@#0h`,��d��s�yٔ�q����kf��M"���Q�����oB�j�ʉy���3	���&����6�]����} �R%}��`=E��[����� ��P��iv�:s��xQ1I���k�	�>�O:��n{)�K��Fl!�N�a�,��=�p_�Ec�w�U5lD�T�K*��f���O3	�zk�����|bS�5նK��v)[��!e$C�D��Ғ�p�Fo����W&<U9�lv��
HP�17 @H����xAR�3��l>�@��\c�z\C�&&���d�8�δlT�#�������L>R���P1_��~<��X�w\f/�"dP b�93{ ����w�m�����R�T�W���Y��&D��"�}e#O��������YS��AH�<ۊ��_Ɩ�2������O���3��� |�N��A��S��Ej���Wa�_	8F�B��Ϩ!���;���>�{VU��h�hd�`�jE�YV|�4{A˃���FZ�F1�"?'���{:���5*T��E������V�h����7 }��J����2u<Pq�d%˛��-Ϩr@�˜<Ab-�/������4�1�~(�v:A�2��{a3	��8ۜ���r�n�?,)��k����|6�3��mW���sbȜ���X�M��k)�������,x���e�a��a+% Y<$_{�W�N�P=
���9gg�������VEq3�i�By�ƶ�o]��ͤO�E��C:��xv�%��C��{��l�X�z�[����(;[�P�9��1L]S��:&�f�����ݯ�"g�I �����X){fG���ws�pO�{N3Y�c@`}��S�ak�)FQ�GO�]�(3��%j	d��+��`�kP��H���M�]��?�6e!ո��`�0��D��}�������+�B�8u&`l�+f�?ү+�s���;%U����'�����ა��L~����9���2<�_$n�U��������!�������U'k	Ͷ)qoJ������������
l	s)e��x7��tCO��x@M�.�~�����ܻ)�_@6jro���f�7�����5і�bdX�����τ	w-���b�XGqn�E���t��;ܣ�a��6��=̉�P;�2L�v���Wי��K����A��MB���q���ʧ�ǰ�r���K<����u��b�Q�+}����ir��s���]��;{�GB�l���Q�(G�$I�:�4�q`�i(��:��^s�\���IF���T~�jC��x\ep�吏��H`���+U����RCJ����c��5�b�S�a����'�o� [ob��}�k�A|I!�AS��cu��6	��L-9!��C���Iw,�Yu^��6ph"nW6g���l-��F��"���^��S�J�+�G	c�lŶ{x�v�\�n��CDJ!�q��;���� �ʥ8��%Vs�~�gO��1z�rħ�@�j�/,��K��b���\W���K-6���5py� ;>M��j��΀�ő�o��f'���B��L�O�R7ѡ�ou�c'ȃ	��?�O�	`/9*$DeUR�5O���:� lzC罂���s����uн��ƀ����<�\��#�n�Bz�U�4���zo6�%H�Gt���`I� �t�<��
 ��/
l=��v�ΐW<$�4ŀ�掐��t��v����90M�#�`���\c�˕�������֥ðVږ�5�R�8���{�׃�����L���Ƚt�=��h����'/a���n��[dm��3���<�W%
�G86�4L�'�Y���y
�)���nn�*Y�YE6;���+�mUۑݮ�$w���x%ԏS�=�^3�e��#��Z�≖�[�E��Mc�����>�2ryz�|�{��sY�;pQz�s~�lF4���# 1��ϠO��_��i
���>�x;��gq���7��=��T�6i2��an]����;��Rs;���c���������Scx81g0�)�1K� �Hw�bkW	��)����_Y�A?I��>P�?���C���ѷ���
Ld�F�y��6���K�Uc���G���n��+	L�irB�#l<���҂��P��0xC�)<7[��|w��oq(ُ�œMu������,�������)�'��g�#?�s�ݔe�u9�E������8@����M��k{ε򽊌ls���W�e�\���o��dA � e��?�M��?��wg���
p�nh�a:[�/2L���]&� p٤l$c��xЉ�-�M��J9�yGܦ�?:b-Vy��$�/Ld7�vG^��\�,�ؖ���8��%�s.��J7?BU��q�����}���j�^�bp5w��HE�yD���:%c�*xQ�!׺�g�~�QQ:֥ridi��Aÿ��e�b
�4�_���vr�~O�����u�qُj��m3�U驛s���� B'�-� ����*���i/��a��-��bcV����3A0m��Ѿ��� y�������tk6w������M4@��w��B]J�~"�-9�wK�X�����0���4���JcֱHA<��9i�5[J�n.}$�?����� t�o�Q�Q$9��f�`o\IO"�Y�"%`������EV� ��E~#K��[Tf��܅иx���;�XQ����3�M��� ����ˏw��G��)�oZ��j}8r�!'�C��/���d�͏t�h��.�E��_���	�3
�ە
EȨD磻��Z�b��m`�����m�ސ+��������Jg��0H�0��9�}�~���5]?�|�ϴUw�����Sq�[�XͿ�$C���m�������|���{$�ɒ_����h�b������r��|��� ?=Ԥ���yق*l�kA�f�S5h��_OC�t�����E�ҍ�%
�s���2$E0$Xt9T�]�m�󡿐��Xɻ%�b��&�Js"sy�y��Y���躱��D嘜���&�����{O�_Hy'
 z6
q�"t�e@����ƻ[�����0=�,;�gsDy�\q(d(��f�;V"T�Q�o��"ͧ%M����LY��͝W�G`0���]����ʝR�.,�.�=���[a���1a��3Pğ+b��si0SQ1�BI i�k�4�>֜�<�.)�L�ǡ��z�a)v��<D�p���_�֙�\^58dׯ�d*���f�Y�H��3�u�k��Ͷ���w�ܐK'Ks��)v@8!�zC�pIN�L�-Z���e�(j�W�l9��f�t�H+d�7[��[�Dsn���#Lv>�-�ו�o��C��:�W�3���K�#��I�)�ǻ��������&Ne���w�?/K�ckEO��� f���J�m�T���C�uk���W�gK�om����� �} �!���/�T%��ݴ�=�ѷ9\�k]�ѲՂ'0���=�ON���N�l�|�����x�E6�RP8_d������yD�����mZ��z�U���h���dM������t ���<�^�M�Q�Z0���s'�2r�6������TL���!�48f%ĕ�+�7[Qb������]�u�%��?������-j��@���<��-��xΉ�A'���I�YX�vul�2Aca.��������]��/�,�)�F��ⲁ�κAmRn�Z�b�x̞�RMg6�kꮽ���+M�s�B󌙃4�aFc@Y�%�{\��NӜk
ZZ�9b���B&�BH�qN��܀��eo����?�$Eޯ��`W�:eL`v)�`%�eC�y�{�����V��Q�u[VX9��1�?@Sg��&9z��z�9�|[���TgԔ&I�r�kG�XXGVaS��7Ir���oBuO��NN�<�޸�X�S �I��0 �BR�ĸ�<3�}�8�r	߼+z�������T����ɇ�ّ?nj!�cn���0oi�v}9O������=$�@��&{�զZ\�[q+׍��3�6ā�'n��;��c���4������!��BL�-��_xa���.یS�^���C�U�l2ͱ^�o���:�P���g�vJ��D8�e~��x2�t�N��3+��I=��&@~۷𿮚�jG왁1Z7N*��ѱ��d�R��\�Ͽ�Q-S(�]�WG��<F���0��NWۣ����q�=g7}P6-�L���㹙� ��Vv���삆 ��BN�^q�+#%S�k�����<[G%��Uŧ�U��}���~orFg4�1s�].�{�ӱ���&X@t(BT�$�����7q{F�i�o$�,^������IA-����%������}�j�%�}�݌ٴU�d��1�PJX�:�~G�5@�Sv���i�P� V���2 XkY=I �hA�÷cP�)6D<��Ƕ!��t��.�w�e�Y��^삩h���Wq�޵5�<-�?�p�x"r�i^�E�	�+aՋc+�@�Q���qh�ɐoC˲F!ͷ��;�3�Tk�@�� �T���rO��1���"G1@�NQ/g*`��"�]����B���m60����T 	;y�g�Z�Ѱ��ެhI�E����eݰ�5F��ᢡnќKo�j�'�	��C����;e�)e����0��PҽE=� ݽ�;f�Ng�Ϫ�uk�-��Ƹ�������>Qɽ�u�0֩�5��z
o� YxG�(�\�����tzS	���*�j�l=`ċ��>W]�����-���h�QB�,��M�Wf`�P\����P�	��"Ë����SR{�ȁ�e��ƹ�>�,��FL2��Ș[r�xע)r����/��+�);|�v��m;8�\I�Ò�,%�L@81�4uS���B���%y�����n�iZ*���Y@	\���f�(�|���$�k��SǏ�����}�eܖ�#�Zk�>��{E-hco� �n��'�u*�4��{|+�Y�FQ�t	sY��Fo��uD�1���������i%���X�x�_g��6���=���ߑ��2�4snx��M��;�;�sv����R���w��dS��1���)m��K�_�=b�����	�u��Ѵ_N�AZ�,ԉP�Pᄺ?�)��_���
�vF�C�t��VK�ѭ7�{� ϼ�%�+��O	g���r�#G|��ϲ���+n�A߂7!�ﶬa�i(�z� �Ru��7���j���>�`���a�ͤ�5���r#z�x)�p����zs��S�_�t���ɬ{��NƊ'P���]VWpū �^����A�� ��5�@M�9���� g����6����J�
�0�D�]�p�pԑ)l�R�3蕹H�ܱ=��T�k�ּ�b�z�����/���1�w�(��\)j��q҃�s)�%�ҝ��L?�7`�,4<��ܹ}�ڛEP�ӝ�x5�H@��Df�j��ݨ�EHN���Q�� ~���:q@i_�&�y��Kʡ}Ņ4~�\dz��������u��4��j�bĦ��GUd(s�+��;�skil ���U�����iJ0�a<�݃��	V�"�zA+��,x��m�y�p����OZ�w�TՏ�sM/�-���WB�'~= -�0�K��.��G��.��/Q�KZjc���AW�y9��[%�.��ھ���)�{��o��Q?v��G�`JL�O]�ޭ�UD%[c	�yz���sV�H�qs#&>k[�\�4�2г�Z�JC�;k�|l��5y3Г�!;��M��ҴUGɨF)�m��,8M�'�$���g����)�(v��#D�.���kl`����3E�&��Cv�?��Q�M���4��K���%��M��d*�ɾ�g1#�!�*�(�]X�� ]��R���w�a#ʵ�d���Ӻ�����7=m�]��/�|`MH�67ɭ������=���A�r5�f���?����DPٝ��l@�T�j��׎P5b�(�O���O���`��C���N(��ȋBE��Xo͘Tw���(v¡�暙�2� B����J5y�ػ��ώ��"�ED`������f�4�$�Zr�'ei�z񞣶=�e��ǃ�sG��Ep(��02,����"��y�mq�^\���af%�r"��Q�/��}�w������������������l�7]��g�3��R�d�"=;�K[<;F�l�G��5������Rs$�QL�YI{D�k��>S|s��)�)�m���:��aD9B��j^p��"_�d��45
$��
Q*M{�fd��3��kJH��Q�u�r�
���WK.(9)���![eCy�C�T�����*���+GW��f9�T����~H[U7����(n�b���3{�>���R�J�uC0�c��U�.�ܴ"cs#@��ރ��BY3\-�����=Fٽ��w��/����/�j A��,>umG���������������-��ik�}����jS�a��Y���2Xt�2�9�Fj�����`��ف�O�hx��2rB|w�e���Ɍ�E�ѷ�M_�_��񲒕�k���ԁ�wF��BUL�h���d���{�g����*��9��Z{�Z�	~��K$'Hw7��`���T�)��΅W�oH-`�ɛ�7��g�d�4��u2��-�*�-�@�!<�vn��^"�����*.�4�jv���2��"a)�a��E*�s]�����,���!|̗	A�i��mM?���Bb>tr�'�M��k�TL�G�ճn�N�m�׺aa��Y2G�{7ٽN	N
�M9]�םl��YIqiE����|�o�f9����E��'�ȝ: �+vD0�%�A�Cx }{%�[ݎYF�Q���A�[��9�-�1BB�SB6Y&tU���Du�T��g�G�I6���X�T�G����S�Hm���4�
�Ni���YQ�3(�S;�|�_;��=�C�۰3SF�S�c	Z�+UWC��J��>����B�"?)�-!/_�V0JgTWY�}�/����ᰥ���0&��B�!�~���+Y�}�8��1�꜂2��X����y�p���Wk��o�>�(0_����U���-�� ��]��$�U]��ͬ�o ����}���_���aW��K��eyNx-��t�m>��5��d�����ےE��� $j�>��|�7�Wu�t�Z�� )dNC"�7�a��߀-�&�XB2G'9���fP�iT�ɒƣ��"۬�=&P1��Lx�(�H� ��#����z��BT�[��B�1�q�wh��&H_����<�ָ�V���6���}�bVu5r)��Ll�]��g{n�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��~ ��UWP�Hh1�H�f�rl`�9�-Y�s��\����V�N�/zrzl��a��Bغ!#�ra�@B�zZ���^����1B�䜧��1Tt�2�dR��>����{�� �Z�(�#	 �X�i*��*Z�~����AϨ�.�R��%���W]��i!���Qb�;��F���C�MDN�	�/u�1Aɍ�'PgP�� �|z>C4A9ȿ�Y��XT���!�^9�P~�[uK���؊A8�[�{���Ө�^:��$���n�� N�y��x�\��#g"��g�y�"[�>�k%�3��'d� h�I|�Ԉk2���8���U��9���q�t�qumJ^W���%����! Խ���z"mID�L���ģ^s�?C�^*p�a<��f>�Gd�Y!J�e0d�?�������Ƌ`����iJ/��~��j�S�΅�k�J_F�W�8$V�!!_{z��&�w#w��$�ާ�9�l��!�=f_�Sd±_���~9u�+���l�w���}�Ew��k4C�"�'^I�9<�Y~�Џ�P����\��9��&���س.}��٘ o2��5�����e���$�l��(.N�� -|zE�^²�_�5+�z�q[D���v��	�濛���y�W��*Hh0uz��F�ܢ��$�+̓
Ԍ33�	��a�̝c���/X|���B�,by��Ծɔy�^&f�X�E�=9.^7�h#��߻�(;0s����5o,{/|�|_�.J�����@Q�p_�����)��0{�v +bG�����&_�U3j���!��4n�@'-�5�y[���ä��UV�F$�'N�&���/�bO�vD�e��G%	C�)Tj�έ*<܍V]F�0/+�p4���vA��D+	� j�cm�<��+����8���M�	���L	�N�����bzZB�<�ȝ��ǳ@�ݣ�{�|Ϩ^5�Ǚ�������͈���h٪�5b,����(U�"W�𛲭c\����dJi)%+u�ҽ3�T�����ة���Z�����J�7N�݊\���@������\�d������b((M��q-<�2�"��m�IU~�6Zom/��$6�_�W<q���=�CCP�|¾�K�`�L��i��N����ܮ�/�^�X�]�kK�D���2%�M��\g�>%����6=�����U�Ѯ��Emv�}V�LK���+�̛BPY񣎩�E8PV��;��h.ۇ�¶�#HeQ|��P(���W����+}�wd�@���q�ժ�BaL��� 
q���}Y�,B���Op��N��W%*3زˠ
'��o;�������d�SŅ /xW*��\x�ҩ����:n1�[��3Wd�i	#!���k��D�оk�U+�1Ev[�&���LW�g5��꾖�j�q��������1�`qx�����]àS��=�sf�&ӑzQC�=w
����	vKfrr�S�K��&7?�y�7�������f4�@!rbY�׳⬄�_#A%q̠�k���S�v��I2P���pkZf6p�Jz�q� �^�[�=���&&���ͦ�����ލG�k�_%�(Gsft"�W&��s��8o�W����/�!�|�sr����5#ŞP��|�M�>���t~���x������~ql9��5���Ӑ&Md"$�ˠop��R'�d��/��?��%�Ũ�P74�x�U���'��,���y�m0����~�� �'4R<Gٛ#'�r�ѥ1@��l=�]����F0Z�Ӕ�%R�mT�zF�ܸrɎ�@#s����LV��F�a�Y�v�ykS��Q�`B�n-��앇Ƶ��m�G*�_o�`�}z������Big#taR��zKF�62�M��9��N�zB)B��T�:TE�]�U��O��%J�����!�ᙁ� <�Ui���*K����A �d.d0�P���a�W�i�hv�B�;;��~����CT�uD�3��~�����V�'A��P��[���C�
I�0�b���T�M��+^*`P���u|���fb�A������]�/������-���Q���;WxG���TM~�Jn|[�O�W%zV�o3Q�q�oI�5�)j��r���,<�@�Գ���T
u���^�#����%��/Ņ/��d�"��(��+�5�F^�QC���pW�����N�X��YRsԫ�T�0�HQ�Ѐ@�Voƅi�j�|�¸.�K�4�J��Ʃ� D��%C��<�JP13W��_Vƌ�_�KM�:"���w�S�$���*�l��ٍn_YB&d����a��ltL9F(����l���L��ʢ���qƳS�''Y9��~����ӊ�0�WpA�wƷR���a؄H��H� �]�f�X���]8Melj�$_�}�~>.?k� >J�E�O�	���z�&�[�W���Ӳ��E��GȾ�G�=m�H�q�z$�ߍ�����+�%�ԝ��:�ǲҩ���Dn3X-���bj֩��y��f�1LEKAH.�&�����M��s��}�f��{�M|rC�.�(,D��@"�_�ȗ�	g)�P{i� �')�wA��DU1�q#Z��ʭq}R9y�f��f��U�qU'��:�'��&��z/@���<��4�G�0{��q����<�cR]w>�/|��4q��7�]��	Q_�T��<����E�Ή*��)P���{���K�	�<�N�6m��:�Zsi���Z�8޺�nB{D~�/Ǌ��詑�H����hJ�w5�4��8?��v�����5N߂l���bQ�J��=+&����u���-��3��Å�pdRfO�JB����xK\����1���iv�#�K�����kK��:�](���q� Y2������dI�}�6�T�x������_X�Yq}鵶.vkCab���"K#ILoHr�q���ظ��/��RX��|�C�Kܫ��h����7�\%_16f&�Xv�}����ENGIi릲�~Z�f��%R�4�`��2�����c�1z��TȲ�>��{����c�ܴ=-@���^̽B�oQރ,��2�|c�y\��br����<P`}6,�fAٻ�P^?ق�V��"�`�F*�o������"�f���K���x��Q�O6��}&�aSó=-Y8�1w:�#��R�4�lΨ���d6�V]�R�.-���H�9��t�;Ro�_�u	^��gc!E貪�)xROڙ,�J��frzt{垕��gx�-l�Nڹ�E���بA�����tMP����>���d9-�<��/�pA����;v���8����,J��綳�=��� ��Y�(����\ݍ u��^md,���y�6���(��M�y�H��ƭ�Č�c7���<@w�ޤW�gư���NP��6���4�W4͔��93)p�܊�P��il�%�>��!uŝ`H̩�~+j^���D3E����n�;)M��6�lm��^#�ݧ�� {�9��D���I����6����H�l�g��e��:�1��P��d���@>���ڹ]/Y˞��>���E���"r�ρ@�����YA]�	�")��/��.5��7�̸��i��r�O�)l�5���[�D
w�e5� 7��B<e���h����7f�x��D��w�7~e֐k۵����k����3:�V��:���\bAki��l쨋��wу�����Ͼ&q��$l�5��HpB�C=�ŀ��W�Ty�� ���,,~��	�⭺R{��3����������	�)$���| nRKt그Z1d+�"����@�tK�dm��v���|�0��Ey�f�:���YQ���>����]��5�g�Ly�Un�
r1K��%���VS��	TcK<��vC��l7�x`{$b��S#��ؐ"I��3db�-��n�5`y���,�~rQ8�~��85-e��s7�'����4���݈�ڣ�6�Jg�̐oJk6Y�5^F>�+�Y�����\�>!����ܟ�0ӓ��_ԅ~(�n�^qϺ���-��&�]γ�A`2
T޻��~���fn�}kS��Ӏ������Ȓٯi�h����K@O���]��Z�ܕ�O�İJ�x@�픬LZ�e����*"�^%8�R?hZ��hg�?fb��o��.��"��L����4f�Ӓ��|(*����o���tx�d��� ��tI�4�
h11|�Ղ!����cX���b]pjt����G܃�K�œ0��<~:](�/M�24���������	�1���y<����B��Z�V�=���� 9K	9��N]4��b�\Z$�o��6�),�(b{u����jX�����#������h;e�53���g�J����r=�=:����=��Sa+J�m+WP,�U��z�|�i�t�A�rW��JSB^���\H�����={�ԝ旆��\��K�a(/�qOy�2  ٤?{$I7@�6|m�i���DR_�:�q�6����C�� f�K�`�L`����߂��,���/&�VX'o����K�F]�Yy���ʓ\I��%�̸f���X�)^}K��*YIZA��ޒR��K�%�5��
G���N����/���E�������F6�c��mjC-���/*3��Q�D�?�M�lZٚ�Wٱ;����N}'��fRp�ǁ׃��>*Rvj��f*��mq���qf���K��sx������qa���N�8�lGK0��׍����$v�lf�I"R`�1��p�"���G2��`�MRu�_{0^^M�g4Ĳ裧:���.,�����Ct���}�gI��ly�^�b���v�A�t!%qXt������U���M)Z/ꯧAI$Ɇt
�am��?�Wc�+������H����P(f�?�n8�q��ߞmA,J:��ʩ�6@2(���M4+U�����M�լ�ch�����3�O�Ǣ'��a�D��"�Pr��՟���X�>3��u�]�y]��҃��/[�!��`��<��h�j��������]n���M��6����c��.S��{@�L��yb��և��	�6-�׷H٣gEД�-�1�A��!�Ur��Q�K��!>]��؞n��[�S�� �"CAe�>���%���A�]+��"�Z/:�
.�/�7�R��
��wO�R��9o��>�D�>*e�nz7���<Vyd�yʹ��he�\����D=t+��X��a���������
�c�kV	9'㏀�b�f��yk��7���E�=�S �/cv�d���8?���Qp3ă=�p��
e�ť,)AW�z]f�i*���=��mR���3����8�ǊT��A�v��rǟh� _�R\!����d|ro�)���1���v�5〤즕�ܪ0�ڛyB]�:tb��(�Q��>��������g��0yIx�{rKO�zʞ�ES���T U�$lG�M-)�7��`��{��S��"؁uv�Ld���-;<n� �`
���Y"���(Q
ɽ��M�i�-���~�g���$�>Y4Z���}�R�GV�B|_��*k�[0��5�X���>Y�(՘!�ᏝȢn��\����9T�t���o�Jn������~�S&^Eǳ~v2�ۮ�\y`��xnǳ�S����)�T���#�Fi%����@@&B�M̋}e�@U��5Z^�	U�Ev�Z_eŹ���"ºJ_����Zg�Z+f�o�s���"�X��
�'4�1��=C|����שoXHti���� �6@IM7
�}�|��!�v�&����8���(7�EOI$mc��n�k��G��#v2�$�9����8������&0�����2�#���nvyu�jn4������>Xk0yM�U�Y��H�q!���p�k��� �U�#���a�W��׌�"X
P��n��B3*���6;�Մ�����v��͏�Ó)�|�h��&�z��r�v�:ĵ���fvG�U���>b
���U�9k5�r/ۃ-DD�e����Ӊ�>^;F#)P���o9y����}9��>��iIo�
��̃Ie�#P���\�X�&�nP�*��L�M�R�9���Z�fe�cj*�:�7��\6!i?�hc�x���E W�W!�{�X��L���m�	�?;�rD�w��ʒ�Ђ������6TLҍ����Xo���.��m0K���r^�'�B�j�l���(l�����Q�Y�������S� 
bm�, "��|�xu5E�>��g��<�� ���%����kv4�C9Z�F2;����l��J���t�0Ղ���(W.0ZUpa�؇l��H+�޴Ǚ�ՠ/�Ԛ׬lR��]��8�f�%]B�^��٬Y�F�m�%��\���o��5��#�G�wS�=Ҍ�S[b��\�Ϝ�8b�Y�� �]�?��h�2s	���[+�J��c��1�Ql�w5���v_�ghgΐ�W����)�Y�2C�0��+�}5�mc������L2�R��ܛ�p�B'�S��l�hsm-�WX=�`�#���9aa�?��w�颜��MQ�*�wH{��}���pvԦG�E�D�.Z>���/V:���;��Ė��v�S�[�!i�A{S�ط8�(�%q%[���6@H�q?��������?�A� ЖY_�s�BbN>f��ܣ*Ԓ�<J����b��~o��n�'"w2G=�c��*�M도jM<r����R�V���	�?wW�a|I���aԔ�Q�U�}dӄ8kk)L/�-?��5���/F?i!Q�z�ܜ�#�^̢��+��e,�&�˫,�J������Ce8������b+��>h}B6<�Yt���F�@�86�G] n9�gT-)ǵM���s��5d����f�<�	�=��3�3`�׺��@A��a��_CBr����IfV��@���_?1�Q�p$]��'�z����J�����~�Q�]4fpF�RS�Fƹ4o��β�
3
�hR�>�u���2F�+kn0X,bw|�&�A�C9��6��k,������m����V~%�E� ��%2���}^��jT5۬>�ma�2�T�?4�>"�-G����0dS�ba�_��O�i��w�T���u2
G��#L���;���p;!����~TW�z�DG��?VŢ�®6m��p�!��f1 ��Ljr^�)�g�6�I����ړ��%��k��g���m�b��� "��^M���)e�+q������ -i���q��vb^q�C�b�β횬i�����vM^��"�0?��b>OP��Rt"<kהH��U1�nqd�c��?��a�@p)���-J�鼎)7ai�N��q-�>%�4�w.�f����[�K��j�c/�dl�6e���h�(׮G"^sp�H�W�fcR|i�c��:��t��y=!��~+@�p��~�E�NT��a:�����&��` =��77�.s��;��������ʉ��/�Xd�痵{Ii�$���E,��&CWOif �����w��F��$6i����y��}���~�I�ߏ�n�/w6F�U�h��B类�
�F~9�cl���T�t�L
��z�y�S�C��P�n&m��O殥��a�=��q��j-;��@u2�C�ۥ��hj1
w�v&vo"k��� ��`2E����?D�+����`í7�7F�^��)ѥ�/ư�Y���E��M^�1���K$���#�LlG�:�Y����	+hz�ӛK3�<�4�)E���L��Aa��]�@A�᏾�3�ʸNY���4D�?\�N�߆@�N�eN�P�v�'1�����8�{ΰ��A�қՏ�q�P�r����@h
�d�p)"���_��kK~�������_"�_�[9���xF2��P�߂K(��Ԩ��v ��U$e��$N�ܖ���z������0�؛mEΜP�N�Ǵ3�F`����&�\=�I�El�vw  M�'�LS�P�&u��ζ�r��"@M�z��:0�g�����I���ru��:v�#G��bF(�8OlP�غ�tg����#��@s�\��}��]O�;Tz��<�L�6_)N,��G\��T[_��q��Zh ����4_)Eqn�B�����z�i.����%��Mě]gF�ly��k{~$$��P��أ��LU�
��/�VU�]�v�5�k�Y���Vj�[�K.%݁u������04���)�}�?8�:j����|]�se��:��,���uH�<�O	0�H�q��0jR���3��i��V�=�5i���$��Z��֯�kc���8��k�{~l�JV�K���0�; OV��x[V$�~�ki���$�3o}|*�E|����>7x�J�#N�
�8i�+"�B�=�N�E��
{��8ZZ�u�O`�ŬrҒ��7�c�RP��/�,8�M	�*L��$ӳ�q�TS�g�3��N���~�,�N�sG �I\��P�>��
�-y>".���CJ����r��^؆ڲk.k��W�����F���Aprӊ��X�=b%O!p��9�)����46�!�r�{_����:F�4��ۭ��r�����,~�7�� �:~ȭ�H5_L��'p�`�&�Ud�%fz�ه��f�v���a�%�"�?z�R��9�0�&l���*��"YO�مaU�l���3�ݗ�q	;s�<���}ј�>^� uL�{��H�h�Eŉ;����墍���L����?V�hEH��m����u U9��j��|���pU�/�?�疌����h�Q�]pr��١W:D����S��;�/����n@��O�A�;x�X��ɣV|����	�+�L=��<�m4��V�հ�������}Ww-�����oi���m��&V�-;��h�p����,Q�h�L�(�,y���d��|x}�B^���.��8���AB_fD��G
��� ��}W��BJ��O��N8ZW#bw�pl
��oIZ��~����do_�>�IW(ܬ\6�@�]��x�i1р}���5d1j 	a&��߭��߾�֫�/1P;v���������p�x��ӣ�F,��B{�_wY��^��8��f�s�7]AH��$��q�-&����y|=���ML	4�Kr�%�S�@J�$Խ�ĵp���M���u�d @߉�r�<���5u���#�?��f��چ�Q�
Č`^���P	}y�nDZ$/p�Ȋ�q�@�^��=A֟&��p��������Kjk#t���ks��t���&^Q|u8m$�Wz�ŀ |L!�X�sp�����pڄH�M�q=���q�����VKq*�+ڳ�����Mbs=�<���1���'p�����ڋ>6?
m��4��ўF4>��U��'���,S2hy�4�	�>|A���� 4� F��w��p����|�@����6�F�du�)�R�c�x@��v�M�k�.s�\��Jo����ף���{��i2` �w-h>�ӆt������T���&uz� �ِZB��q#����6z	�r������7�`u�B�������TC���2��][�ctϏ�w锉��k� z��i��*	t�GldA>R�.b�����
�WLgi��P� #b;r�l��wCRVCD}}��>��� ����u'��P�?��!<C�����_�#�T��0��^���P�"u�Ny�dLiAg�������->V��`﫡�2��C^x�/�2�=�m�HE�[��A�%Pؠ�mY��/��I���Zv��g�����/m�py�Ømu���^f_=�����BR����A/�"��3������^���CѠ�pU�-�i�_��2Y��|���E0M���N�׼��L�gϽ�:������F
~J~y��}*�YP�B�c���J>�W3&�V�"_�Q��]z.��w�v$�{q���l<�ō���_W-dFɱn����9D�p��V�l��)WqV����ݚ��1C�'M=9G	~u�*�ZA��U�ڭ!�5����C�؂��C͸ �����x�V��We�$�'�|A_.��O �uEC��H�drz!��[3Q��"~�*���y��;ݷH��z��c��[͌��>+{D�����x�Zǰ`������s~Xk�¡��b(��M�=y��f��0E	m�.m4�����t���is0�>��{~�$|0M�.Yj��@ �,_��3���y))i�{g� ZO�� ��QU�I�/���;w쭯�sX�y�,R��mÓ�2U%��Ӯ�'���&=vl/dѰ�D�tP�G�<��d��}�\<k�]�8�/z��4����q`��v�	OpI��<�0��/�d·�����ӑ���	�k�N�E��O!�Z��<���k���{��4�-c��H��l<�]���wIh�p5q9Q��;�����}�*�K��jI�� K�Jx�|+d���G�]�0�i��V[�n<�$',J��ܯ�7e\�W���#��*���a*���ퟜ)��L(<�q��h2m��,�yI�	�6�h�6R��3�_��q{�����C��0�-m�K!9jL-����v����/s�XX�F���-K���&��\�\V?V%]P�f丆X�L�}�:��C��I'f�Kd���J�%P��W=����5���/׀)��{���n��s�c��Z�(-~J�\v� ��Q\�8�L%�����7��D����i�:k}��Cf���ǎ�ـ6a�c����R*�(��w���'fc9LK���x�C
������aVϺ�;1@8��>�����Í2��fO�Y�[�7�R�P߱�6?�0��T���
R�B_h�X^�?�gaa �p������,�Y��$a�t��Օ
��gv 0lFl(�o���]�A�=wrOgt˴|=�<9G�"5�κ� /�S)A�I���`N�C�v"2��L����F��#�������(SfNɚ�#�����m��,WX1�w�26Y�(�7:M��y�F�p�C��B�9cu}�:�X���mǏC����VP?=�B�	畏?����3�b���4���+����!�Nm`����_j�w��K��!!�n�k�M��6&����u��ۦ��S�7{-���Bʭ��8=�p��6�V��qHÉhg�����1O�҃N0X"�Vվ����Y]-�e��v �H�Z�]˫"p]�����e?��']�bD"��/'��.s7|7Lٸ}+�M�O��3����D���es��7��~<#J���R��$���6��D*x��u�b֎O���������1�1VV�g�|!,b%&����f��]�-�z� �9�|��Q-E�s4���9�p �$=j݅�_��Rhy�Ϯ�g8�j�3�	n頫�R�ER3b���;�����.N3�g���F ,�R��z���d)�<L�w���O��b�Q��0��In30�y��:�
���yQ:w�>��"N��M��g�˞y����ȸK<�P�+��S�vT��N�iU����5 7׿�`��
]oS!u��NvM��f�d��-��nп�`�0��欛�p�Q�F;��Gz�v��-c�k��S�������<~���J꣺��LO^�̎N�k���״@5��_<�����Y�U�.�~�<+��B�I��n����~�<��n����?��+�N&���k�2Hv���e���sQn4_�SŢ��!ʟ�/��J�i�񻲁Z@���̘S����=ւ���N��Ҋ.Z�ƹ}Q�"p�}W�:�P��Zf�Sg�.�f�Ԩo莙����"[x�|4d���P��|�t:�Xf�o���t6�`� �C6I���
&z| ��!ە�c횲y�3,�7�TI�x���(�ԫ%#�L�$�=��Grv�E=�XG���0�\рx�#����;S�u�4��b�K>���0f2�U/���u��!�k�S�k��K�����p*���S��O=׹r�X�&t��x$�O񫜩A�;CKn����s��>[+� �)J9h�`ر'��r ��'�@�'�HvtM+Ui�
>�;��ڣ��J������Q���,�3��׶>�B�#6�]PVF�o�������9e�t�%�5����w���5eH��7]��E{׽�@�*φm�5�����g0e{�j*령7��6�N�?�GF�E���7W��$_){��)VL���m!t*?ho�Ds�*�7HЏ�����J��L����L�ޅ����O���#A�l�x^��I�j=Q��%�����>��pF����þoנk� �a��!����x�-,ESx"�͝:�:�� �� %8Y���#�NZj6�;�`}͸�T�՞����p����($�Z�|X�r`l��4x�E����-g��s�9�����28���ҕ�B�O���pY���F5%V��V'o���a��ƔB�S�����[�J\]��"���f}� �P�?+9�h΄�	~{�[Xb�f
p��}7l��5c�v�0�hT����:�чYYwV K�85f��/���p\RV`�FA�r}r�ݢ�'�[����s�l�D*�=��<wpWaΎ � =��Of�/�.>�3�̜��r��t� vA���R`g���~.�wS�蒈:f��hw��c��v�d�[�`?���%����q�X���(HU>Z����ٝ���ގ��Ѓ��� $Cb{�m�M�*A�I5��� b��o���nV�Fw_���0*i�����</�l��Ce`��juw�4N|"�A�w���Q=�ʎS�%��)� Zbo���ޜ��?Y�Q��)�*#�oI�";�+��j,����8kr�W/��@��*�8͢��VYZ+K�а���}��<�� >]F�a8#�]��ʔ)��֒T��sɵ����4��)�;���+�`�`_Ty�dW���������C����e��x��mW�,911%�p1�d����zԚ@�|l�Ye~+��]� Fh��Smo�ᎈ�Ȓ���
Of�k����ߟF�N�+x��X�ޠwj�2��ZAk���AB�܂� ����ˬmSf�����2�ŉ<�2�k�JL`���?۹�Gm�m2�`?!��>��:G�wl�����%�_�<�z�S�!�IT��Ou��QG�i�L����x<��5!h���N�8TD�u��(�l���oW���k��<�!�Sf~#n��r���F�v����n�v�ߴ�.�ܩ�Dg��Y{����M,��ox��x\������-�5F���pR�b��C���{���c���	�^���0)�b���TBt��R$�(��6��o���8��N<��@"�*���^J9	>�{�*a��wN�<-N�EO��wh����
�Pv_[�f��c.��d�;��.��` (���GoL�p� ��o�c�:�n�����KtN>=�4�~x+�p�~�Ң8�#ah��.�p��ъ=Y���`��%@������//ӆ!ܔ�{�N�$�G_E��P�$�lio�������RĲ���$#��Ɋ�?�?����*�~j�[ߜ���Q�6�`��U��Bt���7����~�j�cy���į����
�GyH>L�p~�P������\y�3:p��� ��#�jZ�J�-2��+�����Bj~��w�sv��K�� y��2����tD�:��xh��Нs�Ĵ�s���B��^�	�Ypjf^<�:8�1��)�T#�Z���TRG�P�YW�z�E��+U�d�`�x3�"m4�����Y�x��[4(D@�T��P�3���������D%>c	)�N��@���e�V�ңXX1�AٚE��{���d0^���^�uޠ}���W�h׳$�ݥ������o��K�y��o�CQd��e��,t�9& xS����I肘����0b��l���[ؒn*������"�,ޫ��  �?�0x$y��z:���K@hQĦh>��CX/.�@�gZ�y�2����K�>ʵ�tS���T�|
ێ��>�/x��7�X?`C� �`S����X�I��5@d*ļ-�o+n�¡`A��p�����Q�A�F�O� GP--���������UEQŽ�T�~��̓����Xlyk��!m�5&n"���G	Ygg���({�f��Ń��s'��B�kȜ�F��nR�ς����'b&����� V2���S�g���en~�CSO���D]�Z �i�hd�|�@��[���"�����֌f��@���\��ZV�)��E�"�3�����Zp�9g�80f*(�o�S(��&;"Zzˇ�"34.�]�Z�|�(@��MoO�-t@����̺ i6�I�)�
0��|JX!�T�|���_�}�27�I�旎�U��^�/#m��$�ٷ֑�޻�ި�"ߊ�\0���
t�#~l_�EYEuV��4���,�>��$0���U��v�?!��.��u�k1���w��z���.���n�׃3�X� Њ%����uf�sW�;M��/�5-��F �&d)^�h�����;r
"��q����$v>b{Us~]>s�#3Z�����AF�d��[�ދ�����>\]#�;P ��o��?��j9�"�����RQ���A�cb�e��AԷ���ݽ���*�k�$!D��k���FteE�(*��47��6#�]?���O���`��W��J);a��t�L�0�m��?2VrD}y����*����=#�TL�L	N(�5l*�O>��w�$40�?6@M^�����Ihj�Z���٨��ț��� �O��N
ת�� A�ޡC���4�x�+�E�����%�g��D� ��%�6��b5
���Z��s;"��͂����K�-���G8;�vgx(.��Z�o���YlN�]�Ɛ���շ���g��C�����8$с���B�M�5Y*V�F�A�%`P?���o�3��+*ƞ�eSӷ�ң�T[Y��\g	4l����� k܋?5>}h+�	�h["ñ�p���8�ld*�5-�1v��mh�M�n����Y�:)��&��*50���9���jܙj����|��'��'#T����sį��΁=4���oz�JaHk��J�7d�9w��Ս���@��{#�~�v�����, �?1.��Q�2�I:����2���mM�v?r�[1���#�/o��_{ q<D��BLH_����2ԌW��bo�ޘ����Bx���xbEQ^�WN�*�?>Ӎ�M�b|o���n�^�w)a8�:�L*���U�<��v�O�� � )wNw| VQɋ@Bk& Q�ԷF�o)I)c�f$g� ���G�?���QfM�3W#dD���F+|��,��zނt��aI�u�;�'*8AE����+Tٰ�3�}��H<%���F��48m]�]h�^��)����� sS�&۽)�>�Y�s�Z�T')�*8$`i����^R�����^�.C�ȁ���}���7��6�-1o6�p��M�d�z�?��Ʋ=��h�~��?]��F�����1�����%�͋A�N
����5 ���cF6T�+8zX�^�wt�>�A� 쓶���ʂ�jB��-d`mC��p��|���
_2�r�T�J�!Uu�CV(mؕ^2�)?k�%>9�MG� �����) _\�D���+8.T�c�uI<@G�<sL�+ә����{�M!2���X��T��[�<�6Җ�y����}�!a��f��c��ru8
�^m'� v�Y����9��@�s߾�[֬��y���Ǫ���`3Mv�e���բV�O"�-����^�z&�bbC����E瘚-����9��B�}��0g,b���Ǥ<ut���.���+˅݅�G�Z�d������1@��ډo�JC�,����a���N葇-X���4�w�$	��/Y�Z}w[O-ځMc���d�G�+j���(N�nGy��pݒ2nK�cI0b�x����yt�� =��~�vp�Mb�\h�K��a�`�x�M�tL=#R���i��nRյϥF���#�@��/]��^}[{��@$��6E22��?i�H�L4���K����$m����	�P����~���&�
�#�6��kß}�B����J�ɰ~�c�c?���E����&�Tn�yҕ��:ǫP�ݤ�������G�4K�J>���d}j$ ���i2LB��o�pv�j���w��Yv����� �12�ج��U@D�,ん��*�N��=�G��O1�\t!]��Y:�Vh�/��nP1�V�E��d�n�?�G�Y! ��O�c+�љ���I3{=[4�I��c�_��W��>�D@<߬�#Q3���%`��8��D���Nz@4�ee��m�&1��u����{ep�.�����Qߨ�R�*%$���~h�ee�'�=��9��K� ���a���V(��6�s9p��x�?���a������c6��!���y%e��JN;�p��~����Or�@��%G!Y�dpS����NG�034r:`�NH������I�m�@ $4N��ڬ瓬u7�	wĨY�~͑Q:'0:�t	�C^�ㅃAu[k�:�3CG��oF?"�Oc��Я�æ�g&��O�.��Eu\��}�T�O�f�T�{��õ���)�=�LL�\MrJ���n�1u���A!`�Q)|��n���iIz|��$Ra��������]��q��}[�����4I��'hU?@3����
l�m	�R5.��P���jfX�Kª��{.�X��g���Â�tt8��jΡ�Ϟ8�|�rsʡW�H"�C�j�����	�'H.�@�2E6RgH�j�iƶ�V�
5@H��v���m�яM���c=��O��k��5lW��^*�%ӛ0!^�O���x��rġ�k`Q9�p�[��N�|� �E�;3�>�x(v1�:�X
��1i�W���o����E�
��o�0����i�����I*�7�������l�&,8��M -�CH�$��gqJ�#���
��1��k,B�ъ�@�����m����`�����_>y�V���J������Խ&X��u�kń���CF����9��X}�Ӂ�OX��;%��0�ꭈ�������Ur�2��e�:�D��A���r�vl�|�~�f����1~:5�o��CdL/��~������l抇+���p��T?`[a]��"�W��z9�ٳ&8����)O�6ka�~��[��3,�"�A�;j��<�4��4>3��a� ������HQ�H�\�g;���}�ڍ�� L)[���V3�H�2�m����l��9n㽢pwP�g�gq��ږ����
Q��8��H}�pI�}��cY�2~��
SC��f�t)S�e/�&y�Aağ��$�騊Vi��@ǡcР�3�m>V�%շ!9��q��������E�)w���2��q�VH$%;V
�hy{ɇ�n���Q����P�(��������w}j/�U%�&i����BVq���p~
T�"��}�<�B�3�O%εN5g�Wth�GT
\T�o�<8J���;d����U�W�/\�&����u�1H=B�0C�dh 	x��������Ώ�O�_*7b1���vpa_۵��E� ]�~	���d�F��v�﶐��Ϳ������)�J�`]��:j�
��65&�p��=�W����	�#r�toSxff囬^��,��f���ɿ[\�@�Dr�R
׈M��y�#V���U���Ƙ�H��cy8u_P��Ù�*Z{�%���q���^���=_N&[h�����\�ޢ:OkZ���5	s�t���&�ȸ�=�8��W�	Q�7jH!
^sgFK�Xp��ӡ ����M>���U�f��3y�sq9`�j=����M�u��!$u�'�Q�����B�^?�#7�$��(W�4ubPU�e'�D2,*>sy�)���7<�Q��5��4u����g��Ǝ�֍m'�GFE�9�Iz=R�b�o���M��"ǧsw���=��[���<���=۸�`׿�-��j��-�\*q������z����g��B�gS#I�ȵ�8z`�j�˘������.�U�B^���)@1T�k�j���˯�z�����`I��Λ� � ipR�*`���~ �AU��.Y^f������}W�UBig���W�;��ʺ6�CI�DT����bx۷}�'Vr@PV�$���Cz�*��.s��-�T���9�(^?�CPDy�u����[�3A>�)�A�7�Y�9����*����q�E����x�T���"�5��"�[O�Y%g���d���IBk	���]����f�{�)�햺`fusL�^������<.��RJ�x�Z"�7+��\h��K|^9<1Ch Qp�S;���� fY�^.���%0$]��(�+�����ƑA������]� JuV�����UP1�ٷc�1*Je��Wj�V��_��s�����Q]w���$5���?��ls���×�_N�dN�%8}�A�9�_���l��n������q��莲'��9�\�~�I���d��oL<�����򘫈�����k���Q 52g���UM<���e�o$48���d�.T`. ��%EZ}ڲ�N�;pzؐF[�!�.�m��a���$��2��Hn�QzP��b�	�-+Ҥb�Re���lBǧu�̣�"y�9X�㡈�2b��Ԅa�y"�f���E�m.$*䏌�q�7���.��sg��%m{u�|��.'6f�@�O&_�f���)@��{^/l 1x�ͬ����jUy
����ˈr�m��)&���ya|X��.>�*eU���*M'�}�&T�/��|{n�+biG���o��Ԣ"<�#M]���/qd4�݁<JE�2fd	�R��i�<��&�F���~�ƭ����r���):	]ժN��ۆ�Z�)������Ö�xO{�6��S�ǟ����Vđ4�W���thߤ5(g��� D�nY��(�q�a���I�a�����J/ʞ+�l��y����O⏠l�յ�e�F��"Jw>��cj�\5�:�FX�a�m�x�&��V,� ���o�f(ӑ�qs�^2ĝE�c�$I�ֶ6��W�����_-��q�_ܶC�`CJ>�Da}K��L�������T"1�/�)�XK����K�y���\�W�\��%��f;��X�'`}�|]�:A�I�<����;��%�>��t��0P�L"��&�&��3�2(S����j#�c)e�0%-����S	sא�Q�$���4ِ+�����{à�ߏ��1��}��Ufv���%x���������*1le��鴪�f��Kj��x���d^/�2Q�am�#�2��8�\�ooĵvǍ�s�νE#��t��c�R��0�t��Fyu���,��S�R!�_�j%^�HgX1�G_\^�$�,3��{i�t0�j�!�gm�Vl�&�&���c�A�ɾMt1TLK3�z��wP�q�5/���Am1R����en���{b��9��]���zJ�l�_�n��(�NFɱ|�S��'�m:?(,�����~;6���(�fVM؝�=U[;{��̸c����a_���C�ƹ�����ͤP�F���O�,�<�%��3>^�?�����������p!��P`T����js���O,�8��n�YJM�b6��M�f��R�s��{d;�Y|*��-P�GE^6QeR{l�H:"Kg�=%�Q!�1f��E,0�.�uw���:�]��8��W��s�t��"g`���A���˜��]O	�">�x/^�P.�^�7V��Tt��v-O�����.-�p�HD�:e��7�/<�D��
�ȴ2����ҍ��Da&��O�օgV��,������;:�(�V��J�db��\���=�6��;��I��w����(#��i^���3��_�p׻�=!]����A�ɱR�G�������� C-�wwKR���3���\�%���ۗe�~���O� ��R�Փ���d�Z��J��q�fޚ�Y""���^� C�0�w<yf��:�۬82~QQ�<>�Ɲ%v�a1gg�eym"M���Ks���BZ�S�ȳT�@5H��K�%"77.;�`0ǎ
pSŜ�%�-�<��d7l�-_n'�#`.^Å��'�	��Q�|��8r���-ڤ"�"�o��g)��7�~Z)�!]�kb)�N���k%�p�5�Φ3���'Y���'�&ޢZ��B���|��߅�7n��	Ϗ<O�Eb&W���]�2_�ջ��h�zE�n�k@S\FF�B8՟���G�
i#�n���i@�͡Ȱ��/�M�d����3��-&#��H�Z��O�T�"'Bk��ە�؃Z�N�g�L�f��o���O?"ǼT����4�.Aӧ��|��N�or2o|7�t�+�,b v�Iq�
}�/|7jK!*�����q.���7(�pIH2��T�B	���#��$�y.��()�ܥF�χ�3V�0�Biї��#���v�u�^�4���٤�>���0��[UF���l3�!ku}�
Ik>�S�$&���G��gd��gװ$!X�N���<��sŜ :;�����"�i��5�����)�!h������rW�*�^ְ�>��vk
U@��>��ɟ0��]����Q:t�Xq�#�r�w}�>���#�p�PͰ�oݞV�Ơ 9|�]��]O�.:�pT�e�?��}(�|�c���*�[���R�]�}���Ce�,�*B(�7�V�6�X?�#/����Y�W���(ϣ�*L�=Cm8T�?_RIDJ�k��&�X<�Fڡ�L��H��S`�|�0�~Ŧ�>����2^IA��АVjT���D���ަu{�-G�:S���� .���v����\x�$�E
�x��VD�u� ̞�%O�������+�Z!��;/��/���,���������\(���Zyܛ���l���W%��w��D�}���c�.���Z8'��IF@B\lQ��n�Y���F�H�%-=�		o��2�����h�S����0�[�e�\4s��P��Ȏ .?��eh��	���[O�W�=k@�U�lq�5�,�v%�h�<|��*��ȰGYN���T���ϵ�5������6�i�U�v�I��� '0�.ԐH�s/G{7=��rs�G0�a�_!��$���������u�+�����Z�K�&v�2������=C).�J�.Q:}���_�[�:��v��{[>��e�E�|�k�L��qɁ��2�H,���ԙ�R�-{��+�к:�tvbr�$��*��N��0���lbQv o�f�nm�wV
����* j|�(<��	��=��zХ��w{��|����x�Q��m!"4�\��)��WQ������S*�?�ѪQ0���8#��9'c+�4�,�&m��s=��N��"S4�48/��ml*+Bq����	}<�<2�b���F8*�8Z�!]�PWʋ�)k�n�%s`#��ʋ45�`���LU�W�`6W������D���C�#I���C
��d���#�1ܩ�pȹ1�?z+�*���4�~"5]ح�F�����-�XD�r,t�.�
f�1�bnC����F�+�XP�w�Y��+��A�#���Y{���|�:|sm�)�����i6�Š`)2��!���<u�P+%m��26��?Xgu>�&�G�%s��;���-_i;q��^�x��T��Tu��G�%L�S��/�؈%e!������T{!��N�c���F���Z���C!3�f�����R�r�c��	�����������|�������,3��#Ā��@M�'�	��OfW-�L�	-D7����GBb��C�>��	�Pg3��wf�D�����0��/bbs[Ǳ<�tF��{�D��������$��ӵ�i6@�|y�:J��n���uaw"N7-%6�!w��f�3�eΧ�[��W���c%��d��Z5���=1(�G��wpʊK�@�cvט�E#��^��t��B=ELs~�1�p�ⶕ隋x�a�����#����9=�$��B��K�D9�8�aCAʭ&�/jY2��C{�"/$ئ�E��&�-.�B�i&�:�Y_	��p���$Z;�ɡ*�6�0�s9�~!���3����36��Ì��B�,��.����ƺ~]?c��x�=���d�A�y_��g��Pd�zJy���v6��{���MS�7���5�jQ�����G2�3���w7jշw�ػvɬ� P��2i禗�1|DA���ϦO�����wj����A��ɟEjmoY�@3����q�F1��Ȏ��1<���9G,[Y�7����U+��ͪwn�3�cX4�5m��^?��#�ez\��a@)3k�3��3�D��Ⱦ��^D�����Nd��@%Ue�"�Қ��1[o����{r�C�"��?��ߕi޷p0��h�Ȳ��U7�*e��0-K""I���Ch~���p�9ݖ�x�F��tJe�����*!��>����e`ޕN��'��B*�C���W��O�#���v���WN��y3A�`Á*��𨀇�Ix���W �K�p����Zu�6��Vl��Fns���:T>ҙAݏ��a�~�uȺ:&G�WF�ۮO�{`�|Jx0�g3�G�@ ��4~\��}dK�O/�T�mա`KI�ڋ�)r-��8�\����}��:d����9��GmM))*nQ�6��|�z���o.�l�~4���ȐB�iTH���,7�ܓ��_l�U����@�z0��8��y5����}6���j�SeK#+ݥI�d8b�Tko�P�ҷ��8���j;�.ϫ^�|�Z��5������Y��ڍ	T]H;�p�߉bR�"��W�kiSX�V��5���� �C"�~1��S�Tc*����h~k��!l$^_˙v20B0�\NO�ʏxP_Q�Qk�޴�=I�W�0|��E��ۆ��Vxq_���E
0�i^��f�#��E�~
�\�E|#+��i�9Ҷ�7�d��v샹��,%�oM��spl$wWq�lv�ع���ʺ>T3,/S���m�4���J�:y�m���C�c>�g���'J�8���o+Ԋʡ���k�Oј{p��TTe�&���ӮZ�X�%s���=h�5��͹��j�D r ��є�:j������0�'rI3��&~��t�M��L:�T���E�L�)���9������&v�I}f�}�.ي�L�a
/x"9m��v�9LWi&/gZz!��v�O���ay|���h�3�k���U;���<a�f�	k��� ��WH>o"��x;@���J����L6QA;�AV��}H��am0�ڙ��9;o���|��tu�����[A��2�}��u �p��������f��SN��SZ�������A���Q��Ƿ�����-9�𻄎``�m�@�V!��.#[� ��`C���u2R��������V���;c�6h&ӇY]���.�Q^d�Agq(y����a2��u�}�OY�����n+Ռ��B�e��Q�+
�Z��s}{ B��Op�N�FlWGE��K<
�$�o�����@Rd����/BWL��\�i ������1�9�}ՊdU�	�(��զ��� 7�D14�v��7�.��.��:��^��8S3�#��]��ֹB���7^��]e�wu��J2&5���.=Y��ܤ�	��r��S���Hתh#��ٶݶvf
��[-@�)�r�1וNd��G�#���Bl��~Qa�u���0d��!P�����U�Z�d���t�q�o ^��=�=�&� ���E���#�﷘kG�u�9�s3�dt�V�&,����8���W�5�$.�!�OJs����%I��@�^���M�.[�7iɀB"��L[��qΎa�׎i��ƣM�HSCsi��':��a��گ*&?����ѹ%�u�R4b��U��'O6,���y8sи��T���[�4�B��}�uƔ����[��C������_F�VH�6ORw
�ۜ���Ȏ�Js��ϠnP���2����1�[�o�匔`��-����w�۵��"���~��{B��z�'5�4�OB%%#V#ҵ3Bz�{��D��/�`�[�L���B��4�6h�Tg�z�C��|���G�-��;� ϐiـ*�Y��k[A�0�.�s ����.��W��8im���l�;�'ݺ���Cv��D!�Q�b����}G�\�'��PC��ȖC�Q�Ȓ���G|�T���3�^��P16su^Y�∫�A�Ϊ�8��f��Q�s�w�����^�3���Gxn�@�Vf�/�	�lz[j���OP%��b�������KI������
�ݒG��S_������� u@��^��߿�����?'�ޣex"��|���qM^�'Cu�py�&��t����Y4��اR0����r$f�8�������ނ���U���l�J�0��Q��i������RKJ��WW�5V��`_�G��]DR��w��d$��Ì�_l`Q5�P��_{�d�gڱ����N�9hB��Q�5l�������%[�>�5�U��'�F
9/�~~J��`��q�yͫ~�-�Y����ئ! ��*z "���H�Sz/���{e�$A0��^�.��� ���E�K�+W�	zEX[׽4�����\H�Nz}�����_��H;9Nz��@�o,T����+��?�!�a��7��p���gX�ѡ5��b����qQ�y��f��nE���.�H���p��!��{�sTQ��HP�{�m|��%.}b&p@D8_27���C�)�{��� ��6��ی�t�U&2֖�Ӥ�_�j�Sλ%��y.x��8���7��UIhw,a'��L&��^/A��I�p���G�����!�<�$�]YY/���4g~����?	s�0ʶK<�*����Ϋ�٭�'��<?�����	
q�NN���s��ZU���;3���'�bR{&��QL=��\��.ȑ�c��S�h��5�my�������u���NU�0\��n���J��+�>�&6J�X���~z��$@����.J�~��p��\��u��]��N6��]��t���l���,�(���q _Q2���PeIh� 6����!��W��_:K�q�)�����C3���g
KE�-L������^��W>/&X8:�%S�K�.:��kx��L\�OC%�u�f���X�Jv}|�7�g��I�.�o�ƓH��%t��j������߰�S��������G��a�cvX�~��-"����U��b�Q�݃��au�=������h�A�l�q�^�p}�f��2��٤�C�����_�1U+T�3t�F��p�=�Ϸ�t�w	pW�r�kMS>��x�� �]�qX�;�� ��@�r�~]�-��D��#;�.��%��>q�x����K=֌PEr��*�!Z`cf̄F^q!t^��=}��&`�\�G'�Q��އ�~k���2Vms�B�t��&ē�Li�8)�GW�����/!!/�Os,�k����ء�W��M�Q�ϯy�� ۥ-�7>��qfa��o�ŻM��M D�`���3Y'��P���x�Gh�?F���i���?-4�F�U#�'�^�,���y��4�E�C8Ɛ��4����g�, �+v���a��/�rG��F*�����R���4��ܲώ'��s2-����@�B�?w��g�}�`<�-$��ӵH %�Af�虥�ڵRzw�o��Z�B�ڹ#���ˀ�zE�"�PH�Ǥ���ciH?�Bc�����T�(A�Oܜ��5������榔�|��x� �g�i��*ExƜ��AzU�.+�JcD���W���i�0n�<�,;.1��[+�C�D�������\F/T8�';P�$T�'�C?90�*�/�ߩ�T8�~'^$t�P�omu��� �RA���F~�������U�ge�˞~���(x�D���	Ǟ:��T[3^���%�GZ�)���k�IG���#,Ѣ���߭f��g�N[\��u�/�^"QݿPҏс���``���2"S��W�\�/� ^>�DCF�p.D���?��Y���p�0�jh�
�;���-�#��vy.�h)݂iEJ:����FZ?��~� �v�<JJ�W��V@�_�JM�4���u	w/�0$z��$ �l�J0��B_[�d�r�*�{��c9 ���*lB���D��P�,��{B��h'�t9�"~��j=���D�w�G�G��j�-ѹ�>���s ����Cc7��Wv�e�gk$�0N�8r�.9A xT�E@r��v��#zݽ[o��s����a���d�$=x��VH�czUU7�]�_$,+��&��A����}�l�d���~9nX�=����bd��	��yG�f� �EE��.)�-�1��|����.s�
���<`{:�=|lC.(���7@ܥ�_�59�Q6)e{# P ��Lͱڢ�QtU��ʖk�-��������nHy���Й%��0�U��2[�'N�&y!�/�v��᮸�0�GP�2��uM�� r<'>�]�_�/6��4��A�����	}o�N{g<A\��kA��C�T�#]��|��It�	�tgN�eN�I�Z�>���B^�2�.���9{�	i��gPǄ9��X��Y�*�z�hD,]5-���9Z���r����������&Ho�\!�J4sh+�6��������%Î=隗*7�`y�J|x�	t\zP��+4�����ŝ9ܗo䎜e�c�t�(x�q��,2��Ф��I ��6e[�r�{��P�_��wq7���(�,C���itbK�'�Li�t��0�.�(g/�DDX� ���wK���b[�	�\� {%9�f ��XFT#}:����Ic���ꎓ��t%�0ꓹH�l&�q4^�����Nc`�7D�1(�įT�c����-�T�U <UQ#4��Z.���Ϛsi� K�L����}0&)f{$�ʾ��<��S쫚�<*V}Q�VNW�vIf��K�xT�I�N��a�:���`8��Xt;�Zg��x΢���U��
RI���K����ě���?R��1_$�4^�;g,��Tcɢ,U"w�`A�t��ϕFg�g2�Bl�
��+���{�Ac����t���y���"�^O��va�/3��A�
����o
�-���W@V-&{��W�_�~�F�S�u(B
���Z�r��()m?m,���3B�6��[(UM�V~�]��p��/ac���������58�K�*�Ͼ��P{���;��9�jY"3#[����$�B��ϻ�4�8��!���`�*�`AjX�j�~��]d�nicM��;6�݈�����OwY{�S�~�@���'��/,6V�� ��H.�g�����RL1�
߃
��^�^�z���;'I]�4D��.Ӑ�d����",�c�VY�!?Z�A��]��%"#O�/�Yn.�j�7��r����	LOJ*���ԛU��DD]ie�b�7�/u<_���J�Y�Ώ,�r��D�+����J�� ��'��S|)�}�V���8�eb�̕�b�%�3ߞ�P_��oϸ;��� ��WD���p<�K=&��S�����o��#�m�A"�Ŝ0��	�R�k�3B?š����f�����[�Q�� h��R�鱷2w�d僜�Ԣ�3��͋=O�fb������^0*�y�,8:�F��u5Qv��>��3��)	�8g]y�5,�I�K����gc�S���T	'lM��Ťj�7��`�t�DhuS��M؊@�Ax1d�T�-�wnHb`��օ"4����SQ�E��U͛�i�-��X��a%�@KCg������p������J�Hk
u��<Z5�+���9wYٟ$�jo.���Ң�>+�������]��x�9nģE�4y��}&�P�'��2��p�E�d�ߩn�\�SX���~���#���śiH��n��@I�W���Ԅg��E.־W�Ȳ����ZHbl��n",�����	�Z���gI��fܿjo���s�"�L��SCy4 �gӌ,�|b䳝��8oA�}tr<5�� �vI�2*
b�x|�)�!O����|��T���i7�0�I��E�9P��}���#_�#$&\��X����8���<0Tl�ѼS�#pB{�w��u��4=���">�>n0"�aUk3��1��!Ёg��-k���in¬�(Ϡ�� #d�u��X����R_�B�ezH;���1W��E���)�X.T)��h;����-r<�����S�c��v0�bU�Z(>��	���L�����槃��j\>�������>�0#r~*Ps@o©ĘK09�n9�ṒS��3��7�e@!�s�Q�ð�7��*����V3#�b�_ӣ�`e7١*']�7h(G6�	�?�j������e�W4}�J���a�LQ�zm]��?$�|D����ˢ��r��چKL{3M�����A#2��_즖�NN2'(�8^.�O�U�jy���8��W�z&}��R��*��� �94�������hx$�}E��^�D�YK�v Q��%t��T���L4TZ&�;����t���C��ߞ�O�h�(`CZ~&�LSxl@�H�۴p<�i'ŧ����u`?����8������BAI/���CY�U�F�7�%�g�o6�݁����Z�SEۡ�US[KI�\���9��b ]M�?g�bh���	��[]��\��ZRl�
5�;v�@�h�� �f��~Y�$m�Y��ti�5"��kP?G����U�9萮��4'�$�����s�t� :�=�֌�*S��a���<�l��ҪkN9����@OY��]I����v�$׎!���z.�w̻��!:����$^�ğ-v��[������aj>����q��%���H�@}y��>pНT�����P�?���<,b7�u����*�[��8��?�b6%Bo^�Ln�aw�Y�lK�*%0(�͑&<��ۨ��\I��Y}w@T|R���� N��Q��������C)��5N�>���XZ�?W�QX���e��#t_B�^"+n�^,9��ؔÓT(�g�̎�8��xْ��+�����}A�i<�d�%�FB`8���]���P�P)�S���s�(ͪn�pa<�嵎�G��N`�nl� �%�5:դP�BC�e�nE�/P��)���h��1��pm;�V�sz���8H:�Y�{~�]�]=�F$�������G��W�����z
��I�'�Z��m�F��m+��X��3w����UmA�h ���X��o���2��Tm���UQ����2ڢw������I����Cm�n�2�0?�n>��G�"��9����o�_�!6��]A�TN��u�Y�G�ZL�}��4b��-}�!$I��cT ��P�(xCūQ(�_�8�&!S�(f��?�byr'z��P�K�R�Ю���DP�2����bHҖ�+xy���Ӏ��JM�.nX�Ք��Fn:F-2��ӱ����b���CV���7�s�5��D�٦?:��o�D0H�bg�O�V�Ft���`4켝�H�7n�Lu\��{��@^Ҳ�aD�Ju-T�7Sa2�N�#q-�sPwP�Y�xj�Ό�[���3��c�?Qd��_T��D=�(@G�h�pO�� �c;fE誊�ct@��=���~��"p]���:u=��aC�����&�x=����A�9N����cʲ�	/�>�P �{��U$]��E�'����Li(i+�������9ղϷ�$�(G�ơ$�� ����~&�I��׈�J�6���)�B����;I�Oy~bx�c�ᮐ�>Q������k�y�A��,�+P�k�O�ܘI�����]�ؼ���Z��j��Ik�2���g��b)j��Cwc��v8���H\ ���2n�ϗ7��D�� �ੌ��� ,H/#y�"������Y,ǖ�	x����1ˏ3��k��uW�NGс�Y3�����+iͪ�_�3my�4�*����˕�M����p�@����X;33�ƸW,���ݍDag��y�NI�@�oGe�-�_��1�g���9{�r }��$~:�iP��`�糢hVҚ��H���R�+ uKڊ�+A���L�H��h�9��x���������p�}���?�?����eŕ%N�t��9g����]����n���V�K� �N�x�3��`�z�I�[PI�d�_� Vl_�u����u
�V�;x:�����C-L:����S���7"TuM�:�FxGBMGF�ɦOU.V��U$5��g�$A�k��j[\;�}���O��ATu�e�����)�/�~�q\uj�$s�� ��c���Ȧ(�)n��n6,��_�0z����8���B��Û��.��.����"��T�Qy��Ј���U�jB��ݿc��8�{�>5���B����3j�ԃK������I����@�u�ӷf�8 U�j@p��P�2|ƥS�2>ĺ����,:��B��E�	YHQH�'�$J�R��<���ix�V��5r4���kZd��fI�8�nc�I�T�ky�Gl��O��o�%f0�O߽�x�Uv�kR#}���\e|Z�?E��p�qx�u۝�B
�iYi�y��k�a��B�E�y
ϓ���jf��Y'���һ�79�9�&;���,�L�M�>x5��$��q�����!c�~��#�U,�v4�<���2����O�?w$   .    ލp�F˸��%�R(O5f��p"O��Q   �                                  �   �	  �  �     �(  ?2  =  'H  =S  c^  wi  �t  �  Ί  ��  �  y�  Ӱ  ��  �  ��  z�  ��  �  I�  ��  ��  %�  h�  �  E �  t �  F' �- N4 �: �@ G mM �S Z �` Ag �m �w � � Վ � � +� o� s� �  x�y�C˸��%�RhO5d��p��'l��ɶBy��@0�'�F��L��|�t���pd��46b�Z�4?NNqhs��|`I4jE�M�6��"-_�7RN�wk��uGjY�7���
/Y���F�6=b�l��wm�u5�@%=,ĥ�t�X*v�"@�#�0 ��'��O���]37�,����M3����U�̳��A#['�QrDM[Q��=�2�I5'�lÚ8+J��E�Ql�6�\<9I��d�O����O����.~� "G�zʤU ug�%w�����O�RP޺/�pʓ�y������?1e��RfL��篅�t@���ɮ�?������?)����'��$��fe��"�[�AߜXJ��[ !򄟤Y?P�����{ʠ�z��+K�J�"~d�CP��(e2LIcP?���=O9�)�7(X��yr�Є:���1h��(w�HBĭC��?���?���?����?y��?i̟����Q�T����H6&c�hz�'w87����M�ڴQe�I��M�i�6�|���WW&`�sK-n�h��AfىzN��Ї��j�4�rt&��,`�O��f���d-�.���Q0ϕv�Dʃ*��p���I\����҈iB�R�x�4uqNN�I�1�aD�<��2��h{�_�b�u9�1l>$F�\�L�|��� 10C`x���Ȋ�9�"�G{��	����D�ǢյO�t�t!ʌ��=	������oX!VW�=������<��)�?�M>�������`������j0����*U�<B䉵1x@YA���X#N(a��ԃ{/�C䉉"p�]6�ψ���e���0��C�I�_[.}"���̲̲�-�3t��ğ�B$�#����V��Ir��#;��N�F���^	�^T��↸6D�z�@�5���'>a~¥ܯp�xd�5k��9l	 `#3�y"����a咻�xc�&0N�C�I�C�L)�a�Q�Fr��2��FtTB�ɫ�E�P�	�$���J�?����x�����n�˳H�	���d�4���S蟈��d~��K�}�ɋ�l�H=T�0�y�藻g4^x���P�Lɰܪ���,�yRM�P��*�ꉅtİe3�b�*�yrF۲���(bJ�q�4��y$C�c��A".
�jdԂ������VG��(���:D퉲? |��ń�72f�1WV�|��֟H�I]�)�S� �Q�	Z����җグ �B�?e�P#яG�-��)�`��M�B䉬D3ĥp6��30*��9&葭��B��-P���KG��"ОѺ�+N�32�B䉆a~�AX4�T�H
s%�E���OV��>�� ^�Tl��'fR���[�~��S�C��l�8�ʹ]%[�����ͧ<C$����Ie�LK�Y���HH�[��¢;xH��I4=\X��0�	�Q���P Թt
�qq���!U����Dֆ��'���'\F��Ua��^LAPT'g:� �\���I|�S�O�p⢚�/5`�I��B��x��.�"�]�r�6�x&CK22F�q����3�?	,O.T����O�?�����˧l]
�$�d��P���lVޟ��I� =���3I+�)�'<�0�A.ǌ7|�|���Z�p����'-ܠ1��i�S�Oņ�u��
�.�q2��!.Py�OTU���'pr����� ��ݐ�%+Ntt����.[��'D"�'ݾX�AnŔe̐hq�(�m��$�F�O�8C��M��xQ,0}��Ի�{���ʌ��O���'���/
n��6��?!�>�Ӓ�ѻϸC�I�s�4�c"S-LzE�47��C�	�@�0��hS"�ᯚ�K3PB�I�7�
�� �&o�D҂ϓ�l�B�ɲ3Ӏl�P×	!Q�D���R���˓ ّ�"|�s�l�Ԅ��&T:a�#b��l���?y���?H>��Vi�����<������b��z�	�f�!�ݔ&��!���A+^���k��\�,���9�O�%��H�,N�`C�g�iK�U��mz��'l��'��)�<�,�<[,����`�"I����yb���+Q�	�a%��tV*5�6�X ����&�'m�	�1��	v���A
�Y��EL�ߎ-��$��?�L>����Ԥ���O� ~�{"Y�@o�IB��'$\)���'�4�[����O(�,8C#�<er�ѣ%F
2ax���?)��|�"��X��X����y�$�&��;�y�J�s�^���L�r���g�4��?���'����a!%0T���6��O��L>qAN���'���'<� �lQ�r9RU��K�7�xE�5�'��B_*̜a���o�8��\N	�鹢�O��S�M�䈙�	�<i��[�]�B�;n�s5H*&��pЯ���Π3���z�'�}J��Ѝbrp�(Â˧<�&�'�����~{�V�'�2��4�'�\��bH�}���Kr!�S��L��'���'��'���bF���g!�%7��Ę��d�g�O�TaBD�	A>�z�E�70w�(xf�iMP��b2!d����<�	k~�"I&H �� �ƅ+� ���XCvD�O���b��	:�1�1O���/�_�V1y�mO?=�f�z����	�J0a�)�3�e�` ��
-(�H%(�H��{,�D�O��Db�d��4�<���p��ױ����E�
?�ܐ��'#ҩ+���k�Z���a��-��`�,OP�EzR�O^�U�pI1O�/:�Ęi��`��}�t���\���4�?���?Y+O���O��Dϛz��U34 �*z+0�����38�x�	ċ@(SP˅��p>���;{�<��$��ޠ;�N�d:���Y�y�Ђ��	&g� E�&�A��uHu��EeRP���PG�)��������	��M�����O�㟜�)�e���j�^s,ѣ�Wx�<�6L�'����M �ޕ"�oJsyr�'�r6������'��)��>��D x�卢m�Ҵ[ei+� ��������Ov���O88P.շ$��勅��<PǕ�4`%h�"�N���i�z�`��mO:��{�뜼~�2y"�͖;�ԕ�k.u��HVZ}��,�e�'�&���?�Եi��i�OR�q���WT��$�7bn�	ٟ��?E�l̘<�z�H��H"9'�� ��M����?x��$���>z�Ƒ�q��N��|R�'�x����U�� M�hX�4
��lN���b�O��'�O$�p��o�0�F�L&~��Q�"O�1FA������d-;�|"O�0@��/Mx���,W�6>̼"O�љ��3p8��b��4�e*�����h�U��#1(<��ƭȺYY��'/���4�R�d�O��8�e��D�:hD�z���t@����<p�&��c��jѫ%]D���z!�a��+����}���!y$��ȓS�RI˲oD
%����C�!G��ȓ7�I��� �'�bt���U*+�≖'�`#=E��B��*^��8wF����Q3�+���g~,�D�O�Oq�<�B���.��Ze��2ffԅ@�"OH9�W�;�h�����*T�Mj"O���tnX��ҍ'=FVܻ�"O�=�wC��M�Y�D܌}&��k�"Otx ��MT��&�՟uxh� �|�K*�E�J���=��`#yZEs����0fj,��W��֟���O�����>Jh�Z$Ky�uc"O�]T�_�T�b8�Ã�{��!Zr"O�h*�e�!"F�T�Q�dw�4�u"O�LgIB�wa�Q���-][�L��'� �$��+Q�%�2(K~M@!�=Uuў(rP5�'(P�\ۧd�:[#�c��Z�S���A���?1�pj �ST�m�fp��h�!K$樄ȓ"k4ɐ���&6rx�@��H!���ȓA�vݪ��Y�4�H`�S�Vf�m�ȓ/֬�텶,�.xР(*�PD�/4�'q�J�k2�e��B��r%�O��+B�i>%�Iޟ0�'Y��{��w�B�PCh� BhD(0�'��ase�&H�>)᢯GK28S�'�~x�3�
C<d�7�T-� �p
�'����nȁ^t��F���J��	�'��s�43'
IR���iV�*O2aGz��	�{��d�ͺ|u���M
z;�I�I��Iԟ�$��>5D��S�^��D� 7�8,�T�$D�� $��l�8�0���^�ur�"Oxh �
fڅ�.O dct�i�"O$�@Ch�%\�H���MD,jP���t"O��`�/D��u8veX"/dd��|��'�h�L���g^��s'�*,HNZR��^����~�Iğ���O�PyfCKB�h@�3l�%����"O��Z���HR��,|g���"O��	w�N�I� A���įwg�0 �"Ot,�
-s����Շ�jTHH"��'���Dφt�������uTX�J��L�A�ўD)D�"�'r��RJV���ɀ̓3�@DR��?��C؂P!e�B�xl������.׈8�ȓ2"����͐"?�R�x�����ȓ�T� B� �x���e�#b|�Q�ȓ|�i0t��__�����ʥ{���ER./ڧ`/nM@ ��9�9(@
�Jo�8�	�{=�"<�'�?q���Y)i��r�V�0��2צ͏y.!�{�>��(�!�80!6&O85-!���h4����[�]�\<��.�)'!�L�C�H�B�K
,�t�b�O��n!�d�8�@y1�Z�<�6�`��Xs.�	�HOQ>�j���Q��`s�(^	Kԭ���<�t"�?Q���S�'"��Պ��H85�@����`ppC�)��	��b��>��`[�*[:��B�I�F+^Q�5b�n^��z�����
C䉒4�k����jf�,h�ņ�C� ?�5�p�4�dE���7�1O��F~"ĵ�~�D��D�(M�e�ý$�sc%�?�L>y�����IJ���B��5l1�G/K�B)�B�Ɉq��g酌U�}!��^G�B�IV�����-�����	�A�~B�	�<�Z�#��͟LF
��t��o� ����ş�Iu!ȃ#ü��D� *V�2V�1ړ9���G�$ڥ2{&)����k���b� �6k���'Na~r.ȧIc Y���A5�a��&���yr*Z�����:Ѱ�X$*�yR�S�hi#��o)`�k "e�ڼ�ȓ*��`
2���[��`��Z !OJ�Fr�7ڧw6\z�n_���0�Ȁ 5�r��	("<�'�?1�����$K�h�T�ʒ:��&iM'7!�ġq��!��?���mՌ:!�$G�p�f `� �� �+v0e�!���U�P�ր� Z��A���4nN!�Dˁo�p]�c���nt�(�W	ύP�I��HOQ>�i��<b�e+ro�k?��b�<a`B�?�����Sܧ\�e�F�J�\��E 2'�����ȓu�Z���M�Q,����!��J2V����<���B�>ĸi{� �U��m�ȓq�j�`��?)������*G�Ԇ�7/R�1���-<E�D
SzA%�����Z?VB��݋wߢ�������iu��~��|b�'���O.8 ��Ä<���+ba=zN�@�ȓ��Z%��$=���-������m>��y�"
�+�.�괢�5h/�ȓ`�j�i��� ��阮@��]��	*�?����1m�}ؗ$ ��T�0��J�'Վ[��ɘeۺl�c�̃0��(y�f\�@N$���O�����'����H7[��#�mER!�S݆x��܅Sy�m+�I�j�!�3���26OS(��H�!/�!�D��Jm�a�U�D�c+�4
�џ$Њ�I�[���iD�P,4�Z-��J�_�"�&�O��O��d7?q��Wq���&dM(O�m�F�Cl�<�.
5]^�	cѪݬq6���a�<� D�r �M �)H�i'Rv6��S"OT-I����y���ϢM[P�P�"OJ0q��	&n֥k䍁�5KH��Z�������G�$s!�Q(@k��W�K=:˓9^�P
��?iL>�}C�N9Q� �,�ڜ2CkP ~�j=���� �oª��H�F�l:�t��\Ҝm�"[�"�|�pWL=+�Y�ȓ=��XJ_�P�BE	�7bzpPQ� =D��Mc)�p� �dd��荹G��'�#?�)\?�ņ�3vuBo��B�t���x'����w�g���/���&!�ҀTb0C/�!���_�p�x5$�DD\���%3�!��=�đTg�h��D��+|�!�M�K���0U+��#�����`�8\����OZ�7C������W�M�A�8��v�	iz"~�Q��V(�4C��g�FH�+��?i��0?�e`��- �����E�L\jؑҢWc�<��B�2Uۥ��0SF X���]�<�T,ۻ~�.�R�Q1h2���\�<�`dA$g^�R���*.��("�X�'nb�}�D&^t��ץ�RZfx�Țٟ�7��|��?��O:M�����NQ����"\�4"O�0Z*�Wc�8xsK"O���#�"O��R�V-D~�tf昰p��R�"O�uJg�^�qo��٥nQ�X���"O���O?1����F��\x�R��+����/a>���c�CN�֨(5��4@�p��4Q���?�I>�}��`Vd1�@�6���'�x�<)b�
 8�x�r��v,R#LN�<��%A-.�l!�ܰo1h9	��_�<YfԢ`�lE��n�#x@�X�k�S�<�0��j]�d� G���4��1C�M�I��Oc��O��	�	�^ʈ�F$�j}�{$�'��'|"��>I�`^1<R>����P$�l�"�K�<�-<y�����BI�l���C�<yE�D��]
�E�$-e���U�<1�׮VM���h� ,�05qգM��,��<��DPdiʐc�p8��@2r@�E{b�� ƈ� ���C˼KKP�!(��W�N �r��Ot�'�OL�H7��I��	!j"��"O�m��Gt�`H��FN�k;��*�"OJ���6
U��dR�O�N�W"OD`ڢ��Ʈ�!$$S+g�[�I��h�<ԀeL�j0X���Bړ(^ْ�'�8�S��4�b�$�O��7hdAL�6A�����:�b���)6�Ke��Z�� 
�"SZ�ȓ��%��o,�V<Z�F2)�j��R��U�3�ʁg��ةL�Z�6a��Yʺ��p�Y��ԙ%ǄJ����'��#=E�D�!R�i"0�ޯ]�����T���d�@t���OƓOq�6X��"��AifHN%Ѧ!��"O��7l��p&��[`�AS�"O:�s�'�ly�@�����*C�sP"O*x3�˴'3n�R�j�w�f\ d"O�öd�xs��q$H%O(q�|��7�k��0�-�ĩC� �U�h�Y���=8�h��~������O�X�a��|>�Bf�)qX�S�"O� 0vP>Px��C��:M�$,�P"O>�##L�!�����Q�_���"O�����\�HcL|D�	1&��r��'�n�$��:h�5�7#��3d�Awo�3�ўh�TD1�4&�!�)K�9D�q�R<������?�i�&�0�@@�6z~�8E&�
���-���O~ ��@� TG�Ti��S�? "�٤,V{ �)vG$����"O~�{2i�-!�
�ħH��ta���	�h�̸
�e
R�B�1Х�0Ē���'�x\ۊ�4�����O��G���yg�L�Y��ʒ�)j7f-�ȓ_w}���'�I"�$��8�H��bO08�p�\�q_4�6+Bs�^�ȓa� �r�k�nl��I�mw~���E�y0�m�.WY�]zs��?����'D�"=E��-�':���1D�?I'���RK]�����v&�$�O�Oq�����- g�\F��t4@-�2"OLRsG��hP@Pl����q�2"O�EY���2�ƌ�MC�ei:$	3"O"�*Ղ�zLtseKN�b6�y�1"O�� ��+�l P�d�x���R�|2�2�=���:h���/\�yЪ�H�[�ԝ�	X�	ݟ��O s��|`aXCލ/5:9"Oj�y֠��%��l��"7X��I�&"O:,p�-_'=�.mxB�AH0�!�U"Ot8uj�8q�V�9��:?�]�V�'*��$K�;r!�4�֓.��1@��r�ўh1�=�'|�І�A�f&��U�lU
��?��z�>�RD�38v�x�U!�4܇�~_��e�a�Ѹ��q��هȓO����Ƈ�}S�X�(ԇE���ȓ(A|����j;ll E�ą[���G
-ڧm��u*P�U+����M?Bg����/X�"<�'�?q����� `� $M��0��,����e0!�DJ<h����cC�w��ȑLl�!�<��mJF��2G���(M�!���bni۱�A4-`�у#�@!�D�?�d�;Cf��x��� ���D��&�HO>���&��]Z�,S3�ML<�r�f�0*�%S�y�n�,R|��	
|�����'��F	�,9�bpn@ �J����;I>)���?����wG�QxD�`�\�+q�����F���`�ƋK=}�r���/E��O�`�c%�������W502˧)ZвC�g,Գ��˫x�(G|�AE�?����ODlQC$��O��!w�UiN�.O0��D_:M
\x%J�(?̕uh��t��}���<y��Z�G��B3#�1�:P����Wy�ڬ�yR�'G����OjeY���[�l�Fe���]X�-�O���&_tX��/��s���)�'Qj\Q(W�Hj5����^�mht9͓Z�f�ٵe�
yx��E`����%�\�
8˗%e��,a�gP��yNC�?���������d�4@��oe�X��M֣`tP4:C�#D��:uNϞ�f�&r,(���;ړR�?�q$
ܿ-�t�h��$
k���K��D�Iܟ�d��?�M;���?������O�����j���p���JN:�8��U�L#�q�I�P뜜��F����g�'�I�C�-CBm�"*�F���h��׮�2���.�ת���ɫRP2�Ɓ<�pس"�"$�<�>{*a�I���F{�:O�(�EGU�s?���ʅ/��i8"O��v�؟Q�j�����?��)8��'Xp"=ͧ�?y/O.�:5��'@�!������ b��rr�xn�� �	ԟ��'��'0�ɋ"⹫΍4Bi~I��)�-t!`a���;3��c����L��� 	��pb7f]>�Ak㤜:2@��D�b�š��/ ��D�b����d.ڸ#d��DI�I
������	G�'�d���D�!*D}� !^�_#����'�lb J� K`y3��R�L��,O��n����'h������~������F6#����'���71�m�vnZ���d�O����O�����&�c1�×��4�܉8���8���QƬы�r�a�&s.J �ج+�Z�sJ|
ӧ��d8 �Qȓ�,-�8Fc�s�'f�4i��?A��Dhݔa���"�^�C��%�"��(��*�O�m�c�(H��䒢 !i<H4c��'ö˓Hm����O�8ZE5	��	~��'Z���h����O蒟<�$�O��â Y*:��K6��R���	]���[���:5'�8u���6o��'��OZ��ks��"yVb���i��GH��'���۔�K�<�VYcc�V=�?�0�O[��!R%̩u�!�F�s����/�O���;?%?�秀 � ���H�c�������
�(Q"O������$e{2�B�x��08B�ɮ�ȟ�hhr�Ϥ{"�`Ɂb�c�]3� �O��$�O�aC!������ݟ���^y��'f`Őr��&#ހ�� ����u�T}i�
2L� �c�<���I�q���@�e�&��=Ӊ��>�@��O�-��^ÐtA�?#<qF��&�R�P2/�Q�^���o~�^��?I��hO��(�FU����1;"����Իb��B�I2.������u�Bt��FQb�h��Oc�����'g�I�p*�Z�
���I9ǯϔqBx則�U�M[���?9����D�O���`>�:��Ha �4��,ߵ��U�W�/�Ԃ�?�0�
ۓr��!�Խ
;ޜ(��GZ�8��%$�,��К�A��eia{����?�S�¨#�Ұ�#F�dlh�Sg�4�?����.�8��C�J�F$�*@.Z<e ,��L�1�gB�2�M�"��EQ^����iR\�@8�'}��R��"�����c~�!�d�˃�H� �Q����?���^KŪ�`�r�Z��O�C��YrQ�՜Q0�qÀ'��6��8	1G*[}$p�i�.�<P���ʉs¶��6g�?Vb�����O���O���l>��/�c���d�;n<j�S���O��$9�)� r��\�9���薁* � 
�i��	�@=����E��L�F��'��S�X��?����?iI~����D?Y��L{�υ6}\�qϖ�Tax��'|�Ov=!��Z����dL5k���P��|��O6�{��d���b�`^�0�$u���I�����\?���`�T>�I�,�E��L���ƉwZ~�IDJNK~�!}Rb���I;�ħI�.<�hT _��H���d�\=�=}�̭�G��'@�-���O�]i�u� N�>�TM���ܲ��I��	<���'���.�Ը���Z ��gU9��<��a�'=hy���M�u��e���M�M������^����_�*��FP�5�6��O�lڕV�h؄���I��<�rF]��v�o&��O��G�T�G?��l���"�A�eh�W���	���ҧ�9O~X����0���C �D�"#��}/�,��&	2X�'@콠�Ox):��Ҩ����d��n4.�
@$��^"�J?��!�@~ʟ�d�#-�����N��C#�&6�1�
�bD��Q؟��Q�W&I�$�4j�"k� ���'D�L�ED4I� MX#,V4��q���dӂ�D0��I��O��禵��m�m�5��8���*Gp���$ ��`��y��M�ë	�>@��B�˅#(Hs7c�^��W���OZN�ч%�!>">x�(Oa)�р�'�v(� ,΍=�|����N<W�,0�
�'cjU�Q{��q�K�H#�'[�eC��ţ,�<JUܡKHx 
�'���as�)l(�ZQ7R�	�'�N�8R��q�TXqI0��	�'�<��g�-��mk �͢F����'z(�����~И{RK�D���S�'�����#��&��G�;C��,��'Q�D��-_�8��3�B�5)U4�X���ON�D�O���O.́�̋C�8(�t̞-@��p�U��柜�Iɟ��	ҟ�������͟H�SB�� �(��B�O6G�<Q���M���?���?����?����?���?!@�2��+S�Q~kȨ�A
%M����'`��'D�'s��'���'�Bg0
ݎ��ʈ�s<�`1%�
6K 6��OX�d�ON��OV�d�O����Oj��Ց;�l��R�j�<BG�I3YqqlZϟ4�	؟ �I矀�������ԟ`�ɉ���MK�\�td�C��\%:���4�?���?q��?����?���?	�i�t�"�"Z�X�Bp8Äѡ���f�i�B�'`��'�"�'���'r�'�^�(�lC�Hj��#*�K&h=�W�oӂ���OJ�d�O<���Od��O��d�Ovl0P��P�d+C��`D ����玲�IП|���d��؟X����p�	ן���I�:}mp�ѳ����كa��M���?���?����?��?����?Ѧ�ζQmdM��I�	.���Z&՛��'Z��'_r�'�R�'FB�'R"��	Q�b�(�lK#|h*��2�M%Et�7��O����O����O����O$���O��^m��t� YYt�#@ $Z�=oZP~��'M�h�O�d�����r"���6A��6lcZ���'��i�Ħ9�_�fd"�$G�?��ݛDټ{�F��I�� Γ��$�)�(��7m��8��c� m�	۵0wi�t/�O���?s�1��|B�'>yR�G��IXѣQ�rZ�ā����D%�$M`�'�?a
� ,��-!8��Zq��[��p����B}��'x"6O��/5+hEb��#q|,Ԛ�G>r�T��?��(�'���������ӱ2O�j�ϭB�s�Y�"M&�H"R���'L2���I̎'��D��ԋ]xN�bK�O�,�'��	��M�"�O@`�Y��Ok3��yBM�"{Դ@d�'I2�'4r�Z�|������̧4,�Ķ�(}����r��؛�LͽC\6}���	ߟ��'�1��(KE�~��8�,0✕��U��O���?	��$�C}�Z�T_6���T/V8ꓪ?���y��i�+ٚ��i��Z͖�@���%M�&�`��'�j��Ăǔ|"Z�41�Q%:�P�FI�"l�f����R���B�O��	���`c��N�}JqPC�W,6�`�$�����?9�]�t�	��0�.X�(���E��`���#.:]9ҤAĦ���?���!N_����3������,UL����Q=G�`���yR �D�O��d�O��d�OD��:�'4��A�� l9���%j�	ʁ�	��$�I����O��Ě��M�<����4%A�mM*wa����K�Iʟ`�I˟Ȓ5	V�-�u7���\{ѨC�gUDՒ����L� A�O��Oxʓ�Oq��(YZ<`k�����81��$�L}2�'X�'����-�@����ZA4}��ϐ�S0˓-0�������v�)���*��b�M ;����S	�J�"�����M�S�\���V���.�$�(z�����þ2㾸����N������ �C:���!��;�nT��OTʓ؛����v}�/a�T�1^P�*ʓ87^�X�bn�'qҜm���M[#���M3�OD��
P���b.&B`�ZP:HAٰ)�+r���Jៀ�'���'���'
B�'��85�6�����p�j�ŮK�Eh @�'�"�'T���'^6Md����h[�q�Pq�BCrː�1���Ov�d5��#�	��7m���%(�.�H�*�!%�P�$�OT�򲠑��~��|�X���	����p <=$9)2�O*+��3������ş��	my2ɡ>a���?���Y��a�r�VC�A�W��qo.�#�R��>���?�O>���)����T�T�y��p�)����S�d)��@i� -&?	#�O��I�u&�tR3D�4u�X�R�D�����O����O��$<ڧ�y�K���(�rO,'��at.��?�A[�(�'�~7m'�	�?����r�&����Q���S�۟�"�4Y:�& t�8����nӐ��>d�F�ҡ�Hǭ@���{�+wO�(�7�������O0���O��$�O2�W�r.b5�4bM�:6��o[������	�$?��ɹK;p�C�Ɛ$��!�Ƃ\���O���O�O1�zm��G�6SR͈B"D�{$8!�E���r6�Vxy�	�5
�Ԑ�����$U:Iz�̣�$�ZD�B�+T˖���OJ�d�O����O&ʓ���ßHHw�R�Bƌ���?s�6�;�@9ܴ��'
��?���y�*�$Y�)� ���p�Vl�W�L�h ��4���_$a������U�0����ק��F 4��O8��O\���O��D�O�"|"q�ma�S��Q�\,��Bc��$�I� J�Oz�'Hh�6��;q�v��]�V�Rɑ'۰y��'���'�bhE�h��0O���2`���p�l�<y����.OD%|'(��~2�|�X��Sן����\ a��x���	�"�!���j���	Uy��>����?Q����390�e�P��.׬���3h|��(���O\6Gs�)ʁ+ZJ�<�!W�ژJ$H�,Ŝ�%��m�rZ����\ ��J��N�Q��ߞ�t��U���*B�Ԫ���?���?!����'��$��D�%H���<H��*�4A��O���O2�l@��g0�	џ���a�Y?
1 �$ֳs��s��I����l'�Eo�H~ZwQ
�ԟt�3��J#H��63��j���9s���I`yb�'�R�'�2�'�b�?���W�&)��U*(�d��N�a}�'���'���yB�u��牉!�8�"�Bq$9��`T3y����I�I8K>%?���殮��%�Hc�X�[9��)�i��=����ɀ4|����'���&��'�"�'R& �]ذ����@�P���@�>SR�'-b�'�������O8���O>x���Y�*���"�"K&�]��I)�����ĊǦ�0ٴ9��'v��`7�	�� (����J%~���'*���n2�sV���-k�	�?����'{��̓|��-3�J�`�|8��/%85
���柌����I}�O��d�]�t�0���n\Xؠ�ǒ9��J�>�*O�%oZh��
��0�p�d�:)�h��d��=�?�nZ�M�2�iɀ����	��	�i�F*��O���
��!W����q�		'��$*7+�~�Iy��'�"�'R�'��iS�M\F-h���5<q����y �7��D�O���O���
�D��n)j���@pӤ'�
�*�'���'�ɧ�T�'����6;��Rv�ת(��J�Z�x�`�;3�ij��'j�♊��O̒OH˓3����aKY�f�*�a��U���2���?y��?����?a(O���'��� &�#e��a3�A�	^#-@4T�'�\7-&�I?��$�O ��y�P�Ay����ݓc�Z�"V���چ6�&?a�J]�7�h�|�wkֈ��`Ga��6|B�X���?����?a��?	���ZH����9G�f����C�j�8�P��'���'�Z��?���R����$V
#�� BR8~�j���T&�'���'.��B�,Лƕ���u�H�,�
'bY�(�-Sg��]"J���O�O���|����?i�mz
ԣ��� �l#��܎8�B�����?!+O���'�I���O�֙�A
@�Sy8&�ϡ9���*O���'�2�'8ɧ���KAD���ӣ�z����I�`h��/6@}y2�O-������t�P�
&�޸[5��Z���1��?Q��?i���'����ʟ�f�D������kQ�"��r$��OD�j����DP~}b�'���@�A#
rj�޶\��i�P�'w��V*�������8p�'��i@+Q�a�u)݀ n!�+X-bBU���I�x�	ڟ0��ԟ��O;xi�m�"v&��a�ԑF�$�1�P���I۟�Ik�s�l��4�y�l
^S��v",,��|�k���?�������@dpq�4�~�oti&���R�$���v��'�?Q��_$.��e�Syr�'����N��كB��8�r<ڢ6V���'TR�'�#����O0�D�OT����0U�B�$НyP��Ǩ6������O��$�]�	)��t�y��e��vD ,�-O��c�E̍C������ӝ�a��<���3I����,GH��LP0A��Iߟ ���D�1O�	jB
��d�ܬ�q�S�BbB��'����?��8�f���Y��ꟿIT�X��7?Sd$�H�O~�o���M#�iW�TX��i��Oy+7e����[w�$��SK��,�<^��p)����d�O����O$���Ob��H�m�ҕ��!z嗀x3iT�3�z˓UX�	������&?���/}�<���&;g�����$0�0��O�0o���MÄ�x���Û�;Z��SQ����J��\���#W>"��)�'�~e9�'�SD�|�W��Jv�ِ5|*4�%����a�*�ɟ���̟<��ٟ���Vy�B�>��,u8�G,F�Yצ�yW��(�x���_ƛ��$q}��|��8lڭ�?����a5P����K�o	C�K;���nb~$̏/A�h��O�'�yW� %�ũS��.1�T��1�?I��?A��?Q��?���)��p99B��,l��}S���)�2�'Xb�>	���?p�i�1OzTy�]�~,�!) �Ǌ5�TP��'�D�O0�����h��`�J�j=<�oۇ+~2vPs�D`0C�)X����������4�^���O��ă�9V��2��&��W�~����?�+O���'�B�����}��A@�_�v$��D��x�|��������Sy�'�v�?��?Ɋ��3 n$��.#lEqŊ��U�>�K�A��W����?)z��'��!'�,�'G@�S+z����пj� �1.���|�I�����ğH&?ݖ'����X�����so��!�|)##@ʰtb�'���w�
���Oho�������N�2��f�:U���4;�V��5y����̹0�3�Ė�(�:=g�E
�'
�]Ԑ��!n���?�+Ot���O����O���OL�']T�]��V�0:Ԓ�ǃ��H�S�O ���O���:�9O �o��<9ā�5F�l�M,Gd���pETޟ�	T�In�}T in�@?ɐ�A2%���{F�2�� ��(S��5g�(��<�'�?����
Dy��L�m'�l�dL�?!���?q����Ĉb}��'("�'g�0�6	�1��!Y�>@ZY
����k}2'g�|5n��ē�����#ӹ^~-��	U�"��d�/Or(������;��6����?���P��%	a��Mr��E5l�Be��O����Ol��O2�}�'j����%V�v-S�'�<P�F��;o��Bym���X���(�R�꜋t���`)�!Z����	�8��ɟ(�w����'%:�Q�Vx��l�0;�<Т)OU7�,J�X�������O����O���O��dM�M:��H�~�� �łBSf�2���˟����%?�	�0��� eT;(��*!��l�
]�O����O�O��O��d��s��В�%	��B�H)��13Hd�P�
��`���&���'�Z��!�\6 l|�E�@�)3p���'\�'��'"bT����OF�$%��Ac�I;7x�I��Ά.	��d[ߦ-�?i�W� ���̓R%P���)�|W|�K�̟O0�\X������'<Y���H�OU�΋�sب�!_�{�r0H!:K�'>��'�r�'"�\:�5!��G1<�Rq
R�ޑ9z��Oj��k}�S��9޴Ř'�2��UDR�t}�0���O�*ox �I>����?��U�����4��䆩?�:;4�D'�ɻ��/\n1{!��~"�|�Q��Sğ|�	՟<X��~��s�9*�b��siß(�	ry���>I��?a�����A�a>\��I�`Κ83���2���1��D�O4��&��~�#�A�J�Pd!�F3]aژ��	8��3���Y�'%�D�x?aN>�A _� �6QC&e�Fh.t�R͗��?1���?9��?AH~.OT��)� >�R0����L���E29wN]�s�'���'�Z6�.�ɨ����O��6�T0 �� ��Ɣ���$
1��OX�䖖<i 7� ?i��?�b?��`�;ۄщ� ҀI���Q@�O ˓�?���?!��?)���)*<���� �!++2���Bʽ\��듑?i���?�L~�<P��9OaCČN�(	"���C��iP��O��3��0���(9��7ͣ��(E�P�u�P��t�2k��Qr��O�h�����~R�|�P��S۟�:�*�9n޴�y'�14S��c�	۟���ԟH�Iuy��>����?)��{��ECU.ej�m��	y0b�BJ�>���?�H>�ud�+]~Ҍ��d
m`X��N���^�4�%Hr	q�:��|��੟�ϓmFBED����A0`�An������,��ϟ��Iw�O���J�@y���ł=>�l]Q�G��2��>�,OLUm�V���R��,t�D�`B�CI�	M&�?A��?i�YzZܴ���Q�C�@���� �m��	*�@R����67��ڗ�|�X���	����I����Iڟh�M��r�1��48�"ex���TyĮ>����?�����<1�oǡ`��4a�]�Y���� m�	Z��	���IG�)�Ӻ���d�1	��7J�X��`���B��C��)�Ш�O�3K>�(O�$��h�Oz�[���.$��f&�O:���O���Oٴ��	u}"�'���iC8K��f�	W6����'�26�)�I�����O.��k�h�uG�1\E:c-�| �T�X�57M4?�l^"�t��y�ӼC�+ϵD5V��T��-��XO[̟X�I����Iğ��	���D�ģ��D�q��=�:�S��?A���?��]�\�'8V6-+�	�),�8��-��w����)ƕ ��O��$�O��ճ�6�:?��,�x�ƅ?	�&��$HV'G:����ڇ�~��|]�l���$�I���[0e���&9�Qn�3N�¼IcS�,��Vy�$�>Q��?1����)��IV:�� b9=�����Bk��	���D�O���+��~rԡ8}���S�S_��I��"G{
`A�Ц��'��4��h?aJ>!qߙV��FK�2H�@�܋�?����?����?yK~*O�\�	�B	0��� �;	d�q��%v�^�$�<i3�i�Ov��'O�/>������G32�a�%�+K��'�r��԰i����"�"���I�'z���w)ͮU�\��	�~:�P�x�I۟���ʟ�Iϟp�Okzu��f�5`��i��	"�\�Y�U����4��R�s�H�ܴ�y��Qi����`S	�bA����?�����'�F��۴�~�'�/�pIVS�VYR��҂2�?��[�u4<�IU�zy�OW�N� 3�T!�ŰÒ��T�y���'���'R�	����O����O�xZ'F��WE�2��J?;-`��
8�����D���0�4/��'R�LBQ�NtM�C�,�d`y]�,хh��'��!�-?�'(L���y��Fa�� �B���բ����?����?y���?��	y�[�O�������� m�N�05�O"x�'�b�'��7"�	�?A��ĘL$0��F�2@Ϫ³��柨�I�
�4p*�y��4�y��'�U�2I�?�;M��aBȋe� �b�
� "�Ե%�Ԗ'l��':��'��'r@������q��H�77
`%ۑS��K�O���OX�$9���O����J6~�H9�&�  ,PY�QA�`}B h�r	n���Ş6�p�`¦X�&�d�P�I�:�����v>��'������@��|�X�����G;��s�G1L�l ��(O��4�I��,��֟���Vy�
�>A��/l��"���{h��3n�,�E(�o��V�f}B�'�Ҥ�O��T-�6tK���g��?X�D�B2d�����d`�%�'D�T�Il����
����e ̈́|�����O8���O����O�D�O�#|zu+X�{n������G�ȥy џ���ʟ��O����O��n�R�=�V�H���+F�������Jt�K<��ib(6�⟬��N}���z"�P��͂����ꀀ�K�&�Fɳ�H�O&� H>�/O�I�O����O��Y1oл�|hǄ�|Jpx��c�O��d�<��^�l�I؟\�IO�a�=a��#e���p�<��c����Du}��'���|�O��H״GA�!���ɰ]�6�C���^qt�{��L:yܛ������3��9��F�D�� ��H�v��mc7gS�[����O>���Op��*��<��'j�z�O��Z��t���Thƅ���?��`�����A}B�'L�����C�H��4IV/ ��q�0�'�!C՛:O��$��`�(I?�	<!t�`堐�%>Q0UC�d�H�	JyR�'n�OsB�'Nr�?	!��Q'[��UZd����"��\}��'��'��m��<q��5e�=����@���0(M͟���A�Iퟔ��џ�8�.��%�4l��Vθ%�ґ��'9�6aq��kռ�+2I���%����d�'���@	��KK8�4$�^a�x¥�'���'{2S�(�O����O"���!%=�4j�����P�M��x�0㟰 �Op1n��M#�x���x�a��^�FR��#�B�'�)*���D�>��O�i���?q��{���"�)#eȜ9�o
$5�^9z���O���O(���Oң}B��� �\hr���h=0I3䗴A
P4���'d:든��Ц��?���2�ـFAQ�"���[9�rD�(�V�t�p0lڳf�&�l�e~��r����1�d�#� m����!� �$��`�|R���	쟐��ğ��I���7�)�2���f�f������Ey�@�>9.O �$%���0C�H��O9��De��c����O��l�	�M�P�x��AV�9�E�Lf.�I��a���b�S,C�.��'�:�oJ�8�P�|�_��jseD�=������*��h�G"C�h�	����ԟ��IEyb��>��	���jw�Փc�����O+8C�Ԡ��[��V�$�a}҉� m�-�?���x��}��3@���DmL��$l�^~���1`vp��m�O{�_�oz:H!fKH���aC�-l��'*��'z��'7�������'-$�#�OI�E؆���O��$Fu}r�'�2�`�`b�d �O�*�`���*Q��H�(2���O"�D�Oŋ�Gh�T�ӺS-N����V�O	,��c��;5%F���'��'��	���I�����k�f	yd��K���C��� C6$�Iğ��'P`꓊?��?�˟��S�΋��h9i�[�G��C�W�ĳ�O����O֓O�{�&X�2�>��9�βYB��Wo3P�Em�+��쟀���'w�'�60�@	:\�*C��u��`a��'�r�'NB�'��O�ɧ�?����d�XjDi� �����LI��ԕ'v6�&�	����S�ՠ�^�.I0���M�.���x$AӴ�M���i��q�i��ɶ/�0ɡ��O����Oy<��(@.f`����Ŗ�������O��d�Ov���O��D*zULԦ(\�;¥�%Cc��ǃ������O"�D�O������1ϓX���ц%[sl�!Q#Z�E�6���4'ۛ6�<�$����)�.,Z���;O�$B��O����AT$̑!��O�������?iU!+���<���?y��@�= p�Y!��&��튰���?����?Y����L}��'G��'>�q��n�"3V� ���hk&B���GDy�'E�v�#��I(X���� h�&\��D摇�B�'Ѷ�c2�\v4QH�O����9�?�x��ؖ�Y�%Bάs�h��cK^$��j�O��D�Oz�D�O0�}*�'ϖ� �eY�Eȴԛ'G�5b�E��i��|yR�y��L���~��ّ$Ǽ	6ܲ��>'V)�	��p�	���� ��榽̓�?�e�^�|B�'�8�ڀ��&}��q��
)���&�t�'���'�B�'���'��L8�F�e5^���_�+���WY�\��O˓�?�I~����q5�H(n� �K�,��*�b�Y��ݴ4ϛ�7���
,��c�C�Pc�����]�B|eK�0=&�I%!L��R�'pLx$���'J��*�@��T3��4C`��'���'(��'��[�(�Od�$��s�A��\Np����:��Dڦ��?a�V����4s��O�9�u��� ����5�D��>="�/�y������D�Hf����f�eIƋ�:B�9��HD�tĖp����O���O
���O �D�O�#|R��ۄ�
w�M�*b��sӌ��h�I��*�O��d�O�o�m̓zM��
5ý.`�Eɱ@	�>ἀ�O>��4`~�F�O���x0�i[��OZճVD��j��᧯Jp�np#vDA�*�Tԑ�{���O\��|"��?���n84�A��0��1�% ��A{��?�+OD��'n��˟�OC<��"�ٿo�EBË+q���A)O}�'b��'Yɧ��'k�v�ɱ����(ȁ�ۏ*�dy2��%8B��������Ju�"KV�I4�@0aF�R�qo�в"��fb2@��؟���ޟD��`�Uy��O���U�6d�T����**TzDCA�'��	��M��b�>���@���)	�=3F$�����Qy���?1DN��MC�O��:2B�SU���� &~��%ȕx���WM��?I*O����O|��O�$�O��'D�Ȋ��6W<��۲�ȴ3Uʅ��O����O��� �9O
�m��<�p*�	"s$m�/V%�+��I����q�It�
p/��nZ{?��B�.F�q"n��9�����H�(�rgĘ'��%�Ĭ<I���?9�ꂢE��XZq(�d�|�����?���?�����d_k}��'r�'��u9�T92^F�Q�IuK��K����r}�'���|K؎�Έx�:u�~Б�b�+9��	/j��m�`��ܦI�L~�ԁ��LϓM�(�ʳ�	�t|B���H�W�,��蟐�Iܟ���Q�O^��X-�U�FL�6P��(6F]�`�>I���?��i�O���*r1��z�b�l4ᎊ7={|�d�O&�$�Op˕�l�"�Ӻs�n�7���-���,�)W(UV'���9��$���'&��'�b�'"�'�<�rj�>q�@�� S�en�['X�X��O���O\��?�9�╪@ �/�pP�!��$h�:`��i}��'�R�|��D�ăj���1L�=^�E��K�R����i��_�"�����'���'��`CgM�#��Iȴ��h�1U�'0��'�2�'�2R�h��O���ľM>�=i��̤xb)+��."����RӦ��?�T����� �-�2�DJG
N�FlJ!���'�A%�ߦi�'u��tj�|
K~z�wtF�+��Ӕr��3��3^z���?����?����?Y����� �@a����3sB��HB$HQP�'2�'��������<��L\	J���Qǁ�g���eN�a�������ퟸ�DEȦQ��?y$G�8`���F��O�0wj�� S��|&�4���t�'~��'�R�RBIU#�D�ɧ̓=(��i��'�2]�(@�O�˓�?ɟ��Uo�A,]GNfh�SP�\��O����O��O�'Y[ҁp���� �잘�r���#�ޥo�K~��Ov������ �;��K�}�>	�eʅb���?����?�����������2a�:(�RQ��}��E�O�˓E�6��{}�'b>�3��׿.]dA��N�Kb�'s�t��i<�I_���9���Ҝ/cH,�p�<0{v�����/NBV���	̟@��֟L�Iџl�O�@i*a�E�~5`��^ y����Y�,�'�B��T�IϓjB�`mA.4#�UA�gI_\�����&��&?)�sÏԦ���싷��<q|UI��O �`�	�xM���s�O �O���|:��_)`���#@W�@Ja�ƸQ�(]y��?9��&7��<qS���	���	�m�L��Z�4Al�	_Sh�a�;�����$Gڦ�cڴ`%�'���
��"�MJ%�G�r�< BW�d0� ���� �O��� \�<ɑ���/���j��5,@aÅ۟ �	�x��ӟ�D�d7O�8� �Ke@(�d�l9�0��'&Rꓦ�D�ަ��?���q��j��h�x�E�'�����n���o�ZtlڭiQ|oZB~����FQ���T���q�̃'.d�Y`�\�E^ �ě|�^���I������ �I� �f ��{|~��b�����tI@y"�>����?������<A�O��@�ajdHlN�b$����I��M�նi��O�	⟆�ɗ�[��EX�d<-���e�F4ZR�ʔ&]G�B��\HQ���O�SK>y+O�(����S���0�t(�ؐG��O����O,���O����<��R���I�p
�(p�F�w��<�f(9%N��I��Ms��>y��?љ'�z����� 
4ɣ�ʚ�m�Dka.��M�'��Iڦ���Ox��?�̻/(�!1fbª`�x10��LĤ��Iҟ��ğ��ȟ���~�Of�|�C/�Mr(��@I�x[T�Z+O&��i}��'w�n�jb��;��٧2�j�!aϾ.tS0�,��O����O��	b)j��ӺK� %^
5�N,?
�cG�1{_�@�'��'a����I�x�	2t^���AV`��i�SI�9��d���\�'�\��?����?ϟ�� ���ض��b(�7u��[0U�8ʪO�d�O��O�.���2	�
��4kEL�.E~�����'F=m���d�T8��'��'/��؅MT����	�&I$���'�r�'�R�'P�O�剜�?��'�`�v��("5��Ο���Ɵ$�ڴ��'����?��ĕ�'���"�y����d�9�?a��bP�ܴ����h�j�b�?��O�A����]�z@��jb������$�O���O��Ol��8bW�5��fʋ�|�:W�$��d�O:��Ob��>�D\���Γ7τLbIڵ^�B��C�ְ{,P���ܟ|�M<�L~j���$�MC�'뮝���67�.̩v,ʖ����|i�S
�O�laH>�+O���Oԍ���L
-M�4#�O�2lYI���O����Oj�Ĵ<ѓQ�������b0r�埌YP�h⵮P�K1nH�?�WY�����H�M<t�?}<��#&��C��q� ꔅ��䘴z.�p��(T��i>ʑ�'�lq�j����&���&��/������`�	ޟ(�	o�O��DJ�[!�L D�+ak����藅 J��>A��?� �i�O��i��zV��`�B�[.���(�x_v���O�D�鈴�.�Ԧ��'~qT���?�;$F���d��e$t#����o���$�x�')"�'���'��'+L�ڵ�6 �����qIY)$P����O���O��$;�9O�;�ײp����'��y�r�:��_x}��}��)lڎ��Ş$�Ѣ�ɝ�
�"
MH<HJC& �q��i����(@�2h0�wV(�O<ʓ
Wfl�$%�&!�+wfҘU��a����?y���?A���?1,O�]�'�B� �a���m��a�
��2Kb�<⟔��O���O��	9FAq�C��ƹ`b)˵p�0tY�@�u�'�¡ð,K�O���֡$p�8���;)h��S.��'���'���'l��S�:�0���2�thH��N?�����O:�$�J}"]���4��'�DȊ �r{:��!܃{�)O>���?���e���@�4�yr�'��%��8 �JpP��>NL��&W�Z������4�����O���Sـ$*&��5�^�zV�Ʌfz���O�˓6'�	ޟ,��ɟ �O�][��|���c�B�Tf�H�-O\��'�"�'�ɧ��Ǥ	�"bi��cQ��_}�-Asl�]g�6-YOy��O�4����^�ڍ;T��,qy^����!idL���?���?�����'��$����#��\�*&��r�
�	��3
�O�˓�v��D}�'�
Бe�J��j���������"q�'�2lO9���9O��Ӕ�h�����\�0�x��K29�Q)&R�i ���<����?���?����?�Ο� ��Ò�P,r��+���� �P�g�>����?A�����?�&�i^��GL��2�萷>�teۆٸ'���'��'d��'�.P�a��>O��уAT�=�: yu�T�z]���0��OBU��/B��~�|"Q�@��џ�k��[$B�L԰�/� U+D�*��Mӟ ��ޟL�	|y"��>�,O��$ќ5`����ܞ'�y0dꐲ\�"�DC�Ob�n!�M+đx�S"q�-�s.�As-��=r��ɸ,�AKdH8O� '?)Se�'�Γb���CS�[�岣 �&@���I��	�����J�Ow��x�F9�A�n��=+��(�o�>y-O&UoZ~���ʗ��5�vy�����O��x"�(M=�?a��?���O��[�4��$?�`,b�'�ug�
LTT��5E��HЉB������O��d�O���Of���+z�~T�צ',��"��&.ʓG���L�	͟�&?E�I�H1Fud+���S@�;0Kʌ��O����O̓O1���@u��g$)v���v�}X��Pj�6�8?����n9D��d��wy")�+I�H)q܃{��pGh��`�R�'�B�'��'創��d�O�áK>zxxZ�Z89�̽)�r�`�r�#�O���O��I��̼b2e�r��!��UnKPT!�b���WA�-i�$�'�y�H� ~�B��Q)�he���?i��?����?����?9����}H ���K*�ب��9V���'�� �>!-O�qnB̓Y��a�0�A��������$��	۟��ɳu�Dl�X~�bV w�D�І��>y�s�V�(�ʭqlDȟ�Ƞ�|B\��⟀���\�K[�4�:�F+YP���.H���	y�H�>���?	����̏E�HH�7�ɡW��`:b� ���I�����O��$;��~ꁁn萅�w��]�pS�댍H�][E��{-���:�*�ONP�O>������D�>���/�?!��?���?�O~�)O�5�I�p/��3�n
��t�%��==����<��i�O
tԧ-7텸R��-1C�:+V��딈M�����Of�i��s�"�o����n�*�֩�3A�/3���%�ၢ�ҟ\�'�r�'n��'���'^�#1� �TL�9��A�*���'��'�2���'�P7me��c���T�XwG W� ��5O(��5�$�i��Ur6m����H�9J䢜��oP�d;���5M�O �#FΈ��?�#-���<ͧ�?Q��̌��l)�h�� ɣ�?A���?����D	c}��'���'j
x[Wa�$ ��G'սv��������s}RCt�Dl���ē
�L$� ����B�-S�l	~ظ)O@4�vʄ"U�B%�a�/�iG��?�a�f�l��O�]+b<��i�����O���O����Oh�}B�'�z9s��F
L|R�ʔ'�?s Z�G���fyit���#PN�= 0��J4��Zi��ɓ�MC�i��6��>_t7j�����0¬���OK��M��j6�X�@��W?���	B�	Uy��'���'��'I¿p��eg�-/��� a�
�"�^��'����?Q���?�M~Γ�6���޴#�y��샖G,��vY����4lϛV�(��)K�����W,޼X��=�'�Vzڤ2���~ev˓Y]�8��*�O�O>�+O��*d3;a�s��9r�.ܑ���O��D�Oh���O���<�D]�8�ɶD��V@ΎXڦ�KB"�<!Q8����M�B��>���?)�'sb H��C����ʦ��c�
����L�M��O���ꆜ�(�.�����I��Q ޟO8����?)���?A��?i����FQ�"$R�k��S2����ZY/�?���?�U�,�'=�6-$�ɶM�L����R����!�3Y�d'�\ ڴ͛��O9Pe��ij��O�l�
����3t���8��ј�
���h��A��O�ʓ�?��?���+�Ơ	�;-�!qD����!��?Y*O~��'���'�r�?Q9�/�)_�ڨ�6nQ�Ih$$�5Ǫ<فR�H��ş�'��O�0�2���Fꠅ�c�ȉkd8��Ζ�vM�ߴ�����'v�' �+�aš<�"5�IR�h b��'��')��'5�O:�Ʌ�?�S��'u�x�Q/�v�~Ȋ3+Sǟp����q�4��'(�듮?�fA[�D] ���
�0�%��e�?	��A�ڴ��PWa`�Z���`�G�"|�7*ҙ2�X�����?Y,O ��O\�d�O���OV�'��z���9 ��1N^�i��آ�O��d�O��2�9O^Do�<�V�W�q����=jETqt��d��N�G�Sd�l�C?!��$V7vI��F;^,l��IşHbuf��hB�`%������'��㲪7I�l��F΄%����'�r�'�R\�@*�O��$�O���בa�X�n�>g0�B��3���ªO2�d�O8�O��P�S�Z��'��,2���3s��O~�$܈V2hP�T�
=6����?����'f.Yϓ+`%@M�	��.L[����̟��	Ο|��D�O+�Dɞ5�o��"�nE��MN� ��#�>�/O�!mZO����!E�+L� ����	n!
l�&
�?����?���k����ߴ��D[�*�����'�u��L�;�*$�MW�O��e�X������O����Op��O��$*� �q�o�40N��NJ5nA�Y��Y����O���O��D#�9ONPƢDlI���F9!u���p.q}b�'Wr�|��d��{��4a��ƴ<�r-Z7�q���i��	�h�,3��O�O��{�ܘ�AQ��"���GE��(��?���?i���?�-O<y�'$2Kޢ%����"�N=����IW9<�Gh�P⟰ �O����O �	��SՂ��f�0E�=^�;��p��0�:xR@&�'�y'��zT�<8����,���ۓ�?���?����?���?	�𩅲U�f�!l��\'��Y]!8a���?Y��b�	WyB)k�
b����ҝ~r\�!�?A��L��&���Of���O:�*�Du����&��ϝ�S��ݚOJh�sR�؆O����|�fy�O���'�rȀ6ZLB�
'&0~�ޜY�"\ ��'G�	�����O��d�OZ�'\�@�S��M��R�e&\Xt�a�I���	{�)���5~�ff���<����ǥ�;6}�XC2L��M[S���a��/���ML� IÈ�12R̫�a�4(�&���O&���O���*�ɭ<��'�,�6z�x}�3̂3tg<�����E��?�3\�@�	Y�ș4i� :%/�l<��Iޟ�w�����'z&���@A�'*	�| �E˱#~��Q_�HD"#��O0ʓ�?a��?���?�����i�e����aɎM����bժP�듍?��?�O~Γ;��F?O\�$�Ău+�b��G�)�Hh+�'��|�'Mb�'����iE�D����ui'fi��T�H�(����]�E"~�P�'D�'=�i>������(��O+$��D0D�5p�F�I�����֟$�'� 듬?Y��?!"Y�(h���*B�)�ś���'����?i���H�7�X$W��4k�<�:�Y,OJ\�"��4�7;?ͧN�:���<	����50d��`�!5�|�X�j��`��ȟD����pF��8O��!�B4sIZT�Ti��������'tH��?��������hf/J�RV���a݂�lq��%�O����O��B� �7�*?��;�ru��O���8��'4�b'�ż"�n�|BX���Iٟ �����Iܟ��>Qehm#GI�8P���A�@YVy���>����?����O��a+�GO�?p���f�G	V{J�(�û>���?�C�x��GQ�Н���
$��ѡ�KL>S�)r*����Q�8k��S^b�O��X��ۦ�Va�]�%� �~�����?��?���?.O4��'��X-f�,��"ΐ1�za	"�b\b�b��� ��O<��O��I�}�R��ֆX_�t+'�@7c��@�KtӚ��,�������>�λS����#�Lº�e@�4P�����IП�	��t��G�O���蟄���A7ğ#v�U���?���as�I_yruӔc����g��	tET& ����!�D�O�d�O>8�E�{���G�}÷���![�=�m��� �J ������4�T��O|�dLg����p
 �F���q�қeX��$�OLʓ[_�������\�OR����ט9�5ڡo�D�yY/O���'ʊ6m�Ԧ��O<���[�Əu
�L�c��$.q�P�ρ�u��ytHO6��d��8����i�N�O:�k&�G�.NB蒀�[��؁��O<���O���O~��@ʓN��i%���H�`�7	jU:���?I���?y��i`�O2h�'�r�\�!6���ř�t��2EĮYt�cd�8�� n��# �:��`�JT��e9��_�9zMQWJ^3q��Z�L�����	埨�	˟��O���kԏK`�ܺ��B���9�[��Iğ<��P�ğH�ܴ�yr��$Ί�k��~���%�7囖�yӊ0%�8'?���7����"C�7pbG �k"�ؑ��O8�"uġ�?�&b0�$�<ͧ�?�BiV	,;`���e�ch(������?��?����$�B}�_�x�	;�B�����y��僒$C�+�&��?YSU�$��4�O*�$�*�S��N#W�8"�^/��˓9�r]�'��02�@X���.�쟨�@<O�T�CU�~���y���#t�j|r��'y��'���'��>��^;X��a��Y�H�K,�[hҁ��!����O�����	�?Y�'AN��`lU�gC
�W��:;��-��'��i�N6-ڟ<��6�3?�w�Һ7���)i�A`DْRy��𩁜ZKͲM<���<���?1���?��?$�z��) ���7w ��B���D�J}�'��'��O}"J��L$*,#��DF�8�L8T��X��f�o�R�%�b>�U*�-�H���86�U@#cɁ*[�]���=?��&ՒV��Ă�����D�F���4,݅Z��<��N��BÎ�d�O@���Ov���O4���	�l��N�;����L=pW ��A�៨�۴��'|��:��Ch���I3C& �D�Ѓ#���xvP&!�2}��cr���B��Q�,��>a̻q#<���$�"��y�Y��y�.�������4�	ԟ��	ş`G����z]�];1�OO�ۥ F*�?���?��\���	���	�4ޘ'r����'�Vk���2D��NH �K>����?��'�,�ٴ��ď�5������W�Z�����KЀ��~|�W��͟D��ҟ�� �I{w�:BV��"b�7Q3Be���'�rP�D��O�˓�?�ɟ�Z����y\�i"BmT$k%Jm!uV�(خOJ���Of�O�'.]45@��W.>�,+g��b���2GS9~�:�l�~2�O��=���u`L���� /�� ��N#Y�~ő��?9���?Y����'��$�ɟ`!CeD53M�5�2�)ф���ON�d�O��n�Q�G��	ߟ�"V�7Ɍ��/�4�B���G����	y���oZ`~Zw��ّ�ߟ\�'CY�(pq�/ �5)qMH�I�Bܻ�����P�S�ì�����Q��0��%�R���NO�U�2|�5�(�٢�n�4uX���̀5sR��CD�( �~8�� V�6u�8�%!p\y�cl�>a9e	��ˎ)K"(��F�"Fv�Й�4fju�dj�&�H)�$f��� �#'T^��ȓ�?R^�pّ�(^�@�i�2����d�"Zj����A�a�`3�;'���$��&4zP�� ��2�W�6r:0�P�D�YdM���/B5ȳ!��h<ڴb�Y2`��o�s�:�("N,��0��h�.��F.��|�"p�� E
@(�m�g�j}iu��o� pC���y��S�R=:����O�$|벡��m��rs�RS���K%�� Rxx^���WI����n�:3:����!+OX5q�h۷@�.1��%��+����5D�J�2���ĉ.��aX��
	UW<��5� gz�8�0H�?��@0�G�V�BQ�fƌ$����0�r������L� �3D�΋A��8�4�?����?y�{��Ity��'���C�+b\1_ �u���t���?11p̓�?����?!�H &��T']ֈ�8�NE6�?���?-���<	����H$چ��l� yp�߁�X�:-O&i�A!�d�O���OT�'O�����M��p���[f'��p�	+��D�<����䓐?��K9hl�-��$���7�	�t1�٧�?�)O��$�O�&�	>uA�H7.B���FY��m���O����Ob��:���O`��4���p%�cU�WV�\J����l˓�?��?L~EY?�I.~�QD��H<�xC'^7t{���IşD$���	ş�HPL�O�<��x��ЯA�TP 6H�4K��m�I̟�IEy��'�X꧈?����?Y@DO�Y�������C�������d�O���O��$+�|�'d���2j�R��d�1�n(hMb[���I����쟨�Iޟ��'�ԍ��C�i�.|����*�r����'>��'}>��������K�ޡ�@ʳu�`�H��K\"�'��6M�O���O��T}�X��F/ݲ8"�ݹfM��2�� f��֟���*?���Oj҉�H����q�-1fbM���6��OJ�$�OL��Y}R���I�<Y����rV�W%c~A@)�K�
���RI>)��?!��3h��U<r0�J6�3_~����?��� @�	]y��'"�'C���u%Wl�8K1�Β�4$�DV��C��ꟼ�'g��'��?yֆ٣Rvl*�cR�7.�)#�e�O0�'�����$����������S� ��5�VG+[ z`��͓�?��%����؟��	s�1��`KѭK�|�Y�\+ar�4����Ȗ'�r�|��'�BJ<��䈈d�pa�,M�i�H�xn�����I��d'?)9M|J�I7bw�Qs���7�t�cM��?!������4��D*
���	|z@jFN�����s"ޟ|��㟀�'zb "��Ot李6v���^���O9x0�4��,�$�<!��?�L~�g�JzU��s�f5
s	��������d�O nZW�T�'#�ư<e�߭{���	Ux���
��b[�X�I�&?Y%?ݲv!��[<>��p�Y�F93��O`y"�'^B�'���'s�)��� !��S�� (��(;�kT���Z|��"|�3�A89�~�a��(&��L�u����?��?����?Q(O��n~9|tD�㶊�4�Te�5/{~lDx����Or扗L(Nl�N4j�`03�c��(�.�d�Oh�$�<i,��⟘h��dS�͑�̝�x��͠V��b�IS4b���IGy�8Ox1g�0H"�3Ab�GR�\�6�'�ϟ��D��?��'���uJM+S`��qN�b�(B�"X*I�'���'vr�����zS�$R��@����	��ѐ!P�T�	ȟ�&�P�����'dd�c7�T����ra&^��P3�|b�'��@yrV>��I b��m����I��Pp�G�=Iz���F���?�(O��C�>�ʇ�s-l�`dfR�
����'ڟ���@yRZ���O�r�'(��T�HT}��%�2F��8Ǐ�(@�'��_�ܪF=�$�bd��Ƚw>�`���_'1����D�O�lO���'2R�<�QE�3#�@`M��P�˔�˟�'�r�'�O��O`$"��0;��əQъ3����'�B�}�x�$�OV���O�'��Ӂ֤̀�Ќ1K,%�@��K��$�OR���O��O�3?Y` �-i�b��!þ:������%�?����?����?)/O�o~RM�4�4pF�%`��2UcɄ*��Fx����'�R�'i2�3q��B�
��ы%�T����'�"�'U^O��U�5G54�CE��Z�����[��-&����Oyr�'��'>�':'J�S"�/ָ��  �v)���	x�Ο���S��Ny�� h��/�(l0�g��`Rp���'�R�0�	�4�	H�ӄ����EO(�!t� �kgޔ*pd�yy"�'�b�|2T����PIO�s�|�B��++x�D"���\y��'���'r�OD�ꧼ?A$"A�'0�}#�$ݯQ\��4%K=�?q�����O����OJX�D���Ӌs�:�щ�	&[d���Ƞ(�P`��ş��	fy�'�~�'�?���?�2�:��!��E�|���s����$�O<���O���U8O8���<ɝOZƕ���:+T����Y&�������Onyl��`��՟��ɓ��d��^�Ӏ�O
�ccEȑg�
���O�d�Em�	Kyb��)��*��-	W/F�P�}�5�'bc|�����O����O���'�	�o8��&\	�����X
J� ��	u�������'<��d�T�XX1g�ĩ^���`4�f�J\o�ߟV���Işt��OJ��?q�'�l5Qfa�X����2��P'>����?�-O�!�6�	�O����O�i�sA�w��$�uK���l�P �O���O=�'��I۟D�'��Ӕ4�lq�@oݡr`�Q�G��[��	#����_y"�'G�\�8�T���!"[dhؓ��3(�%�>�*O���<���?���²e���rj��pa�L�-�U(#��<9/O����O���<��Q�?(&Kk��@�' .z�����O"��?!*O ���OB��ܕO��ė u��D��. �A(>5��C�^"�'���'
�U��0���jމ�rkP)d]�D-lX򉉑cD��D�O�ʓ�?i���?ё�m��>O\�ƮE;u^t���B�Y1d�K��'���'*�	�p��D��O���_�GQ��&��7\ф�h�@�8~p�˓�?���?qBe��<�H>i�O�\���A�>"V�����, L��#�����O�=m����	ߟ �	��䆣>L����/BE�Y�f�V/hB���O���9d���OJ��Ol8Q���O0o�Ȉj7j#[������?!�i���'x��'�b������	��Q�9v��ɑ)Ԇe}x�D3`��L�*�cSN�ɀ�7/c�!f��3^.d��i-b�'�r�'�������O$�Iht]��,�%WvXZׇۿz[��d�<Y�V,�ٹK~J��?q��]����F�9��L��k�2G�Ji����?�u��'b�'��'c����R�n]� �ͽO�J�X�U�(r��"��ڟ���,�O\%���OH$U�G�e��<�����'���':�'���'��Ӆd@3'D2��b#W�S�~��!�XIrT�,�	ʟ���Q��=�z�c��;&̍�Q��+����E�SOy�'v��|�'w��Ѧ�~"$M%c�¼���i��1@�
���O���O���t�&>s�űbl�!+7F
�1�؁�HOڟ��Iv�	ڟ���6
V�d��h~"$U  ��d�˰+R��b�/�?���?�*O���H��4�	�)�d�GO��v�F4ɠɓ�m��H'�0���`�����p&�L�'��$�P��D�����@���	Ry�'�d6M�|����?�S��C3KF"U�l"H��K'����Of��Ov b�3Or�OFb>�{#͗���]��UrP�YSc��Ov�������h������N<��]`:9�ō� �dPg���u��a8��@��4�������O��	�v�n��Q���ACN��@0&7��O��D�O�d��។�I�<�$�A�#��l�Pe� �R=ze����'�P�p���'\B�'��nF�X�s���%��	�� '���'/2D<�$�O��D*��k2��Y�(�G��B2%��r���t�@�����$�O��d�O��o ݚ�a"`��P�i,�ܴ����'��|��'�� �cZ�9��k��V��}����8b�
9B�'��ӟ��	ş�&?i1�'Wz�Y)�[*p�hl�� �W�,e�'���'�'���'��	�'T��F']v��r��l�P�"X�t�I矤��`����'8=���l�����z�&´������?qO>����?��ŗ�<a�Ozp:�G��Ь+rj&!d�b��' ��'�����I|j��?	 -ʧ3L8���OG {���6���?q��@3��"������k����z��RS� ��0cS��?Q(O&�$̦��On2�'	f�H����'P!�
e�����DA�'<�ğ��?��Py��Y� 4��s�w:q@��'�R.sӰ���O����Oh&��S���c��1q�	zZ�D�b�<�����Oar	X��������+97ș�E��2F��'��	ΟP�I��h�'YB4O�0�]�[�^�)�,ۏ$M�T�,�i���$���O��D�O�h�dDPj`)�E�J;Y��8`��O��O>��'�O�Ҕ�w�<n�"�:�F�9U$ɓ�c�<Yc������?���?����tE3�d1�'��-^�-2aaO�?�+Op�d�O��,�D�O�#Pf��/�=�V)9'D�N������o�Iʟ8�I埠��j�?�|I��,��Q�&@X�mK�$xv�'�R�'�b�|B�'��	� -@8�Q� ΜH�V���MYl�Z��y��'���'��ON0�'�?�Q��l#��'ɞPgxEg��?����?�b� �1O� ��)#Aȧ|)��)w�˩p�0����',�'���'@�'(2�'��'x���&��F�ġH�c˒�(��|��'��%C��"<ISe�;ki�}�JF�c�t���P
��F5�x(�vAC�D&���$=et�����ug쒅���
�wd�1\� ��ç�y��OD��~�fl���?���?����<MtZ�b��(Ad�I��_\(�˓�?�7�6x|���ҟP���1�uG(=c_3̵#��Q�uR:i�l��N��mp�'[�F�F��Bq��J�mJ�����U��Q�R��S��1!V�K.�m:�v�M����h��ɣi��`��@ܱQu�0��޾n�lԫ5ʃ�Oa�*���Q�ƽ�'IC�@�TDI�7��D듏A(��e #��J�̈ (C���t`��R�ְ��N�����L �����f�|���C�-��0⫆0���HB�,u(�|�!ՕI����R�Ɠ��$�V�3TM���H,.���'��V��
�l��,Y<Jdl��ℱAN�D�j�@y�G�L/Mg��z�&ӟ�'�ħZ�L��[X�bw�H�	g��'_��1*3 m���PAQ?��D
�$��!�"�?k�N-�&�>	��ߟ��Iy~J~��Op�"��]+��	I�7+�=��"O�F��0��I:b�L�b���������R�aؼ7&�Z!/E!;ϸ����O����O�8���Ϧ�������Ty»i)��$�ϣ?���ˆ��#i�$�G�0���-v����!�]v�3�I�P�D��0�؁f���p�[/f6�vj�>a���T�:����}b�^�<��
����`�f�[F��Z"��I���G{�;�|���H�K��I��ާN����ȓqp�#�˟.��e���Q!P���!����dK'�p�q䒢�8���N�>I�2OG���I̟���Pyb�'!�9��%)4E��F�+W4�B�x'��"%(�ʀ�X9{԰�z��(<O�kNբKZ��*'M%^�`��P� h�Uc�V�qQ)<O.d�U��UU�8J��q��"N�s����?)���4ғ���CH�I#�9!JR�k.�ȓj�Ѳ)�^�Ű���UJf��OD��'R�	����ߴ�?����M��W�\��-�*�ҕ�$ŝ1����0��ğ@���Y�H'���� ����+�� ���hZn��L s�B�iG�(AoH��I�`e�硎�j��c��b���� �OB�D[_���:s�� ��'�>�!e̓�%[8���ɟ�?E�$�ƆQ.�q�gJ.@�3$m9R���B�)�'>��ֿi,�ةD-u^�kc�>S����ª<Q�I�'z���'\2����'b�FCS�nct��Z��j|��(�.4��dU�wCn�S�Jm��u�#g�%\���O4�O��*�J��	� �#A*<�邭OD���.QӢFL�Q۬�m�"��T'		 ��@��`D{�jӳ��k`��@��Y����%�OLn���M����䧨�޴P{|�1bТ.��=!��=`;�
5�'H��'�a{����iF��\��v%+pc\���O Pmڜ�M3��Dj���T=ab�e�B$�%��6N�
�Ii؟C�F�X�6 �"l��d�X�=D�0�EiR�掍����?+��T�ڀ]�8��xU�ć�T�6B��<f|������C�I�h�s�΅LnC`-	�!�$C��>�r�8�eI�Qӂ��D�5.�C�	>
g�a;��wp�Y��-�6S�C���[����]whm�'���B�I�-�jE:�J�Q��h��Z5q�B��$Q\�X锇 lqRQ�s�V�V�B�	.40�Sb�X:8�8i�4G�$C��<W��|��iA8!e�mƼU;�B�	�n}�c�N!I^��c/Ć5[�C�ɔrm���&'p�%�1	P�C䉓=&��ZaJ�O���"_���B�	aj�I	 �Kq� m��F�+"�B�I� u����3�<��s��01�C�+,r\L�g�ҷ3 -��'��8B�	�I 
L�S��j��DP���C�ɿ7X�aʔ���Y(e$یs�C�	3}�=��D�
-�bѱS 
�> xC䉿)���1v�V9~�6 h�K�%ZC��^l�$�Û><���WĊx<C�-q˘xb�b��;�ԉ�Jãg�C��>pرP�L+��9ᎇ3MH$B��"(�h�O�9C	u��S�A%B�I�t����&��K��(��F�*��C�)� �1�F9 x��r�9B��Lo"O��*�R�h�4yz'��L�UQ�"Or	T(M�hV��G�G����"O��2�O��  (��hF�r4�1#"O�(
�۽E���Q&g�%	g\��"OZD���Ҙ1��uEɖF�t�"�"O�0`�ٛ,8H��I�{�D��e"O����Һ�|	`Ş�G�<��"O�x��ĉ8sv������� "ON�d�0-��C�J�p��q��"O�y`�L1"��``�HU��� ��"O~��E@`��Z���fl���"O*�R���y�H<0�LMZ�x�e"O�����D���S2��kJ�q2"O|���h>x�T O�$6x�B"O�}Z�e��y��g��-q ��*6"O$$�!jذ_��T�� J�}���"O��R���(-ih1���Ӏp5�7"O��hu/^m��Yɂ�@�h��paw"O���L��h�p
K
îb�"O�CG�Z�n���ٳ�N�ZB��"O���6�`��ÉS-oH��!�"O�I����!WKа��"�&J
@z6"O����A��K�~�IǢ�>:"hH�"Oب�gM�}��� �	\����"O��`'��SO�9�Ot�T"O8��R:D#���b�pZ�"O����� �2��M]�M��"O�Q#�%���(�Û�#���%D��  Ўр��ïڗ{�fa�L6D�x��fW��V�����l��)�D 5D�H�2�.x�\���ꚩ6�Q�'1D���w�-@���w�_�-L�"�/D�D���O���C�T�TIE�8D�<�!<�����RR����l=D�� ��ًc�^@jqm�o���`s�:D��;��"�Ɓ�a�t7Tݚw-$����lC7m"���&��u����A<�y��1:�E�#�(j��p�c��y��êƆ��!T'j��������y2���$��H�C*�Q��8�t��yBM��(v�0����-AX���Ǣ@�y���2*�<Pw�S� ��h������'~��`���w8�H�W���4<2�Z1 ɺ�C� �O�	�F�]�֤Ȣ��n�vԚC+�P�$ȵ,�
��?a��B�����c�|K6�~�'͸QPP"��M�T��C�)�|���Sg��z��q�Dk��5�!�M�|�xE2��H�n�@�"��?3�rΗ�r�� �ƮT!+���#���9_npсO"�
��$[�o�Z�<�0d۟n�X��$ E��$d¿�B�2�&��
�@�'C �1��0m�QqA\>c�D�e'bP;e
%7��J!"�bS^�z6bFu؞ g�*Q�V��%ǔ"�����Dγyb$T�KIRbPR�?XM���C^>@�2�JxB��RBGY<3�������-J�i׈_�eh�ŉ��N�'brȡgߔ!� �#D�^�6����'Ht����&�'<`�8���]�N%�Xc�`��/k�|�S&�K%�ݨ4"5
��ڒ�O��(��|�f�°7��!2��L�xy��EJ҇m4.K��_ ܈�'�[�"u�^w�ڠ��(Ć1����ϿC#��v���v
R9]P�c����6f]R�[�n�.�땁8p����O��p�?9F�[�ݮ�25	��v�U��Ϸg�uCЍ
�blF�a��uzTǺ?qoڨJ�v�K�[�A}�5�0��$R��c"O!p!�se�ga�'U��B�b�#t'�G|�X�x�2�KC�Ĺel� Q�n[�K_�[N	`��Ȟ_��u�i�z���J��$�3k�<��� ��V�}��j��A�=Q8�w��t�8���Ǉ/�阊�P�+T6�J�&� s� �5$��-� �ݔ���٦�:�4���A*Fr�c��jT�q�@�M�@�"��?3̆��e_�	8��[V�H%���m�.�a�	ٍeT�Dz�+AJ��i� ��R���@F��%�4�t�'+����Qigf�9iY`���=C�Ј9s�ٔsj��ƅ@�5�c$�M�0��->�l��)e��b�7
��\ySC�$I�Z�P�i� E�V�W�.`z���e��Re(����taS#U$N�X� j���U�۰\C(��l��9*T�zM�3��#>Y��M�7���'�lۄ�9@Oެ����r��-MB,��6Mɚ ���J�*)���DD��j՚�i~ݭʲ��6�6�`j�4%i�����"L�p�@&*��i���˅6A�Y�Nɓ�D��ӕDָp�Y�	��*@kȭj��9x�DޓB\l���٬��Ȃ�K��fO�-a!$���:P۟�D�#,4�IV'r���4�Ȋ���rWG��o 6-�B�� aQ�ѶS��0��m�O�.�S�Es�O!`w)�"�"��	�2�	�dʃG�5B )��-���9��0L����H� ��=����I!��8���+^�����)��~؆�I��ΣL0��UH�e��
^�!t�ʣ��FyZc{�]��Ѱ@�P���)ӈ�������;�g�:���ՠ��a�1���Z��!H	.S<i:6�ށ,��4�5��Oy�I�~�4ˢ�WDy��">�<E�C
\3U�3�W���O��R�'��*y@��S� A{��:ԤN+At!1!Ǉ�!�:����UɎ��`��8�N[�����O>u� ��hՄ�b�5m�f)dQ�@�Lאzܪa;%�'��d��l��i�v�O�&`��۽.�Q�)|di*(�	9n<�;�b[��t�$%O�OϾ2 �(��89����xj�mа�D	U牉�?���ϥb�93�4����2�iTY�g^��!&Ȗ�>W*m�v"Op����>h�(��G�gRAc�S��QÄ��<'��$��S5? ��(�Z������-�ڰ��J�Pf��Eg"D�؛����{��%IŔG%�ᛲ �dE�E ����- O�i�qjEz�\�b� �����O�a�Q�R6-��pS�㕟_��1Ƨ�c1*m�
�'�ȉ#�i�yM4�,!c�=��']0%����xrf1
�H8��k�'�@�4��I��e�g'E����#�'���F@�m�&�kp�%Ӣ<R	�'6�D[���@��aq�I/�u��OrB�O;wJx����S�ȬBt�Y�𣴦-P�|���`�JyPŦ�&8�D���9�1�ՁB�s��E�ȓ~^��cE��9\E:�ÙID�Gx"Ɉ�c�����JF)6񟰬��g.?�f|�DIɜ���"O��(�DCP�=�FR�:V ����\�AE�9`���!Bm �S��y`O1J�F���Q"/��A�I҇�yE[S�Z�F�:!�$���`޽�yRU�o(��sR/
�y2I]�&���� %�Ȍ��(=�0>���A�����7@�ٰ��D�n����uEɻB: Ic�'��4�#�5x`��[@��k�i��d� ǚ�	��W�i���?K�NS%i���#B�O`b�[��7D�\ж�ڢZ%$��Ę'�Z��M^o����Ӛ^G�ѕ����ď�Q����D�{�h�jf��T�!�dX�G\,
�-��d�r��@f�~���E"ߜsF��f4���P*1�p�1E�Z�2��P�cH��|�Y[5*��
̩R�^䲣J�RJ���!K�,��"���.:�f�"~�a��v#,; ��aܓo�zDz� 0R|+哝S�R/�>,�9	a*Q�8��D\!w�(i���?�O Բ`�P�6���A2툑r�����'I�	"OP;�D�I$PHdж�%c|��X��V�-�B��
):H($�Q%��R�
+Z�b������*!�|� �S/+Ńg��	�N���:� B�>Rc8�"+2i'�12�Be�`�s�(�[�O��D��O�y���r�n� �x`0��4"O�`HP(^I���n����5��i �{�)� {e�%��	�.m��3�^�w��Uz���<<u����:I�N��'G�?QGƖj��������RoXa�tML�<�w�¸P7�mJe�K9s��5L�L�{�t-����3	�F�}�V���B�e螶Dgtl��ÏM�<y�R�^L��A/P1e݀);��=.ӥޟ��I#�H���	aT�)p� vy(� ��^Y�B䉵Y�"�x��U�R�`�S�}~b���uhTQ%� �O*X��J�;h�,`�N�3o�1ˀ�'��Qhs�F?�$F}\�d@R0h�T���fY�<�ǉ�'l5���,��2i�s҄�L}��5f���Y��'��pS@B��x,�4���	�D�p�O�">���J"3qT"!�P�y{J@�Q�$D�胲]~P���!}.��j� �[/H�w�ǋ�����ԊSf(X��
�7m`�e����y
� �c�NJY�a��L��	`�i��A;5����4�<�p�S��y�C�op���&�/e�,�K�*� �y╓i ���n�>\�<�BO*�y�B�>٣���&~�y���91� ,[�طZ� �X����0>�W�F ::xV�欸�p#�q�h`�O�d��	�'u��H�n,�L��ɖtR2U2��
'I,& �F��\�?E��/R�ʰzT�Y"�L�@7n9D���DS�7Z}iC�V&i�j#�gJ-O$���T�22`m�����:��|ۓ)B�_B�%��Q�l0!�d�%f�IQ�-�A&(Z��C�$���e(b!w����d$�R9`�F]�DȰ�
�9�|2��z%h�0CI)Z����W
{���D@:�t0��S�,l���5��YZG�[�D�=Fz��l��q��?��[�o7�"��FHY ��B�	)fp6�X�!��nX*�q��[�/�B�	2��p�1KׄP2d��(c�C�I���sO��q�WD��L>�C��ڰ)��Ǒ�N�d}�ǉ�;YE�B�I<I�۱!ߨv,"�*7\ C�I!|�(Y��T/1�-R��@�0`C�`�����Ƒ|��˖e�t��B䉞b/6�� # �v/d��\�QhhB�I$$����g�`=fĘ6&��!�6C�Ů���"��<�(k��3��B��	�.��U��9�D-��S�&���DG�4�)����*��I�KX!�d�h���/�5
�p�y�m��>N!��*hwz����I6_�$�
�b!���
}S�M����0S"�i#h�3$!��t�Ҩ���H�IPp4%��D�!�$^&O�
����3B@T*��/G�!�үRQ��0c�\&L6i�ЏR8�!��C�bh`��s�ԽNLA1�B3�!�$M�`��  &� ����@��5s�!�$��S�N�;2��(B���c�k| !��ƣCސH�¤DO��	�1�A�e!�D͋~�
1˷z�*)ԫ�Hj!�dK2l���?`@��@dն�!��49�Z�댭zbv4zQE�R�!��-(�� �j�}h��i- �!���X�hقpcQ��!�	��!�� S�:��t+�)9��K��/Q�!�ۃt��S1(�	�δ�g��qy!�R�&у�	�<�
�9�/��8X�TX����:��ܱ�J1|Oy#!�8vq\U� (��"O�"O4�¡?V�
����&y3*Ѣ�"O��Ec��?���T73�U�F"O�P"�� <2��4f��X&�=�"Oગ��r���8S囐s���W"OP� �&A�w�h� ����@D"O�y�3h�'b~%(&n��v��(`"O����-=\�K��ʌ=�h-�2"O�\�,>�Ʃj����42�0v"Ox� Q��l%c���,�8�G"O�\��/öN����p�ˡ�R)��"O ��1�_'4���S�T��]Q"O*�a�2WdàD�c3��r"O��+�,�kp�,@�ѮH)��ڴ"OB� F�J��H��O��>ވB�"O�]�զsU�X爛E��XF"O>Ђ`"�!dP�s���d�ˤ"O%�B	�#tm@����/R��*'"OQh����`l ����K�7�iG"O䝃����^h�])#�����"O� JY ���&\�Vcُ>p�,X�"O< �!aSX��0�O�)q֤+�"O����W�8���K�)V�M$4A	�"O��b΅G�:̂&H l�x�A"OȣPK�	�ޕ��g�]��"OlD;�j�5�����ņ�'��#�"O��A��@�	BZ�gDh�"O����5N+Di*�@

kIFP�5"O�͂�k�&mʘqǖD;Ɲ(�"O��y1�T�l˄ �7UZ�Xz�"O�[�OU�k<� 1 B�7Z,<�s"O -�H�.�� A�Β/QHHa�"O�hF$�S�i5��:aHT�Y�"O�a�G��RN�!��,L�nC4)r"O���M�v�\�)r�!YZ�"O��3ri�	mٲ,;��dԙ9�"O���V�{R��ah kj�zu"O|�1�(�_��I�'��:&D8�s"O As��-:�2�F�xF�d"O�=��Ea�-y��D]9p*A"Oځ�t�@��&��'�Z�R@���"O.�iC�BO�0�R`OR��L�F"O����a̔c��� �9�E)"O(�qf`�*I�ZW�P�A�'�!�$�p��Rm���v�zgnC�!�D�' ��ٲf@G�A���״�!�T�EL�Y�A� L��<��#�J�!�ܜV;�YR�6r������-�!��-� �!��Pj�噣/� ?!�DV.kR �0b�V��Ä��e�!�I��n���N���f��E�7"OJ��a�	 Q[~5��c����Y�"O���s��_�^,S�h��S�"OָR�M71�l�h�G�伹�"OfB�`ۙD"� ����I������i��	�M%��;'@;y���#j@�"+C�	�I-�%��G(,���8��ʿ+��q�`J 	���ӝ&�y�MŖ)V�8�M;%(ax��
i"�l�=����9��L���!��FM�<90➢���r4"ДO��sӯ�I~bhE�-?�T�=E��@H�U���T:U������6�y§�V�,E	0�ܚM�t�0CN0��'S�Uء'9O<	�g /���P��Z�y�"O�0k��&7�lPh�	�?��C"O���2�̴.��y��� �z�"O����;.�b��o���a��"OF�"0�ʟ'!Vi�5�ߓ?�z�+�"O��GB�u84�W+�.��HД"OL�+�Gˊ3�X���ɔ�%}A �"O���	� �d�	���>ej�D��"Od,j�NJ2~��Q�t��d+�5Z�"OLi ��Q"vH��b<�ꅨ�"O�4k'-Ҽ\|�@�7�S"l�q��"O����	!��ҡY�9g*�z�W���ON���L%��|:��V�pj���.bEV䑥�Zx�䒣X�P�#@0v����AA���+gGe4%!����'݈���.�W�<8h��:Жg�')Bt �K֊ �^���~�B��<U��ٓmEG�H+���!�d��T��}QƑ𬝔RkN��$[hY�e+A�ɪ[9H'��Pq�!��h9Zs'�c)`�(��d)E�ي�8
�/���n,x	���@aZw�n�sE��+~C�	5�h���gY�)K���A?���,p8� JQ"$�p,���854R�l#�D(H��	�!�H�S�X�>��c1VX�����[���d\�2N�\H� ��/m򁪀hٍ8��9H�$��z-r���`ɭF�r玣t���*�����j̓M�䨨�S�@���h� ��O��Fy�f��-?d���K� FL�j���+���G�j�? �1�Q�\�-5���E�����p��X��$�VL��ș8D�'^�-ʶ,.^+z���'��'�(@��B�ᳮϻ/�R��v��2T�,,Ȳ$�z���/��O��)B��j�\%*��6`I,�h2B˒H�9�"O|@���[������L[k���9>�kR��L��aȶ�I�f�|A���K�5��!�LY61+Єg�Q�nҒ'�`83�D1��,�vi+�O�Z���&
sBL��yE@���bY�A8�dcwM�
�8=�U 8�?��[6W�a�ă�3�����jIA�W��p�)��e��H��
����Dz"c��1�8傒Nɂ8�%hb�_�!rv����B�\s��L5AEܰ�����r�Z�)�ƕG��UP��I�Zx��I/=V04��舽2o�	�ǡ�4U�&�[�;M�(�*��zMP�bZ}�05�����r���é�i&牫,��س'f�f�q+&*�D�$B�~��9d& ^�\;�JԠ)X��Q-V��2 S�ǥ#������.>���$e�z]8�F̐h��睜$Vr5�V�&�r����
Nv���6.���Jd)�$7*P8� E�"@0Y��X$��H3r�
��y"
�%��B��c��Q;�U���'�to�&��$��I�-/O�@����-Snl�ֈ�4�ȳ��9h^x�C3AL�!���%��$v�xHx��ܞ?j�E�
ڿr<M`ӄ7|O&�h@/:L��T$Õ � �j�6Od��HV�,��]
� P�v�&�j�'���P,ӵ@H�4��Id��VJ�h��ԡy`,xC2"O�ͣ ��o5�x@́{��"�K�J�zA�R�a��eN�}?�O�^ w�%w���;/<��,�H��iYf(�@l��IPۼ�
0�œ/ !�e�A h�z1�����剹F����R*R�DAi�,�+r�<���I�
l����%#�1�K�e�'�M)��Z;����w��E��:֭С*��z#%Y�1�6�x��V�܍wҒ���	Cl��ɢ�B�`-2��Ѧ�;"�&˓J)����GV�>o�q� � �p������ʧJ�X�����!Kj↟9Ԗ��ȓl'~���7f�h�J�IԮ]�r�9 n�p!B�������3W�\��'�8q(�+�)	p�:QΪ<��'�8�X�/�2�����Y�O�I�ĝ>a�ˑl
!��[Q����88�&,ÃkJ�h#���A�4\O���'�h�H��LZ�lЛ�[�f�����"| ��1��ya2�1Vq���,�>a��lD�AިOja� L����Dh��4�܌� d�0[�T�b��)�y��/ REj������@��kC���$B�$l4r"��S��R�Y�fЙy ��"��B�F{�C�	�k�������N�����ɕ>�rC�ɦ/��A! /M&m1�� �đ�hMB䉎R4�[S�G5a����%�;��B�	O֜P0�ʇ���r� �(�~���TE70X�f�-|��Ar�G�A�P�Z�j�
32!�d^��:,���O� T�)pI�>X���˷�V�{�"|��	��)��-Z$��)/��rU��i�<1���q/"��4B[?D	��\�<Yw"�O+���<E�D�Ջ'߄Ԍ�z� u���yr�ԡT�,$��,;hq�!�.�6���Xr��i��'ꡒ$���W�AOI�&�nXY�F?����&	(41���G_��s��%�xY��Vm���T�Jk��d��H�@.D|B�L���|i��TG�5B"*�e��9� ���R!�D�/T�#�NM�gX��6j	�G>!�$ԑ^��5���\7sI�ً�I
�L8!��U�KŐ\�t�E�W2�4����)0(!��	�q��� ��N������!�$�jH~]����. ÆF�%!��4'�5��a�F�X�a���m!�d�5L����� i��mMH!�䉙GK$4���� ��� u�!��E[b��y��G Ul���BA�8�!�D�9��\2È��CR�3���"z�!��r �:b��9+�����%%�ay������󄅲]�Xفd�Ŷh���sΔy�!�ہ��@�����Α�A��x��'/d�c��9�)��$LI������,G"5�0%Ն_|�B䉹v+�����N�1�Ͱ��
U�b����C��0<�!��M����0/�-d�8ЖşWH<a3'�Yx���b쑤,j,����+9 Ri�O� �d�cƀ�������)H��Y`7�'��ū�{R�7�R� �<��<�֤�(�y�A��m~���)��\�y�I�=�P �v�ɚx����rɜ��y¤�4�i�@Q�5R�� ��y�dH��^��+Ҽw�lK�F���y"��6o��I[�葉u���(ш��y��||�`�"o�hQXX��B�?��>��A�,{��cO̿j��� ��?��"�J�$C!�DO;�l{'�X*0���,M$��Hb!'�t�����	ڪ\�,͓A���K��T��!�D\���`gɎ�9�B�u�,L��"B�<�1��\j��s�J���K��zu�Y�-�&0�d�D"O�XE�5pu~���� �R�S�R���s�M�D�P�'7t������$"�䝴;�R�1	�?�B�q�Cm��8�7i;6�$ 1���2��|
�O�	�'f�,@TyQ�
�e_hP��"Oа��JCW���`Un���"O,�yE���:�
�P@(��'ZP��T"Oj���'��aEN�I�� I����"O��3sG��M3L���0xȨ"OL�1u��5�E[�W�k�ru�"OBix�)���@KJ�Y� ��"O��b2G�r��L9�/��l� �z�"O� C�U�Q����%�!~@���"O�%�E��Xn��7B��`c�e(�"O�P)�+Y�mN��"���(�"O�A�&�]���`�`��S�*m[�"O�h�@�&���#M� >���q�"O����H���leR�AV�)τ|R&"O�8D��UF}�r���jPr"O1��+L�N%D�7��F��m�@"O�TZ��4�8Xc@o�5�r]�4"O�p`(�]	@ӣL��Y`���`"O���٣^HH!�J�:7�X\Bb"O2p�hֹpx� ���0u�\3�"O�1�䬀�7lߠ.46��"O�A��.�@�R����P8�- �"OpIq��x�ܻ���{���"O��ʒ�]�_�L�c�gָ�D"Olp���]�O����f�TB]�hA�"Of=Ʃ��s�д��-��6�P"O6�P���
a�Q��&S	c�����"OLq��9s*{�E��Eg�T27"O� ���O J-�M�N�p4"O��XR��9� ݻ���%d.�M�"O��RG���,����J� � p"O\�*�1'f�9k�?��i��"O|s��˲�4(�Uo�&e��B�"O�����W�9®M� �C�e��"ODف$�?X�T��ĮԖ�ԣF"O�=�W(��t�2U@ݽW8=KQ"O iaq��4nd��n\ �+�"O�N��G�.�v㈾[���S"O���j�sL��9��4��6"O�	� �V4S�١�0�d�d"O�s���V��XB�_r��yG"O< 0�O�� ����f )�"O�q�co˾$Ҹ\bgn�$���"O�$ӳFgؕ��o��H�@�e"O�X�UE�>m��Ts��%#��u�"O��XFa�׼��ECQ
���"OXMq���="n�B�/:S��"Or�x�H�~;�M��G�O���#"O�  hz2e[�"V���>1/�R�"OX �R��6�B�;} X�Y"OX%1�"E#0칱ABT���Z#"O���P��,s^9HU�&O�����"OBqY�-���<	j��}�T�"Oh��p�.1�}���<Ja���"O"�AB�%w�4Ap�*[� "O��*���$��s���2�,�ۤ"O4ٰ��ֵ:,����\�z�	"O�����0l��|)�}�vtj'"O�1j҆.U �1�1Mݾ!�e"O28��)��pՆ�y��"O���5�L�Ƞ�h�&��"O�y���9�8	x�M�&��(@ "O>�
Q �"H(Q�W�`� ���"OFUsA�d3hh�� p��u��"O�UcNE��1���F~ �B�"O���% ɌsǪ���)D=�u��"O
� Wϙ�w�>����G� ̜("Or��gZ�SXH9��؃Q�a�2"O����ϋ	E�,���y��[�"OX,{�(�d�*�'�ĐsBr���"O��/�Ô�P��+�,�E"O�A�[U����qc݆+���r �G�<!1*N/K|�pF�S+n����~�<�FZ�:�Z���LT�
�~uc2ϟw�<���(.B:Pȳ�"F,yJ�G�l�<�VoJ� �(�B�@���Gi�<�t�;wcD��"�|b��u�k�<��*)$��5����'��(�"�j�<�3�Ή�Ȓ֫K���Ar/�j�<��$[*�ڭ�vb��_d����i�<�E�U�)�88�B7xB���b�~�<�p��$��I��
��0�hL�e o�<��ɫQݦd8Pᑂ?5�9�#
�j�<q`�At�2�$^=&}8=��Pj�<٠I�>8P�0�]!b"s�oXc�<颉�c}��ꎙg�$�Ґ�\�<) @,qv4y'��%*U��*�W�<1Qj[(J��'gJ�n%Ęc4
J�<��ŏ�x����"n�N܁$�]I�<1��IW�4�ʴ��X�h�q�nUZ�<��1[l���-�H	��	���o�<	@��"1��1HӣH.d]�����m�<I"mH�m|���B�=p�QU)�i�<i�Z�w�҅����,���k��f�<i ?E�p�(2�&E%֌�`%�a�<QV��f��L:�C���0{ �`�<�5i֚~ʺ�[�ܹ<۪H��)�]�<AE���4>��uoX�HB��9�cSV�<���R�̐�g'�+aoΑxЊN�<�FJ�����*!KW�g�r�P�K�<�EFi��IpB$$!E�D�<�b"ʮ?�d��P�,V=�c�C�<i���[)����݁Z҈��$�[�<	��]�81P�S9Q� )�7O�}�<q�CY;RN2�aG5v|��1 �y�<�׬R�n*=��Eψ*]f�锏�k�<��I�R9�L�S:P��@�e�<�#���l�� ������Tȕf�<a ���?�Ӈ� Az��'Ly�<�F�э`k� �n�6)���� ��J�<��+Y?X<H�a�*e�L�ЅˋJ�<A�])]4 2f�]5@\pc�EI�<� X(:������O� i&�aT"O^��$�7�X�a�`�-|Z$� �"Or �#�G�^dpa)��//�"O|�q��D?P(�(�C7Ms��r��'Q�d�aKҒ_��a�ܨu���S	>D�@��ܩ>���U�2qJl���=D��8��5��T��=|����%�.D��3���^���c��FP�~Z�--D�lFd](��ks�E[�d�9�5D�`�0��{& s��#�$$��4D���eD��E�6 �& o"��'D��BZ�A�x� Q�IK�!{C�"D�|s����qJ�I� M(?�tLbg�>D����
����p� �"� pԌ<D�L(B�r�L����[����a:D�(�p��BŢ<#Gm<�,C�D8D��g�_5R�R�-͹Y �M��7D�؊5��z��d�����2d4D�H�r/�!w˸͹��ݢ��8�O6D���㙢^D,�2N�p���.D��b���	[�$@��؅%7� �tD.D��j1�Ē��MBMթJ�V��'�-D��R�, ��	� �ԫ��a@��+D���HP�^�z��0� ]jq�*D�$)�!ŏb���9�*�,\��Dz�(D�h�nW�f`�5�ۼz�0���(D�A$�Ԣu�B���X���(�	'D���' o&y
EȂ�P��=;3�)D����U,s�����8\��X4�!D���9ۂl�'��Xq
�) D�x��kW sp\=r&�n,�c�=D�8��Г!�P �E(A�r���8D��Ϙ�^;�U�s�ʅd)�e��1D��"jÌ72>��K�	��mУ�:D�����D��H��A�@h�:D�t����@ |�aF�I���6D�d(m+_��1�w��t��׈ D�pڣhU-?�Zm�& ����Q��>D�09'	Z�&������3[����;D���B���91�����@U&9D�Tb���/db,C�
�#&z�q�E:D��X��׮
Y���T�^:70�Z֣7D�h�&"�6\�0)VlR�Uϼ��K7D��8���-|�1�W��rm��
5D��s�!����+��E�R�� K4D�$s��E�_���F�Z�/2 �#�3D�t�B��at�ᤁK����$D��K�+)y��D��<��Dóe?D�|��T��)S�5]Q�>D� h@b��@eby��B��P<D�4��e��pY�/ ߸���J;D���dm��Z���0#�Ayۦ�x5n#D���͑�"�$L�'-�X�n�`'D�4�@�dl���ϑ3G^-��&D��ElÈ���s�l)BTJ�b��%D��#�Q����J�F��:�d"D��{s/��Bqz]Ys�k�>��M!D�dёA ���3�a�5
(8� D�@f��%��0ID���>l�*?D�`դ	+~��A��Qe/�S �;D��I"�P-o�ژ�$K~ؤq��9D�8:�J��&>�rÊƀ!�f��T�2D�|9׊�Z��QQ��Z"^y���/D�iFj�!8,k`+Ș,8Jň@f/D�� ���Ȟ#Pnu�A� <]���#w"OnY+�eS�M�]�0�ԧd�t[�"O��8uIAq�DrUjJ=s����`"O�;桏�U-Q	��@�VŦt�V"O���b*ؐk�j�P�h�sa���"O�LH�43���!g�bi�UH�"O���"e��-i�}xuś.�����"O�DG����p�_�j*̊�"O�P�̿P��ċ#�iJ��"OX����;��t�WA��q8F"O*�ٔ� 4~H��do�G|`Cr"O��: !F�)���&�2;d2�Q"O� z�^�c� �ҕd�16U���0"O�܂QD�?8��у`"��[T����"O踊 B�cJ���`�S;ZHR#"O e"K	�pb,�R���.du�"O�!��Hy�X�P�&�g0�q&"O��W@��"�2��2��}�)�"OT����3oD���+_"���"OBu�U- >�D]��$D�HC�q�"Ob�K��N��J����#%(�a"Op%+�DI�S��y�b��0��b�"O� �qbڎj�~=��aI�	X0q{ "O�{����3��z���J�4 1&"O��2��'$������\a��"O ��ũS�����@��N�`|��"O�@�l���(��a�
F�h��"O�;0	S3oh���@n�N���%"O��s��A�5��� 'N"�,:D"O���@�F9Z�(´�
�oV�@��"O�,��3���b3�!=��aa"O�p�s�� ~$�16cB ��#u"O\T���8�&	y2�V(��8�"O"u9䅑=*ǒY9��"���4"O�h$Ӭ}����f��2��aU"Op��
γ3��%R��I�G��
"O���"�D�2���F#��7"OF%��
R��<%�c�윩�"O�\" LLb���Н9d���"O6��wg��{�v-�E3&2[�#"O�cU��T�M�e K7<t"d�'"O�T� �,8.r���@� e�)""O|�H7�T�4�X=;��"[O��"O��{�G�v��,s�� 65�jT"O��s�]�p#���*Q��l��"O0��'��ojxEZ�I�{xl�"O@� Dqap<��P��� �"O(�Гc�Xr�Tr"�-q��eR "OL������� ��dM��x�"Oځ�Q���:�J�X�߽9�H�"�"O.aq��>� �K��ٌ�h�""O>ٹNA/�D���I4Qľ�Ӏ"O��A�Tl���S�	�ML�@I�"O@A�0N	���kH�7?(��"O�ّu病y���B��y*`-�!"O�H l��~����B��R��(�"O�u�և�3W� p����P@@"O�!����L]����5�~�"r"OL̠�D�����QTʯDР�Y�"O��Uč���;��/5TĄ�G"O�R���&Y`�-@C�f60��"O�kuA#Q��/� 5"q"O��U�W�����ϝ�B>Nt�t"O�<���(4�Ը�.��U4����"O� �4z��R@�zi)U�[89��"O�E��KR�_bNZ@��0l8�"OLe�`�h �}aE�â �x���"O2��c`�|�c��[���"O�ՃeP�$'0ԡC���UJ6�!�"O�DC��C7��誥a��.�����"O�`*�/<U4$�Ѐ
�"@�\2�"O�S�CE��!K���m�p�s�"O���FJ�'Kl$�7j�+9~��c"O�dkP(MJ�4Q�P�H?��b�"O�`;FD�7O�i+�䋆&�]sA"O:p"g���'
��d��Y�:�f"OF�ے瓸)�Đ[�S�V��"O�}���^&[�(�p ޤ;�*q�U"O�lk%�δ>ab��.�a|�hҗ"O�TZ�톴6D��`6Q���sb"OX��`Z�;l�2��<v^\QӅ"Ox5��C�_*z�A#i�
[hQ��"O(f�[���7�-�
t��"O\���CM�3�(�#շb�F��t"O`�R%&�t�ؽ�rEɘ�&q��"O$�p��?�Qc�DE��t�2�"Or�I��q`B��d�ƣFtp�1�"O��1���_A�8��9@
d:�"O`�D�Ŀ$�@��W�0a�!H�"Od��a+֠D8�h@u�����sQ"O��Ȓg��^(FU��^�U��{u"OL�
̎�c�rx�@
�%�`d!�"O�}R�[}m�ɒ�)�+�8���"O^�&H#g�HU� � c�j�"OP�2p�P-!�6��ʒ�^Z���$"O�$ 18^jL�@�*��jVF�8D"Obi�s!փtA��x�I��(3�9��"O��R"#T(`ͺ��_S+(!ha"OT��
U�O ��a�'�	L���"O��cHK�8�NTb����qcZ�� "O��ɷ��]I����Oï`��+s"O����)Hp����ᎏ_�r�b�"O0�g���qF��� ˶h���"O�h�q@��`:���#�H��Qy�"O�a�0 �1��!R*�@iN��e"O��+1.�>=���ޘd��"�=D���GI��0�)���6���نO0��<!��#fbd\�a��4�p�
u�h�<i�.W%.U٥�Fj�\���_�<���D�2��l:r�͓E�\� ��Q�<�7��2H��wt���OAB�<����t��  -еm��Tk�L�Y�<�4���4�ೱŉ��(���QW�<���Z%3�T�!O�0 �	�S�<Y�̩+*�Qd���\F� ��M�<a����?�D�Y���A?��I�G�<I�/K�9¢}��	f�k�`�F�<Y��G�^B4"�.F}z��c �H�<�q�>�6E����i`-*�l�<)F��S�`�p��Cx�����M�<ɵ��'��$���ܤ_@��aw��s�<G�;��]��_6M٢�a���s�<YHͽT�f���(X�dr��� �n�<�I7��ڶh��2��Ԫ a�g�<�&*�b4��gU(=�z8�D�g�<�5/$d
��a/%=�&P����L�<�ӫعf#��0�`Z�&���ƜE�<��+�����ʧ S�]��sg��A�<� ���wϑ�E�(��5�-�"O�l)g���Z1sSg&ض=d"Oj�W�I;&R�m�ȃ�t!����"O+�
�����*:�D��*�Y�<ig��Q���F
J�<���_X�<�CIA%7��9�n�=*���1f&�S�<Y��9P�$�k���n$����BM�<92h�3C�p&�8��J�a�q�<�$�^�Os~����H�8����3�i�<��_���9bRbQ�`��(�v��b�<a�螡���c͜ZX�R0I�v�<a��ں/�|��b�"nt��R �
o�<	fh@���L�V����Dq�-�l�<A"��XgjmA��I�Z;vP���a�<�cJ�ݘ=�t�]{̠�тgT�<	b߲ ��"�@
��1�@W�<y�k {�6Ey �X%e�ܳV�[�<��"&׆�;'&��i�� �Ea�<	W��&-8��q�e�	_ .��3,�W�<��Za|yi���&��0�j�U�<�`o� {Y(`�c�G !1^0s'�[P�<���R�l(��A;J�$��&�E�<�	��0�<@�r;i�Ȳek�I�<�1�Ґ� ����
�h�2�/@p�<������PJ�m� ����Ps�<a�bǐ	��3L�o�"��@MYJ�<�-tK"iCÆ]uCly���F�<ISh	�(�l�s&?,�ܠ��/C{�<a
ң-Ox�����9LX ha u�<�%� _K���:b��P��Ɂp�<����/%\��BO2�T��PH�<ّǽ
�b���
[>�a�.�j�<i6�	q�a	T���1@�����h�<���ӫ�:�@�g\7`�e�@\e�<Y���G�<c�A3e�&�2��X�<i1H�^6�Q�#�E���ȣ��S�<�����j����Q�1PsB�M�<��M�EH2) s�;�@lp��SL�<�,HqV�=�1l֞!}�-0p%�D�<����DW@�8!d<�^��J�|�<��	N,2h<-� �D�,��C�a�<I��ްg*�����Z؊��g�<��Y�����ˊ.5��9U-[�<A�'�<�e�n�-M� %a䨗P�<�������Ğ^�^��	L�<���5,�����
�i��P�BJ�<�&�>k�"9���՝A�@�EYF�<q�'�U��(�ˮ�i"��@�<�R)��Z@�d+I�!b�jEG{�<���)D9p�FXA�! Q��w�<�,�:�`<��K�'R�B��v�<qnȇM�8	Y@,�/Yi�)B�k�v�<i��iwd���"+7�*�)�a�I�<��Ti��CWO��kr.�9���B�<a�,I�T3�-��	�2H����S	�z�<ٵ$^i�V�r&X1CL,ĒC�v�<�`�ήzK�St��1���1�g�<�#�L�>br����ѫ.��ٳ���f�<�s����
� ���Q�G��c�<!ԡ̥o��T��E!H��E��D�<�W�A8vN*��s�vCz��M�{�<qԠa���hwAƟG�*9"�f�q�<�'M�=��$��|�OZm�<�Q��q �t��J�~�`/�d�<� n���#X&~�����ro���x��'�����S�2��ٶ��3G�$1+�'o*�jń@�^m�h&MA�>?-b�O��dS��.Պ��A�YJܚэ�>C�֒>I�"~n��T���특 ^xp���"+hB��9F�6���K)��ѹu�v BB䉌!�R�@d�Y� ɬ�����-�lC�&R�*���k�(,d�L�ω�ybdC䉤]�&�g
 z���2�cD;ȀC��(-�d�� �ӳ$�\a�P䆯�NC��-AH� E�C�wE\)R�O��SeC�_ȕ�eb�H�@��(V��B��	l��@@��&�~H(�iߩlo�B�I5pm�@`4�⺉Z��ǊGtX�3�'�@�[�HL)3� �Ŋ��EQ$�A
�'�
1pNU+P�De2� @���P	�'B�Ba�8N�q��AX+=�@8
�'���h��NTN�Y��3�(�:	�'��р��;4�v��9/��ݛ�'d#�̈(th�C'E��'�h�'꾉ʥ��3N�l4b�$�K�y�'�\$�"��1#�l���E�*y�`��'��Qb�+ OѸ���ƤX"*�'�p�Xf��D�pEBa�S�~���)�'��$��[4�q�%�
 5vA��'�3�B�(q�65�WPs)d��'�~���Jٱ��iAr�{D&��'?d�h�B�)Y<�)���XB
�'�ڱ!�K�FOJ�� �)5��2�'Cz4�.J�[�L�zJJE@
�'�Ա��J�r⤨�äm'd82�'7Z�q�"U�5i��AdKK�kreC�'�����́k���hP�Ba��T+�'��@a��*K���F��4KIN�s�'����@�\�4z<�Ђ�1Mh}p	�'�������kPH��J}�Z	�'��t��ž�4A�P�8{�~�9	�'���E�D�-H"�1��v��Y�'�Ĭ��L�!`��p��##Hα�'�	S ������ץ�$(�8`��'_X�؇L�6�${���-U�dѸ	�'5�d�&�I;ے`[D�I7] ~��'�"����!V�����Y�t���'��T�oM,R���b��� ">��'�:�8�`>n"`Y���P� ��'"XL�囊5��Cc���G>9#�'ڸ� �ϣX��4pB+OB�1a
�'/
�0F݌���a!К0Z.a
�'�,㱎�.05.��䁩's�Y
�'~< Js����y*��I�i T
�'Ѣ,!a�žZ�ܪ�mNfV-:�'��%CE��V2�����3a�%��'��=�C��jfȊSHId<���'���+dLP6!�@8��
�,XQ��'ڽ�vc���3nM~]P��ŀV�<�'b��*�6�㷃P�f����L�O�<�����^Z�5���[j��p#Bu�<��W�� R�ȃ�a���E�<	���XOx5K� B�O�f�J&�V[�<Y��Bk��l�@���}��Qǡ�M�<��:z ��2�@5_EL�P �VM�<�Cg�	�pc`�K�a,��٢H�K�<)�$�>�l���� +ࢄ)���D�<�@.VM��)֤@�P1ᣀ�<� $@3��%n�n0�6(�>G&:�ڦ"O�`��B>Yb��L�	��+"O�ٚ�㏉J��<����`�6��"O^-r��Y�Bz=Zt+��`�1�"O��s�M:�<��r��=RHx�`"O�躕Ɯ:9�JݺSB��AUFk�"O�l	��ܬJ8,a3S�40����"O��*eY�� �h$R�"O�-a�F�ITƉ�C�E(NpJ�"O|�a�86���V���U$|	�"O
L�3'�6D�6��`Ο+6*��4"O|�XR�ɫc���@�m�"y\P�k�"ORRf�
V�朁glْU55��"O��"�K�W
�x;�A�1"2B�V"O"X���g��ۤBA|a"O�-�F&�0"�H�a NB> �s"OlŢ���X�H�֌�� �*f"OfT��C��'�(W��~w�8æ"O"0�c�����0�F����""O(Dy�OZPTu1L��"�e�"Ozez�%Ҵ0���ʔ��i�\�KB"Od<+sBM%�t+���'(�B��"O*���2gܐ��<Ϊ��"O�q�2E�:A$A2d(�Eg�x�"O.���сW��81���OGhd2�"O�Ȃ�g�Q<,q�Ý"`5���"OΠ�F@�$SD|��LC�$�k�"O��k���/!/�1q����4L�"O���R-J�D(�K5�ɝ�z��P"O�P�5�9av����G;����*O&ma�'�(N��0R�	,E("��'	�@� :x��'�#:9N܋�'�:Ax��ʣ,v@	��Ή~�zܸ�'+��� "��)���?t|�e��'dΑ�T�ŷ7���Z�eA��'veb�\�)v�\cU�˞d?�c�'p��Ĕ�&�}�MI[s�-�'ר�8G$W	�4�4��AԐ�I�'a�!ק�2b|��JĠ��An���'�T�:� �Zq�ӣ�_q?��S�'jtm�"�%�l��F<�Z-�	�'�yb�`� P��e���Y���X��'���ȕ�N4=(�͠�A��wbl�3�'Dɋ��4/jݩP��;c)�Ѻ�'G���Ɓ���)p@�PZaH�'��ோ�7�L�a�+I�O�|y��'�j�JM6!伔1�[�Y�P� �'/0,�w�k/<D��gI8J��5��'�d �����0x#��I�&�1�'����`#� @x�P�F����'hv��挌8�%�TdN�:��Z
�'�py�-�DX ���1�|R
�'J@����	
��F��)�*x�	�'c>U�tGݵO��FcY'x`:I��'c0�J$��5!�;f�AF+�x 	�'� `�����	FЄh��**�����'��q�Q4R�u2­E7#ހ!��'�r<��>!*Lʑ�K)�d=��'�Xz�`_[�,��A�1L ��(�'���BKc�Р���<��؂�'�� `
H���M�-��'�*\[�J¼{��<�Qˇ�*)��K�'A��p�:w���I�V1��A�'�"h�$O���d�p���h�C��� `�w�T {]�Ȓ���4a t}S"O�Q�4��B�jl�!擒6�쥨5"O�ɪ�o�.P��$�uƔT��ʢ"O8��E#Y��ܽE)C-#�0}�T"O~܃�@
3#'2��hA6l%s"O�ū���s�r��g!�=�^u�%"O�TI%]���G��9�,=7"O�q bD�v�Pr�D�:�։�"O����c�_ņ��DnF�!��ԛD"O�P*��\I]� ��}� ��"Op�0#��&�,"�-���
"O
	�����b� �:3"O"D�Q)
���B�v�����8D�l�G�DVq�X�u^�#Ɔ	e�5D�� ���G�N���,&4�VA+S�!D��'E�zpDx�q�4SkH��6�:D��0���� ��| �D�32+R8��>D�ШקϤU�p0�B��:�f���O'D�,�����������d蹀e?D���U�3ۮ=3�������F*D�L�U�S�j���Y3" p�0�ia(D�4���#[3�}�Ŧň�L1D�$D��+�"yQ �'�-JI0xTg#D�hydH	_r�
�����m6D��Aա.K�>a��m�Bi��b�1D��P�i#I��!��W>,'���$�.D� R6�*LN�)2�T6cu�LQU�+D��V�M�J�:	�6�Q�ĐS�N(D�X�2C� 2N�ۤ��A�b�s��)D����ٴ�*h#�G�1M<���#D�2��U=����P5Oؓ��&D���&hF�3��c�㙔k�L�H%D�ɢO֭k��I�F�<��pAfN'D�k�ğR�hġG"�B�@QL;D��#��w��К%ვ;�X�j�.$D�t�cE$e�B�x��b� ���� D�(A�c�*X�U����YB [6�*D�t;�;\���@�IT�p��7�,D�D[�I��R��&�C�@�&d+D�8�!��f� �QR��&,�����f$D�LJ�AYJ��0���ҩvĎy���"D�Ti`���i H"�iRX|����*"D����R��P�F�&� In D�X����9�bl����|����b?D�@���M��J��
&31n4Ҏ=D����M�S�D�����A?f\a:D�p�^��t�H,^�@� �ownC�ɩcDB4�7�
;�L�f@�-r�ZC�I�3�@��� G�M�y4*���C�I�VD�'(	X�4��`����?QߓSb݁�
y���q�I�1OV�ȓ1�Xf�ޕUݴY�,��'P�Y��^Q 4�B��:[�&�X�A$�����C\�:�.��hy�qc�L�f܇�3���a�:�d`�$F��K}x|�ȓd��)�j
/i
mR��Q�u���ȓK����
�8���c��_8�ة�ȓF��}���C�@��B��L���<qߓ!����>� PӀe��HU�ȓ8:,p�d=a��,��BcG`��ȓT����F$��_����!g��@��NQ�UJ�h3x��*� ?c,]��~a,��g!N���@�ϑ�L`�ȓ,�&�)�m
�x�����j�P��S�? 0mq�F��R������O�.2Y�"�Ĥ<���4�؅��N3>�	D
�nz��D��̅�	Zwt�yE�ֶjo2�@-R$�nC䉒�
m�2L�)PA��
;��C�	kT�Y;�HY��=���n��C�r�$9�e���p���nH!3�rC�I����h�Cd:e[f G=M4
C�ɽ<x�Q&cF�?&:�˂H�,R8�?�-O��=!��r4�y���˫(h\���prd���?��I�M}��9�䊝_�!q�`�_�<y#M����9#�i#4~�rrv�<!�G�y[�I;�%�-L�j�/u�<!�	^���"E�H%C�9�fM�<�SbیO���6�̥GV��ϓK�<�6-�=2���1f�G=/L���gF�'$�y�g�/tE���X�R��H�n[�O��$�8!]d���d �>����\,F�!�d�9EHz�S©���j�ߝ*�!��ﬠ"'%�R��e�COģ�a~�U�����߂]�J���=�	�*�f������Ÿo&��4�.L�̓�b�!�D	N�Hs��]�4ŀA��)+C�!�d�c��R�B�0p�4�@�	��!�]!w�h �5Bx��˵�~!�d��(u⦕�Zo�\�g=!�R�x�zQH�(���N�����"f\!��E<!���p��1��AБ �}H!��)�͒��:	4`SG� DL!�$��!��`A	�qBl=	'�$�!���Khj�p��Q?g���\'k(�	p���Fq:  �8]�����Ԃp^ D+�"O��2EW7\��A��1?N����"OFԺ���������z":p�g"O��c0�}�X���ܻ8���f����ɸ1|xX0aF����hw((t��B�I�B5�@�8$@b����;5��	k��������% ��@��&rFhS�����R�S�O�R�v+�*@���W�Q�F�@�'�Pj�L'e�!�]
BXz���'�ʡQ�(�5gJb$[��%+�HK�'(m�E+uAb<1&N�����'�`�l6,��95	"���q�'z��N�$,� 5�F���X��)��<I�FS�Sm�a�����L�b�A�q��hO1��]p�����|a��=>�I�R"O�	���(>j����U��I"O��R�#T�ܺq� bL��"OD�Sv�_7|~E��)йB�<`5"OĽI�E�#i��G�j����5"OҌ���F����D+�'�R�"g �I�"|�'�\,R5bAb�L-h%��3Zސ��'�Y�F W�}�Ɂ�6U����'Z-@L�/��󎔠H�!�
�'f$\:Ѩ��&F��8HAt�
�'=p�� ������Ϸ̀ݓ	�')���R��/l�Dٵg��P�(��'L<�CO7t�̄�5�^�18^|@�'"m���[�z	����$k���	���'�j6�Ȅa�����	��v���'�*L R��_
�{d]9z�ո�'ST;� C8D���9��	��]��'�a{��:�T�Т��z{-��'7ў"~Z��3`��i m'P���F��<����ӌM�����.ą������x�*B�)�  l;łB
�#N	(�
�#�"O��0���H�^]���x���"O�݊Э�)(� ��'"��@��8�P"O|�p�韞civ�y��D�o��I"O�8����+�¨�D��Sk��a�<!J>E��'2`I�σ43�U��/'�+�OL��#�)§)�Ěg�:)O ��@��!h��ȓCM����-.��-I�E�*�<؇ȓ�օE²e�����N�8&�옇ȓVy�Q�O��F�j}�cc� x�>͇�Gf(�3GT� �>�8Q∽A;� ��fe��$�2s�
؃L_8aPx�ȓHQ��`%\6���6n>]�ȓ n��Ϙ	���0��,<{�@���?Ab+�.i�x��ְ=^�TYR�<�E$�#Pčڱ�,17���vL�c�<٢קVaJ�㡋�h��p���]�<ٱb�A%��y#K�=�����Q�<)q���Mu"	�dH�,�.˥͇e�<w�2)�z,�v�ʥJH�B��k�<Q �C�FMPYj&K��D� h<���0!ADܴ:,�4$��î<��'nB����J �`���@]I�$�ȓ���sǄ�/���t�
�V6HU�ȓ���"�NИk���	֧IՇ�7lI
se�89�,@E��)��l�%隼9��X��g� V�Fx��'���H�����2
ǖ!�D�O��+#J�MN��C�?d��"O�@h7� W ���ec�?@>Xك"ODd;*M8�%�π.]�Q"O�8��I��s�m�D� ��"O����·F�Y���Ҥ:t���"OXm�5��6�H�z��ءwZƅx�(|OH �)V[����"�-:C�u�g"O��BQ��TQ����A8ZxmӃ"OD������V�6�!P$�
@ I�"OҸhc��_.��C�"�YB\A�1"O�Lp��K<�Uh0� �>:�`��"O��&�	-L�)�� �}�<��"OZR������ƅ1qW����"O�m�W��n�\BG��GkLE��"O�iW�Վ�b�zWNM2do�Ţ"Ov�?�:R"J8'��T`2�~!��X�r�c"$88�R �c�8o!�Z�E"1��"6�i�QB�N�!�D����e@�
#D$.�*%�Z�!�Ċ=K��ْ`��*A"�����@�!��^�p0B�Ip�R�S/��P��2�!��DVq���FiD2�y32�Z�1~a|b[�@��%w2���Z�C�Z��
):B��:U�:;@���8ܢ,�%.A�=� B�	��)�Wi�7x��C"��/��B䉂%�D8��'l���K�A�N��b��G{����]��0#����B�Bj�y)U0Ak�n��ET��+b�Y��ybC�&<� �8d��7f�bR��ҭ�y�NG�"�8�D&ӊknpk�͒?�ymJ�_��,��a�;:k����
�y��?L>��ڂa��
"�,C��0>�L>��O!~�pQ��P�}S��@QHK�<Y�f��1s0C��r^��f��V�<1p��+a�p�1��1\]�� ��
|�<��oe��F��4�$�H��v�<� ��3#��I�f�Дo��.��h"OФ(�,F��d)������"O<�Wʈ3drָ{�,S8p�%�f�'��'�x�#��2w"�:���"f����y��'��y�dU�t�x،T�~e���Q��y�NʠF`��"&��Ou$|���8�yү�fM����V�X�ȅS�_���'��{2,ߺ;c��aS��A.`� �*���y���~D�`Ȅ�3:�2�s��F�<Ѵ�5^pfL�pHJ�	�>ɡ�&�Y��G{r���p����m��yr(]�'���O��ĞK\mp�ț3*Q7c�L!� L��	3���\Ox+�� �Nu!��:P���V�{2��	s+�"d�0�O�p�K�d9Ε�r�X�I�DT��"O �!���o2��cɗ�@�xH�"O��0�+�dF�y��8V�����"O�T�@M�F�mC'�jD�-�d"O�@��TZ *XS��xB��"O6�;��ХPt�[t��_0�=�"O��c�&pK��X�EG/'�D鰕����	�|<
�zs!�|eh`a@F6*��C�I,�RQƖE4T�b�އ7��C䉼]Nn��f[\���s�a�C�I"+�T����C/��9Z�I�(\4BC�	�BsDT����;9�]C�+^��B��6N|�*3�X�X]�Q獇�ǤB�I6�ʽ��*{�N�RF+E[VB�	5 ��MA@#Z�!\���DEnLB䉒K2�e�P��|� �0�I��s(B�ɲ}���慕�#��F#_�(�fC��n�Xȥ+H�^9�taf*/N4C䉬#�dppw�ε�f��RH�C�%*�bCBBO<V�td���ٺ_{�B�	�@�I�g�R<��	�N�B�;a.LiX �T��z�C�VIY�B�I�Mb$��M��a\X�����)��B�	�V�����'���
��JK*E�!�ĕ�B�ĉ�V�x)��)� l!��Ւ,+��ߖf��=1�&�- 	!�$�s���!�A�L�.�柙\!��8oƼ����M�ps���X�!�$C�fl���7��%�6#w#[�!�d�q�`���&�>O����C�,=�!�$�..y^�J���_���aâǜ�!�-ʾ3G���7��1a�֓ !�$щ,<�Y;ѦPO;��@ݲf!��M%���g�L�]+��V�j�!�$_'&#Q�Qg�A�u�!�-N�!�$U�I���2Qe L}
u#d��=!��b�&��F$�XI��"s	Α]�!�D�ą� k�2E5��`��H�Z�!�d�"R��Ѝ�	#|����!G�!��V3E�8[1�	kk64a��#�!��G:Պ��ӈ(Q�@i�쟳;�!�䏬FE�aQ�ӤF2�@`�-P����2�S�O���Ƈ]�<��8p1�A(l�m��'���ʵ��OXF�QT�ؘ\8�x(�'��y�o�
,���ȝ2VM�,�'�\Qwf3V��{�MA�TЀh��'��S3hP>�.y��m�6X���'�H�c�A�*�4�+"F���b�'~v�sV�jV��"���Fsl��s�)��<�1,�Lz�� �N
U㊼���c�<� �ЪpR0�&�J4bA�p&dxE"O���c����3`��7>_����I|����5I�"vK%�J�SP�r!�d��b�Z�7��A�y�q�H0!��<C�%��n�y|�|Yä�1O!��Z�p1��d#
�0mpIS��>%�d)�S�O�-2�ΞbT8��2d�!>ޙ�'
�`��Nľ;�����̢�hH��'���W>CI0U��� &b rE �yr�)�S�:�&�h5�S�:0j�bUoR�(�XB�a��	U�S�y��v�P�Hb*B��=%A|	�aeI����XRȍ�n�4C�I��,87gʍ7��Aȥ,^�����.D�p���9�t��@-�+a� �+D�Ln�I�XQ�Mܙy��A�uJ,D��G�Q�Hߐ�BeGo����!.+��hO�4}.�S���% �3!۽F�B�	�.}��(�{<�L�$)X�4��C�I�(g��qalLlHQ9B�C�I�E���s��ʝtb��ĥ2��C��4s"�;��K$pX��W���j�C�	�LWv�CFN�Rb�z��B�-�!���o<�(��D�9S��}���;8�!�B�D��ܒ�#ū<�`�D�J�m�!��[�C��5e�,�"��W�&Dy!�D΄O�l�a���,AI	�!�s��1�c�C	0LXbaä/!�D���EId� *��rO�H�!�5�.=z�� �|r�mŷx!�F�zSl������R��5r!�G�W#xX0��bB,�h�T�Hk!�dM�gު	�a�c" ��a��!�H�'�Y+�f�*)L�+k�N;!��&�����P:����$� u%!�$�+Xx��q��31�2��g(M :!�Kg�^�!�ʐ��8�b�� 2p!�	�]�l�����>�@#��#j�!򤝳]�@4"���Vn�����L!�O=�,e�� ��Ji����@�;�!��
�x }jl�b^tM�%�Y�~!�ě(z�@�g�Ŧ#]R���LF!��7���!b�'�6d��Y�*!�_^�mxC�	nl��w��>1�!��.�~�J��*��%��Oݮ|G��F����;�H11�ӱ#�8�TE��y�K�NӀd�FF�/ۂѸt�U��y�鉹30����Y��@�'F�y���G��|�f��>���c`H�y�֣irf���$�'I� ��$׎�y��Օ���Fʌ80��	�-Q3�yR�	e�z赁�_t��(3�K�y�ǔ�Q����v��g�������y2F�)\F��#���4�F�d�ϭ�yR@Cm��@�#�WD�����ņ��yr��h���i&DJ�	���A�5�O|�=�O�$�2��ԭyN 5��&DM�u[
�'� ���ړp� c�#�?Z�}�
�',���-2t�4��L�:�	2
�'�uY��E�j_�U��l��=ˤ�	�'�% �>�|���]�l~��
�')��#�V1�Q��i��P��'u�|�u��R�V��1�H�N���'�Z�G�N�@Q�Ƃ?>��j�'ި�K�+7S�.iJ0.��:�F����� 0�(DF��2�t��7��/pC<1Z�"O�ch
�O�$H���V��"O������nŰx0�g
O6�qA"O�QvfD8���[?o/>9r"OQ������I� ��X)&�Z�"O��H��RC�U
N��"O�����a�B�R�L��YjE�4"Ot�����D6$��T4����'��'��	R&�l�@��pKD�4��3�"O�E{�A��!Ć����
,�I�T"O��!����Eꦫ]�d�j�C�"O���猜�
D٣ቶ<���"OV���]�D)�����B�p�"O�����6�r��������7"O��SWςn9�e@Cn��4���C��'	bP��r��Ƕm�:h��ǆ�r���Qd� D�x�vM��m�t�	�	E��D1pf9D���DJ
9{ݬ��%ױѾTAB:D��suG]ml�B_ 5�ڴ�ve6D��iw��1���]7��t�2k5D�$aV���Gt̐��3H�(��0D�d9R�̽	���Z"e�,�|��.LO�㟤���2*�nݛ��F2�0E)D����B̭!����!�<���&<D����oЅ̌E!���/X���@�H<D���R�	M/t(J�'�!q�A��,<D��і�	�:�lը��[�/��aP�k9D�ġ�	խNK2��a�Y�u�DQ��e=D� 1�-b�:�1Lւ@$
���6D��I�kH8`��jArR59b0D��Г�HK�e(���y�Ĉ9ǋ.D�C���&WrL��e֝x�j]�T?T�x��!��(�P�``��/Q����7"OM��GڸK(8�Y���hl.(#�"OP�F�Y�*��adSw6��"O�ݹt�
N��h�m�j��P�'��'},%�E+DF�H�!�}0��'����7L��e�`��{E֥p�'���H�0�ڭ���Z{b�`��';�PZ�!�0Ug�dQ%R�r�
@�'`��a!���H� &FF+@�!Z�'���FOځ���J�ޝ��'ɐ�$N�.�D�[ŋťA�����$ܽiՔ1Q��*&H�cq�ܧD�!�ĝ�c}������{D� ����~!�T�Da�u��}��*��]Ks!��a���7���		�lV!�D_�x��s�V�o�#�-�!�$M�����*Z�3�R����J�%�!�䚝��P�r��� ��a|B�|"m]?�1#"��^>�@�(�y�B��=(!	�����
.Ʀ�y��׃<G�E�`ĝ�]42x�� �<�y�䚻u�0@�B+�U1����L��y"Κ~��JW�M
Q���Aw�0�y�"�Sll���
XN/^�0���7�y�@��a�ȼ���Y[dq�5͚ �0?i-OmcfL}Dfx�El^%2���z�"O����	G5~ML2���.I�H̙"O��KY! ᲍�7���/��$ig"O�,	c��qخ!cp��� ��"O4I��n�L���B�]�[W���"O�[r(׋EV��1r���`m��Q0"O.���%g���R-�$(R� �7O��� �E�E
2����E���Mi��:R"O&S��	��%aq��g�I�"O6U��L*8��haw�14_��!"O�ԉq�E���a�աο)(l��W�'���uy�석�YR�D��V�E�0j��y",��vb,a��`���X�(@�V��yrbMi��͐�j�h�J	��ykҐ1��h�G���@�V톚�yBo+e��u��@
{j� �C���y2�C� dT���;�`8�s�͒�y�E�B6�� ����0�v*B��yb*:@����!���2H�U�W��y�A̼ "��P~-֭�rʋ=�y"����hZ#�7)Pd��&���yb�\�mf�0SFY�O:j�H�8s��$�Ѳ�����9^��-z",^B�!�d�9�PI�'
L9@\�(Ƌ�(E�!�d<xj8��q.��E&�C�j���!�ӜdF�I% F���m3��+�!�ĉ�5h��Y��Jvɮ�����!�M�\��4 0(P�)���}�!�ʣ7T���D�X�*�"'�-u��$�Of�G�=I9�e���_"JЀ�"O�@��*�r^Vt�:�ޕ�%"OΨ`�
�6C��KWqa���3r�!���C����Μ�B"µb��!򤄶*�j�)$��1[)Y !��n�!�$�5U~p������X�t��� �!��#3�|:�I���Z���e����|��+y���* &z%���.��/�8C�	
��0�D���|�5�F���C�I�B>t4�"�U�#^�%���B��`B��*%�S�NtmT��-�&*SpB�ɸu����L<Zw���@��T5�B䉡[e���v�S*��()]�4B�I�t����\?.`��9�%� b����(���r��->�Q�H̔f�B�I4d�qѡi�Uu��i(]ajb����	�^О��փA�-��	�ďޤf��C�IH����Bo� #�����l*�C�����񣪖�h��c�iXBxJC�8/����+�:q�L� �׏'�&C�	�g�᠃#úE�f���	XZ]c���>�詁I�[���rT�U'/�џL�?E���'\��1�S�J) ���7GӬy�'x�Q�t�X�Qnĸ��G&tUgO��23`�` ���A�%���'"O��q �[�BaDHZS���9��"O��@�P�~���2&���:R\�j@"O�iN7>K���W��1�"O�=�!�>X�̠:�Ǎz���e��lE{��I�"_g|�����e���ѮƣD\�7ړ�hO\��r^�7z '�ʒ;m����"O��؅��8��rI	6i��;�"O򭢴*�*:��,ӂ��_�J�"O�i b�S�J���b�U/_Y}��"O��1e`Q
�p�D@4O
dS"O��oY!�~�@d�-�.���O�d�""��A!@ޒE1`�s�$S=��p$�,��k�I�S��y��nF.7X� �K�?7�C�əB��OeKB���8h�B�I z�Y��8oҘ��H	�,�bC�I�#���;B���P#��*)C��uZ(�P��G^��Hc�9z�C�)� ����UB���v&�P��`J�"O�Xb�Ʀl�n]�غib�Y��'��'�>�x��$���&`t�D0q
�'T})��GEt8H��9n��Ă�'�� h����I����j���'3��X���1- ���Օ���J�'�vu�sGZp���rs�
�!Otl�
�'��@j��9/Ɔ�����:j���	�'�5��N۷����fnؾ`b�����?��eBl���MK�b��Fܧa���;/OR�O?�I�W�l(����?fI�	ha��3��B�	�n ��
�!�k�����ĭ.�B䉃%xԡ��@�^��9`Aßf����z���W.ȳ�p���j��7T!�$��4,�ف 鐿����T�\J!�$�t�
��6z�^��C@�r��	s�Il������s�ݒ�ė6[�>��p���yR+J&O00�5!F�t��C�y2F	�v#����A1F-�a���y� �$ e��j�R<��:�B��y�j����X4jW^��0���yd͉��XbB`g
�p����';ўb>A��(ϟ�J����+�0h�b�+�Ih��ܹ/ɫ	X����M	;����<O��=I���o��DJ�W�z��q�A`�<�r)�% ��T�L��e��Q�<��*�	�΀[�,ͳ-,�)s�
UJ�<A�d�䘰�"Y6g�̸�"H��y������R@W�G�HTqj(�y�b
~�����7?
���LL�0?Q.Ot$��A�3��X���_���"O��y%Z/t����e�+?�*�"O
]�w��B�ܬ��O�2;�ce"O�\��QjuJԸ����q3 ��w- �S��yR#
b�<HG
�>�PqB��0?�+O��ZV���z��#U��n��Ҵ"O�eK����e�4�Y���;�-��"O����/?��R��m��Lh����O8��+���FO	TE��Ȓ.X�m�!���3:O~���cև5�yJ!Ο}�!���r�)��5-��Q$Ö@���j���N��PAl4Pac�~Jy�c"O(Yڵo�K��8�ģ�,�IA�"O0Q��9)�&�B��'�QP�"O-Ñ�W�ř�'%��p6h�<�
����B0kI�U���N9?`�e��I|f��y+����J�b�|�ȓ;��TYV�*8�X7�^�P���Γ�?)���)��,�`��K�k� !�W�ϥ;xaz���ܮd��0���"`p@r���Vm!�d��K]4�2�fC%�Fh0��F8
!���OP!k�u��ĠUiM)�>��d�����	�N�9��?2��0����L`�C�I���]r�ጯ.gt�C���.t	B�;\(-J��D,I�dٔ��,EB�	)n�i�W�7X%��!M_���hO>[S��;�p�P�M����m%��R�����M_?o�m�#�B�\R�0�O�O��y���!�L-�l��4`B�"Oz% ��3J�D�҂�O�Y�̕��"O����S���f*�0 ��,Ч"O���C� <��%�b���3���"O� ���4XR�h��hE�<٠�;Oh�=E��Z�m@2��=J�;���PV�'��)��<� �p�#ğ	l�\ %E޳Ζ��$"O~���E=Q�NQ�`�����f"O��dL�ZF����/T�h�AB"O�B�N�,��+	�fwT%��"ON	����,���JGK,w
��"O C��B���X��Q
�rf$�S��y��� ��	�?AŦ�gh�&�0=�b�J �����<K,�y�'Z'v�'��^�'92(S�l�C�cD�Ȯ��A�&�y���catY������yx0�� �y����1H�q�� �0�4��^��y@չ{�Ҡ���ڳ٪�Gi��y"/P�.�����i{��T�����yrP�/�ȁt�
{`d$��'���y�m�)Z.P�A@xʦ���J ��O���DNnf�T�f��� ���\��!��Q������Q�T⾸x�
�*�!���ڜ{dG�5����H�<!�$J%	<jɸwD�0&����V"�J!�D�+b$�#fiյ)����!`}���l񴘈�m�$n�T"��Qu�vm�ȓ�UR�e��X$���f��%bQp1�ȓ{�����0,&`la�� "uEڭ�ȓJ��)��k�#�h��� �'��|��J���� IV)-$�h��X�xل�H��q����,nQ0��'i��Q�  ��Q}�9�d$�=������2�:H��Z�hu�1��� �90��z�쁅�_*�E(�JS4d2l��P��I\���lx)��ʠ.���o��ȓm��4�be��X������
'L݄ȓ;W�Q��2RR)�΄,ljՄ�$���U�ºp���;��!@ 8���=����a�)�ؐ[��]�%Ɣ]�ȓ-3��Q҂ˎ3j@�����.uZ�U��.�,lRB��9r����K'F0��<�N �Ѫ�):���(�
�4E��y[��e�V4�zE�f�`G�a��/��Q:Ӛ
���+��X�8p��*���J�2Zz�3f*z\NȄ�Ii�	���"�U�%�D!�"i� ! ����7
((c�	E�m$�ke>S�@��Iɟ��'����"�5?��xKV��
ʔ@��)��<�֮םiL�]xD�
�%�x�sTK\y�<��]�=����#�
�-(FTjN-D��Q篘4w�xs�T�|�a�?D�t�Fn'w-صh�6
��8��#D���'¶I�.t�n�;d�u5�"D� �W�B�m�QbңEh���7	"�Ov�pU��f)
([Ćt��e#u�j<��x�-j�P0B��� D�e3���i�����B�)M~}Q��кI�ȓ2(�Qx��R�	��}��g4Z��V�bЏ�1J�^Pc��`"��ȓBh���ĠG ���su�̣	.�	��oa�4�k�XXʨa�H������?!RiE�q��G�N���Ѭ^���'��y��ZRPl�K[����.�yb�@�&�2`
�%�W�yhX>�y"h�!��i:tAٵ~�\��H[�yb-@'��� ��/'���bT#W��y"�մ-��=�%�Hv}�L�c	W��yb���"��/��h�Ƞ����y��= ���ca �*R����W���y
� le{��ȅ;��@J�cF�u��<�7"Od}���H){z����R�^�;w"Ohj��B/GXV�r���s����a"OR	����U8` V =<k~�`"O�5(�(�ռ�H�p�xa2"OB�K���4�nFaL#7�pe"O6��]�j�@����{Ҹ���"O��h�ʔ�s$)[�d)�@"O$I�!k�Ffe;#���<�i�0"O̹��!R�.�%����ꎀ��"O@�#�¨m*��u��|1���0"O`pdY���4a� �q.���"O��2K�50�֩��_�L)L�`w"O��� ��R-���PE8��]x�"O�9�慜4��t{�Z�z r��C"O]裇Q2�>Ycb��F��Yy"O�QX=��A
F��÷"O��G@�e������ݰ��g"O| )�G�g/j�RK �G9Vy��"O�˗�	?�nIRF+ߘ}�$�"O�{&$�F��d�8��"O� �/ƸJ4~����&b�V��D"OքZE�4%d��'S޶M�R"OT�&�!��h!�4Y�r��C"Ov�;rb�FM,`q�A�$�r��"O�ݓ	:@��u��KX�&����"O� i��N��%�&$ôo��� �"O��y�g�9cn�xtB�\���"O5�T�7`բ���XR�`�"O@����-~��lbC?� "g"O��S��ۺ�8P���J���Q�"O�DR𧒁F�U�A�J��%s�"Ob�1�G���LA���(Z�a%"OP)_
�,�樞S�| ��+�y���U1�$�gX���Q�e�:�y��[�T�<
�C��\8S�/�ya�'�8t�{Z���Q�F�y�D(5���@�s�i��(�yf߾2�6�bdo�>p�n@A�	��y��- ��x�o�,l�r�hP���y�j��Re
9(q�%��DG
���X)��v��-rb����*w�P��T6�D+���n,��(��;Ct�Y�ȓi�4	���ڇR��3l�9 � p��Y�%j/C�G�rаa� c��<�ȓH:X�z"Dͅ�!��U:=Ҫ��ȓ:�0�T�g	���(=D���)��D�D ĩXqhq�0��	���ȓ(���Q"�w�4��#	��7D�ȓ%�Z��p��9�}k�+�f�(��ȓ$NT�S�BS)��c��ѵD��Ԅȓ,�.eН<�l��d��o�:��ȓF��y �'� 	[���>Y�X�ȓO;��b�d�N�J���:0�&`�ȓ^�.D �莺\L�M*�FV,ؤ�ȓ`�г� �0d>�T9�n��=�ȓyZ���Ȼva�91�@�v
Z��ȓ.�|����±{@+i"�4�ȓox��1��W�N��0�'m�}
�\�ȓ�L�hqD�Y�Q�G&��х�B�\���]�09�E/$�4AF�\V�<�b��?���P �-�iw��g�<�ca	�/y"8�ă&i� mrd K[�<��6=z�{�摍D\�� �V�<� ��wa�7ː9b ���e��"O�t*�D�a��x��&�+�x�°"O,����կ5O$,׈�	9sp�95"Op(I2�T�a&��t�����"OFȀkv��@#��_U"��fBX"�y��]���	QV 
k*�A��	�y�k�\&���3�
~ߊy�h��y��
:0Z!�6ϋ; �&%孟��y2/MA�� �/x��%�1,�yb"��Ii̩Q�p���y2��&�y�!7p<����9a몝����yBE�R�̽����U�R`93D9�yrLZ����7v֜�����!�y2�J�G�\��(Ukўdk�'@�y�h�=܌����c�0!��C��y2iF�w"�e���M ��R��
7�y� �<j,���T�Cu��F�[+�yH,��*0Δ�v
C#̑�y���qn�4m�&����虿�y�6ih`Btfg�B,��)Y�y�n�9�e�#Y==�� ���y2�(G�P1sF�,LNܙ����yre�I�>�8� IӮD��ܲ�y��R��*IHW�FQ�3p�@��y���)a�b�ұ���&l��.�8�yR�O��)C0� C����	;�y�IX".���s$K�0Q"��[��y#�#aZ���%C����	1ȅ��yb��/Y����2�x0S��	�y���?(�dr�U1f��R$���yr�؟)�VY�P'2zgd]:����y�+N�
��M�6@U�v NI�,C��yb��j�إ�'!ǩt��r�	!�y��]8ʌY���mF��j��y"兴<�%�nZ>v�X��R,�y�� S4,@F�.E�@v�X �yB(�j�.ir%I�f�9dL�yb�մ<����&��*
t"q�2(��y�E7�P}���&ad(s!��y"�ćZ*�L4��2��T�H��yB`�h���f�RE� c���y2Km�B�*�%_�My)zc�B��ybf�dXm3�k��|��ԇ���y"���vڶu*� ��E���F*��yR.Qm(��I:i2�ȶ���y�I�H��EP��P���%��y�H�&v|���L�z{��a�y�-ʉC�b���.��HlL�KTd��y)H,`��y���ԔV�ҩ���yh�QkPX�$�CK�n5��BY��y��)G�I�WN[�B�h�Z��0�yro�,Y�� ��f!�U�W"ك�y2
�� ���g�U�
����6�Ο�y�%Ж�Հ&i�,̨���-��y�"^5��ءh ��ذ��&Ү�y�N5�m2S,�3`��y��=�y���@p����=��{#�B��y�C�U�8�ᰀ�g@�[@ ��y�k�t3Rq�3�2R��hkӤ�y�C�Y�t��)[f��H��<�y��[72���9�l�2O�N<�aǍ��y.޴_�b��ׯ1|ߘqn�y"b^&��X�/@"u�a@
G�yr�Oe{
 ��l#��s7.�?�y
� ��@��;<��5���E�D�3E"O�%WA��yߪed�H}D�v"O�y�p�Qc� �4�Y-_h�g"O�US,܈
K4���	�~Ẩ�"O���M�)=C�a0A��ƙ1�"O�!i�I��*M l� K$���c�"O�m�"���!��� ���+���"O�u��!�6��:��S���� "O��j��6�T�nG�D��"O�f 
	t���F��Z��K�"O�+�X�XHa4�W����"Opܱ���(_FŪp��7d]j�"OHd8�D�2q���vk�$|jt͉%"O����I$z,�q�J���`�W"O5R�
�2�ꙑC̄x��i��"Oh�z'�%J00�T��9��d �"O��Z�-x
�e��ʭ�6]��"OZ`��:w���t��>�zl�c"Ovt�"(�[A�HB�±�ʌ8v"Ot��Bn �baF-�A�F�2"O]����&8C��I�K�+A��`�a"O�s�!� ж-�f�^�����@"O�U�ǩ�4�0 @�Ű tzPP�"O��	b��.f�d�X7��V�t"O��iFK���ȥ�N6%�
��b"O�w憡`ޠ�zDeǻ�Z,q�"O��ywg�M�Ȁ(��ގK���8�"O`h9�L<l|	�JԎb'�p"O9VG=�x\�,90~ZD�"O�Ȁ�׎���2֦s�,�@"O�y��1\Y��`�ze6@��"O`J
C*�H\H�X��"O�0��eF��,0�F5���K�*O0���f�]� Ⱥ�֘}`��p
�'��x���.���py�H��y���^)
�Ϭ*�>@���Ի�y�MѴW�jɚQ���	��5j^��y��X&0	�Hz��4\9h�hH'�y�ߪե��;/���!\.;f���ȓa+�!iA.m�b�z"G#���ȓaT�`�Q�CY���*�jў	��C�ɕq��p�!����@�m�XB�6L(���#�l���,'�C�ɨ��0rg��?��=`ҊØC�I�	
=X�S*e�]���.��C�ISP"�Q�ƍv����G��}��C�ɬk��amX�_�Y
�`�;VjC�ɇ
�x���R�2� QHX	bfC�	��(S�cM 3bL����/4�C�I.x���b"	ܟ[r@���#�;}�C�	�`�.A�d�A�/}(��R�ޯr-�B�I�f��Ac� �­�6�:j�B�ən��!��n�K�|��$�38H�B�	�Qmti�g�'���êߙ�ZB�� Q��ZP����ڨi$#�3i�\C�IDĐ�g��$|A���Ac�E�hB䉕�z�+���\���)
<�C�	�<�E�s %o�88��� *
C��$s!N�C"�G����#�	��C�	�Pl:g�@(G��q��ǔ�u݌C䉳 ���ց����J��ӟm�C䉡��	�BV�9��wF�U/�C�I�j1��rf����P�2e�K�dB�I-.u��E�n��i��H�%idB�)� ��;qm8*
����A�*7�p"O�] ���q#���ņ�̴Qs"O�H��
�Y�>}{�@5W���`"OLY�!�N~ �����]���	�"O��q�ҡ3�L�%�K�|��L`�"O��r%^)�ܔb5�9�B��"O�щf��#��3�a"7��@�q"ORQI72R�ֹIǀۑ|�z���"O�eJg�T)	� Y8���(�����"O��rCC�!���a$�r��`3"O$�B#U�*��`��"ǓZ��u"O X��\�>Tz�,�����"O�����$]������y��-��"OPJ�H�� P@K]�6��"O�Y���	u��h*��)8�p��B"O�8`�,A�q�UiQ"N|dx��"Ob̢�F�v	 ��'�>��A�"O�䒱���ѡf��`�$��g"O2��U�X6�(D+G���5�`"O�%{p�?$ޜ�&*�]n\�b�"O�9����;�y:%��>@^��)�"O����\P�)6h�<L@�0"O�Ii7dxG�ECҭI'>�� !�D#�S�S(ut@h3��&;��2-ݱI[�B䉸Z�����U�R-V�xn,�<�˓L/>���FurX�$$����P��y�`$Y�-�'H�rI�2�\�c�b$��9J�)g��4��53�U$h�4 ��
�к3���q6]�E�P��ȓK<z�!WH�mE��H6�Y�e<��<	3�4�Şs��h�քK�Bmr�87mٕR��ȓ&s��H��0z�a1lX�'ld�GyB�'g��BKK�y�D�������9�'��dY�Z<�����`��J�'\�H�aӨ<!D��.Y�T�I�'J�}�`l�kQ�� -�Y��4!�'Q�����E��ѐ�)ŝOPr��
�'z|�1Mڗ}-�T�v��M�6��	�'��]�Sj��1�$k֎Z�BҴ�h	�'Y����"cJ
�EH�8���'��a�ǏF�s���qb�ݷ;#� ���0<Otb���TMrJ�|m�yW"Of� �-�Y�Q�B���M>�@��"OF�[Q�Hl�s����#&�08�"Or(j	�K=(4��ܩ*��S*OfH*�D�4c��E�[Ԁ��'�����ɂ�QF݊��[TĬ B�'��(ɰ�T�N�:��`�ɀagX|��'+�����:T�Y8�m��_xn� �'XP Q��%}�d|��6Y����'�~<{u!�,0�[��֡H`
A��'Ȃ���쉿W��LҖ$�!*wt��'\���.^���%D��rh��'�
���BF�OAH�Y�Q�;T�b�'
��g3V��p�TGM����'��x��RY�dT�c��J��1�
�'������f����R��5`���	�' ��"�	w�Ĉ�IQ�& &�x	�'�"-ka�W��Рs!*g�x��'��T
�������d`$��r�'�����a�-�r���ӌ�&�9�'���kDFΏ�� U�\̾q)�'����� D�5�ԁ�!*4]d��
�' |<���X�PyCa��0'����
��� ���O�=b660c偞�1b�:@"O� ���/���qnЭ5(p���"O<E�A˧� d ��T=Wh]��"O:��#o��$���O&��'�xU)��ݻX�d��#�A)�'?�0��Ę�"�mf'Ƃp �X�'^���b_(c����ׇzF�X��'�P`���6H5�t2�����)�'���;�[8(��Q'ʙ)}�~q��'�v�[�#�g$LdxF$�8C�&���'	 �ɰL@�L�Z���D��?���p�'z�qq݈JP�ő���7y���'���K�L��<�낎��/��i�'3�yKѭ�'7�-����!� 	Q�'��)u�G�KM� ywI�;b6(2�'�	�$͈�D�m���-a�����'9�)�ťF�+w�]��7WN>͘�'��X�P)^!~غu���U�"L��'"�5s3瑤�h��ǎ�GL�I�'`����bU�����
Of,(�'���	qI��^>�UxHޜ@�vZ�'�>��-)z��M"��թ?5
%#�'vH ����!H`������1>�j�0
�'���j��3oH)��%޼5t4M��'lMz!lۢ������ۼYpL��'�Ak��<��iw�.(C��'Pİ�a�	dc ̡�#շ$W2�P�'m�F��/���`�� �x"�' �$�'A�#�b�a�g�B�b�
�'�nQ��D�C�L�1 .��4V;
�'�n��wE̍.�����U%cB�	�'� *��B<�6L�e�K�x)*	�'�̅�vnL<��`�>2�4Z�'����i�xi�0ԍL
&]���'>}����v�sGG;���0�'=�l��e�,�,�+ ��1}=2�I�'x�h"$���k8~�Ag	Я('�h�
�'�H�br��3J�xx��S(�e��'Y`����;��Z������'�TU�FW)�.��
J�P��5�'�~��@Ɍ:�>I G &^����'�2!W���A�B����J9I��e��'�BI�%oW~��ԍ+l��1{�'Ȏ#���>���	�"՞_���j�'VZ� ����J4����Q3b���'"D���I�'x2aP�.ڍLѰ�h	�'����͔+J�y�ӁZ��Ly�'��(HIގ�l R��Wv� ��'�]����R7���O;I���H�'ۈ�-�%f�*xɖ$o��i��"O��qC�4J4��"���d��jE"O�kg�´4[��r0��ASV�1"O��X��ǿ}�Xe"@
D����"Oޭ��蘛&�8�b�`��%4�c�"O>�ǯJ5?�PW�D'x. �X�"O�@`w�=O
��NO,Kd8S�"O�$��P�@WZU1Z=>���
�' ��W��Vj}���Żf�hM#�'�����Z?�� �ş�S����'o�����I���y�iߋO����
�'~�  �[ ����#)֌5�Ř�'���3EdZ�����q��$�g"O���1Ȓ4JD )ʑ�t�� "O*�0��7ZA��:��Г[ ���7"O� ��Va�.|��Љ0 �4��"O�A�M�g��J��ټqE��"O��s�L ������Ѷ,e� "O�AkG(�<�U(���"�"Oq�w)�|����e��<��|!7"O`!�PB	4{9�����O�q<!	"Of�	��]$%C<%k�cI:'n�iV"O�,e�X� ��ܓ�aAO^�D�"OD�@�K2�r�P����,#��P"O��t�?o�H�x��*^�б"O�A�(�1�|Q��1T��a&"O̝2�O��N�.�1����Б"O�Y�+��	���P��
Q�D"O���H
�SN��a�!�f��4b�"O"m�b�\?6� 9C+_�L���"O0��bÿLg9���_�
�:|�d"O^Y@�H�����M�Jeh�!"OT<i�۾i�LH7D�,OE�A�"OM%� k�ȁ�b�w�@h�"O,��`�]��d�O�< �,̱�"O25�1]�r�#AM� W�@t"OX�xP�4ehcK=<: ��"O��͑��HP�cU+}6Ai"O,1�E!�K#��R���WR��;"O�\K��1^�q��~;6��"O.�BU@8ھ��Q� L@�0"OxX	1�Z�K݄�1D.>}�.�3"O&< vhK>Q��M��� ��"O�̀@�˜I���z���R^*Ԙ%"ON�QpjQ�I��`C�ɶv{�5�"O�`�r@��O�`�V��5`o�4 ""O���efc|!y����G����,D�PGoҏ����s�O� �p��?D�p��"�X��'L|�I#��;D�8��7'��k�
ˏh��Ix��;D��[��G>(@�����u�肱	,D��S%('�5su�@aR�/D��r���H�2]�&!A�A92Y�1�(D�t���Q-.�訚��!��H��!D���Ҩ��&�`�k\�$��(b�?D����KC�U!�T)@D��p*��S�,3D��0�@W�8���N�x�×,2D�p��%I�7E�Y�O��|4� ;D��q�.	=���kc�(�(Q��=��0|�t=ݦ��QǗe8-��ęm�<��Y�e��Z��� ^ޢ-!� �`؞��=�##�Srm�$lY�w�`�SaP`�<�P�L']DF*�͔�Δ���Y쓏hO�O�q�	�F��y� �<_�0#
�'��5ˢ��4�pq��&�RXt��	�'��x���:	����H�4�		�'9n�@C�ׇyPXt�`�+���s	�'|�0��p��x�G��\|0�'C���I�R��hϥ�JQb�'�>hۄeO��
Z�݅�� �}2��^��ħ�B�H��Y�f}K h4]a�8D��S@D�����p��(9\�)#;��0<A�h�aŉ�`ڄ B�A�.�v�'t?�Q��OT�da9���;hr��q�:D��z�J�5v�{�'ۉl�bѺ5�8��}����'#6l�@��$	}s񭓪Wf���'�񰂩C�.6�dG(J>��Y�'�z\�����x�T�B�v�"9ٌ��)�D���XQB� U�8)�h����y
� ~�go�I1ta�Q��w��9x��)��=G�����ĳ ~��8�S�W��B�	�0g2T
�nW*5�&��*�6qlB�Ɍ/�>�bq��`�=LQ��>B�	0`���@����bn�\��
	o�<B�I:�Dh9��إ6�Y�/�0B�B�	�$>D�@#p5�`��hS-:��B�I$4�\����^�*�H��"
@��Dn���BE�b���A烀u�غ�'&D�h�r�)[kTzR�E
`���4#D��Js#�,h��it�OsQ0e�'�,D������&Y���k`��2�Z�;@F,}��)��>G�11�� �|ۂ�0�<=�ُ���O�-�e��,3�pZ#�Թ����$�3lO�${筛1 Х��ۺz��p�O~��D͓>�
�����/��a��BD7J!�E�`oL�åM$v�^0�Bh�Z!�$��j�*<�i(�h���̭@^!�$V�kQb�P'c�=z$⠡C+B!��C�U&҈p��;\��̳�`]�H�!�DW=G�~1#���maܨee�C�ɚ�4��&���j�Y��^C�	'MJl�sqY�AI��!�iH�Z�R�Z�'�h�,L��0���2�,���߸�y�W3<��	��[�~�}H��P��y҉�<B�L	0c�#AjUQ���<�y��-�Ɓ�H�:~J|p7 ;�yB�}�譐+B�,��MKԡ���y����P��2��p���࣏�+��x�����H��ց;��;�2!!�X�l���w��7(J�H��	�!򄈵,g^�J�"ڕZ!�4ÅV�\�!�$��^�)�aԔu{t�x�CA��2�m�e'�$��(��<�C����'T�����"OD�A�A�X>���`��N���r�"O9�7�Ą34�ǏZ�d�N8�W�UH<��`��=�����X @�H'����<� )�I�k�x�C�O��}7�a+��4G��B��65��1q�R5[�I�С�5�b��=���D`]	�j��'N�f��8�D�W9�y��]����#Ň:�ʍ�� L��'�ўb>e#�%M�-Jthр�(�$A���I,*X��M�7`�v��Lƈ�t�'���Dy�Oω'�L2ӢY�͡�.�B��x�'�2hf ̦=KLt�f�#~��Ӎ�'��t�QG8T�EQV�R5Fמ�@���%���:�-@�J�07�NL�T1��D��0=ɖ"W6-lvi��E�l�@=;co�����O�ӧ�g�I� L�JE�rԤ�Q&��_`�$.��AA�G0iJ�J��K� w���M3D�X��Jט{���jc�
-n�&����6D����0o���c�	�5 ) �
e8D�D[�D�"NL�FA�3"x1�I"D�yS�����&��+�(v3����M/����U�T(�ae��%1K����Ej�z�A0��A��^:�=��
8�-�Q�W;Jd��q�K�g��p�ȓ �&��%ԄIl��!0�ޅT.⌅�D�'�N�{�䆪���Qa��L$�<0B�>$�,q���*
<y���)G�����+D��z@��1�e���V�q��0�q)���VЊ���a^�i���I<q�"Or@�c�fC�$����7Wu*�"O0�@ɻ��)�� ~��]�W"O� Dm�E�;%xLK��S)��d"O�U��	�	���s2˔M��X"O��A��PDlQ �X
v	$���"On�9A��4n\�x� k�$�a"O��I���2C�>`�S�Ъ"�x�&�'H2Q�3����dC�#��IA�,״<�|�ȓ7���b� �.4H\@t�������IW?�C*�<_�8h�������˟C�<	!`Е	Z��PkГw^z�!Ak�h�'�Q?=�S�܁xdH��&�G2��d`U�-D�D� lZ"+���2j؟H}�H���)D����A�@���`Sl� `�����h<ꓦ��&�PAW�:@�H4뒊_HR�cR�8D����	&RGxБD�L)Hr���ci5D���@ �3��0�$�W�9&�E�Џ�>i�
)��cGhQ$(�a*�N� \\^����5��cˠKƒ!b���Q�%��;�����	2?�� 
��ґb#f1�ȓF=�Q� �� c�2�0�x��Gx��x���3\����}ZT`���K� B��!^->�x増�J�L�����I����I�D�'����s��sdY)Y�y���<5F ��ƃ�O��0ꓠ�'j�p�+�r�ذ�ʅ�9g@�z��-O UB�	o�C�I�wp����"O��s�^vTl��]v�L:�E6?A�9��h!VJC95��L+�b��w>8u��~3
-���L%=\"���
&Z��<i�H�U����.p@��T�F�`���>QÓ�y�BI,R��Њp���[֮M��艡��x�T� ��h�f�	�HY#BǟZ����,�|t� �$.�#
��PG�Z��ɅȓuF���va�1Dnz 
&bԅ��=�ȓMBx��:�.m��ɐ�0����V&��Cb��u8�!�o��A�]�ȓK�!{����Ҧ<���
j������?�6f�)O�TMX�dμI��HP���k�<�b��7뀔���Ԟ#�*d%k�<�g�ɮ`�;��	 0�&��2��`�<1rO�,<=�Q�r(�|���c��[~��'[p��d��<z
,�g(Ȥ �e�
�C<�	�U�eۚ"���m���D�P
�'�$���ퟱV��A:��4E��-��'.�)��H�smC@�[CU���'���J�L�6c�����2O����'�p���[ Ej�$��J��b�'1x�0Ǚ+��u�DEM|�I"�'����(�*4b��cbߋK|>�Q�'�@�ZxƙHB(=>	��'�L�
f
"EJ}�LV�DUs�'Pă��O�=e$"%�<Q\���
�'j�E)Ȁ|&�tH��}+���'����H�j���OK���ܛ�'����)X?tq�a���I�43�D�
�'n
��$qx�,�$��'.�q��'��P0�BʬS�Y��X�M(&y��'ApHi�$B�?Ǿ,�q�4[4���'bUz fA77����i�h@��'`h�P 	�LP���`ɖ\J>�q�''Ьsǜ�.�|����hD����'���s4�	$B��I।\�H��U�'��9�����]!�y�(&A��B�'��m�U���e�&��IZ=�f���'���RD�<n�mj�pL$R�'.�m���B#8����S'�<l�.A���� ���d˗�lp��r#�Â4рiy�"OPP�g̸A�4#���r�,�S�"O�LzF@ʫ��U@�Ɏ=˂���"O��Å=rh������R(0c"Od黢*�;1����5���]�k�"O�b��G�^�~Yb3'� L����"OB�kRX=�t(�z�b��#"O�@��O��`��D�'��� x
L�U"O����M�?"��!&]`ֈ�0�"O
H�T�W�A�kS�0�aD"O�U!�L�7#d�����$.�B�C"Oh@��)ֈo�Z9���"2��թ�"Ov`�j�Lv�T����>A2��"O�t����?\���[$��2�"Ob��嘮>f�C5�
�0�["O��:�҃C�%c�ƛ	F�Dx���-d�0@􁞱!g����H(��S�P�/ ���Űe�!�d�, �V�A�
�QmRh�6� �!��ւL@4�,ƈ3�x=!�dE3f�c�M|��P�@�!�؍�	�'HL�)���:��`�E�Ҝ#z	��'�P��ԯ� ?xq���7!:P��'�"�H���5��m��᛾{g�`��'�$(�c�!�yǌ	�u��8x�'��cU#�?v4 �Q�D�f^\�	�'�zt�@Ō# �Z,��dQl};	�'̥1���$�@��%���~#zi��'Y^1�� V<v?��SVk
eE>MC�'@*�{׮�8d�Tu�gآY�dܳ
�'
 �`$��:�4x���ZBj}��'���cU��F�ej��\=H�&H�
�'���!�*��i��B�&Tu.�	�'��y���K��)�U$�V�*iY�'�.��I	'.j�GX5E��i�'�$e�@�#<����g��9:��']M��aǈ2���3�-?��8��'�M)R�׎h'��q!T?/�z�K�'¾mY2&W	e�"�b�MӮ'̼��'��m��ߊok③��E^L:�'��C�8:]X��X6���y�%�+VM�qC��*L�x�(�<�y"��"~����v�A9Qa�g�ϋ�ybiJ�G�8y�ϐ=V�������yB�3��0T͏1���XV��y"�Մ8�Ν��DJ�6|!��O��y��M�'
�K��ִnİ0e�I1�y�JY�l ����K�\e���3���y�E�?f�H��V רM]Dh藰�y�˼�Q���@��@�B����y�o�+YR��Ct��(ԐYB���y�#�P.�`-[�r��zr
���y���X�:-�P'Ŕ(5�T{�陪�yr�[�
2pT+�BƟ*Bj�Ě�y�hF�
I|@�!��u����VѠ�y�=V��<bL��c%t0��j��y��F�x(�@�O�����/�yk��j�tK�fU-Z���b�,�y�+�a���&A�,Q%�y�Dq�	1AcC�a
y8Ч�(�y��?`y�5-�=��S��	�y"*
-*���/�>c�LR;�y�`�%n�8q��-�&/0䉢d�:�y�� #�-;F�[� 	&��b�ʽ�y�Ұn�BP�}PqB!�ݛ�y
� 2D��!ӏ#4��{�o�1�ޥ��"O �3BH�b�6�
C'���Ձ"O�� ���Tp��C�	D5�|��"O"��!�Lm���q(�%cZ��$"OL/u~��uű?&�rT��yb�10��zE�"�p���O%�y2`M�"�ݙ�F �Z����\��y"d��
�a(F�����Q�,W�y�-A�H.���sÅ�i��'Dӊ�yR'_z�Q0��x����hɵ�y�N@�'	�������֋��y�F���.
{��@��þ�y"i� Q8؍c���5])��������x"`�,�����8/,�C���<�B�I�g�xhܛi^�+�A��8İB��*>R`��o�a�.��䨄�9}HB�	� >��s$
����ĂQ�<B�I��|� F�,/��"@�Q�a�B�T���rVE��f���@�h2�.c��H�HP���xr�&0=H��W��I�2�sSN�+��?q���Lc4�HaM����2H��[Q��1�%ÎԶ���P"j��h1(ڌW#_184�B���@�c�Q��#ip�kA�M7P� �Y����!�TI��4Fe(�ȱo�����Q&x���	�C|����M�Y�u�g�@�O�(z�-��T����������� �ǓY� ���h�E��t��ɱk�x��UjBڟH��r�� ��LGx��y.V�
m�Kg*�,`����Q��PݠF��u�a{�#ԪѤ�a7��3j�\�Q�3��kEs���x�&�4����(8,��ǦG�7[�����N㌽���zlx��T�L��0�$�3��x�r��\葞�Z
�'JZ�A�r��lt6P!P7��l��šo��8Q�B�_f����lhZҦ�ϒG/�(��� �s�0���& m���|�&�P�o@z9�6mȝX��v�Z/Y���VdWmڒ��E�`X�X��]�_K�Q#�&8����^��"\�FW4hٱK�(ݤ8��LՐ^*�=Kt������+���*�OB�uF> {��zW�:@�BP� �[c"��gZ�p�n�3To��)Ӣ�:ǩG8G�V\�!`"_h`iXj�,j�SW�碈b�V�� �`�;v�T">��`�R����jU�c�T[�M������ě�c��p��3����4��PӶlY���fb��{:���	6k����l(,�bl�A��{��-KWa�."��Gy��I�.�rD���V�|��'�ȯ#��N�1��|bS"P>KJ3d
�-�8Y��$1*٣A$U3F�T��j�Z��h:��?��O`^�A7G�/(�;���f1丗`��tpI�"�D-��@xn�I'Q�-/�[��T0d3���L��%ġ^��!��P����P'@iPZ4�%�d��I��N�p�ӯk}�O}2�̍Y��C5)������'Q�q�ژ�ݴv�$��C�3:��әX���iN�����g�%p�F8kB���*(\��M�sބ�Ǆ�'P�X�"��(YԀ">�!��s�� Fd˭�x���Ǆ�+��1O����*`�VzxJ�r�X�a��X�g�L� �f��d�Q8��X�<��"���%ZkX}K�0� �0���DFHˊ���7��9�Eh a��K�"'�E	c�Z����[�`MX�Z@�eܝ"�\Ը�jH�u�P�u�X���)E	���K�П�DN,h���^aZbD]iWT�R#�?bl6�C�MO��s�� K�EƷr{��hR#C)JG��sr�

��4��P��_@��dA�=��i��B����䟀!N��c�OX�(P$��4�Q��^�3�ݹ%�����BC2f����4{ƙCb�|+>��B�j����M�v�З���O� �`l���[�Y$ꨳ&�!�O蠫a�)N��| S 9G�Q ��6m��r�K��0 ��s��ɴ�Qc�
�e��ID{��L�)��ɴ0n���+�m^�ep��ʜK�h#>��͢R|"���OU�3	�lk� ���̤^��`a�ҭ?~�6-��H8��J��С��Y6�&�?�	F��LrtJ�"o�r1�FfAv}�%#R�u���	����T�Z*-*5Z>%�v��*��UP0��X�f�#��
EIU�����rc1@�l�4��*�)bA
���~r�$3ےE��hQ�R!^��!~��xJcMy��Ӻ�ƊM$�m��@w����M^�<��b�b���s�l�j�����_}�ݺg5�D��|�O2�X�V�py ��	|��r��׍,��͚W C��y
łS�L��&	�5�x0#І����5�p$�)�0<a���(nH؃�CD���@���O<i��R*K�쩔��-�� �F$Z���(��*V�͌d�
����Vz S)5D�L��`��]�A(��t�
\�CE/D���f#U�%���8U��؁Q�3D���aI�[x�x�&ě7b���!1D�� 
��W�e��B �p(V�f�'��T "���B��z�H9�p���L�>3~�����p>�q�D�!����e�fC�Y��.j%96�B��5|���	��/�0 c��~�T"<��h�*��7I����Olj�����P��W�vT޹r�'��ȇP=Z�����kA~y�0i?�h�Qu�Di��)��<�
Ԇ�!Ƅ�4!�Zu	L}�<�U�^%��s�X"	V��R��<��M>!��R0�E-��<q3�R�H�"��d��p��MS��;�L�+j>���&	�#z��%h�a^�]��y���VR�r0�Ɠ+�6��c�	�]�(����. Z�Dx"���[�]�U��>��𘪕ԝF�܅Z�@�.����"OF%jK��s��x�̃�&����#T�� `kW�я�8�S��y\�.�0	ۣbN-T(���-E��y��P�"�6� �D-���S�㓭�y�*�SJ��貫=4=�y�d^	2�L����)/��	2���p>�§�� n~1�w���/Zm0�"�5!��Qo	6\���ePB-qO?�	����A�Ě<Hn`��(B�X�8#=��IK�X�(@��)�n���1A3"8����7B�b����!�'����5U��L�R�ϩNrl�	�i]�����a5���>pl.Tؑ��+ZZ9+�ַ#!���Gu���p�@�p,�����&�O(�1Ci�2��Y����V{����Z+,h�k��!�D�������1zh�׋#�j��W�O	���'D�#}�'�@��DʌUK|�	�&
�L�F1q�'�����o̻{��(X�:�*`	�4V����C� f����*=�Jغ�#L�g N��`�[j�a{Ҭ ��H2��͟���N('���*�� �&�b!.D��c�&)0�)uE�D#�z�0�I��NS���z�>Q!&�'u�;㠜>n�Mۆ�"D���q	�>P�]1��ܗ6���"ܾ��m�SE�U�D�x�����&X� �ᢟ�pҸ�tԸ6�!��$Ll:m��aҮ=�sFF����),��3�'��]CdL2���˦NV��R)A�u�N|X�j��7�ҷA��@�LW�;#�Ad(9D��9eoV�G�6�B�!�[���!�Ͷ>�����*דX��X`Fǆ;�����'~졆�I;��u�׊k+̴9ݔ`h����	,���Zb"O�1�Q��W'&���.X�Dy�{Vቁu�fE[`C�JH�:��+vN^��&@�)$L,�9W͌B�<9�L�=q!@�� �*I�� )q��2�X�C�BE����,O?牞Q�U�����>@�FK�\��B䉊.�>2 )��e��!a�P���	��|:�F"����9N��*1F:m���e^1���d��,�"��N�%MX�`�	�r0�2�%	�(��/4���`�7��x $�AI*d4L<M����A4h*F=���!��#nz�#�M�NE�Q 
��y�i��`��I '�8U��y��T��ȡ�N�zBu�sU�"~Γ�js�H�j�k>`r��`�"O����%@�ơ��l�9E�T
f?OQ*���;͘e�s$.<O01Z�L.+����:7�l��7�'��l�E���N�R<PZ�y9����C"b�.�#qʅy�<�ԉ���@�kjU;&>��rp��z�'��y.-&�
��
�v���*W
]��[�iE:+t!��=Mbб�E�;V���WJ�	�!�DS��:]��MO�| ��Ch��}�!�	t��d '��y���b�_;#�!��Ȭ`�صq�$դ@m�@捛��!��ʒR���	�BI� 9�&Y�`�!�$���V:@Μ�9(�--��9�U"O��zfGA6����bˍ2 8YSg"Op�P���v"� ����[b���"O��z��g��ܛ1/�">�+�"O���r�Ϳ
i�-H�Z)Y6�ȶ"O� j��7ʔ;t�q֡�:�J��q"O�}����yqj $@G`��e�2"O�mI5GL>�}&oP�K^r�p"OZ�#LH.*�P�s�خq��1�"O�Գ������g��Y`���"OPݹ`��*��@«�4X�e"O�tH3�N%+�,@FH[�m����"O�]���%x��H�����D��"O,m�	#��)z�ə0t�b�*�"O�9ãk֍=A�Q2�I΃��x#"Ob��䗢
�Qs�H"[ȱ3"O�ᒡW�&	PZ4"C��H��"O>��	 M���U��2t��)�"O�`	�#�n�F��W�̵|+`�i�"O��Ӓj�JҨ��	�5�]�F"O^�e�j��-�d��`�*"O�uy�g���Y�JUS�`��"O���"��!}%��q���6X�X��"O�}� �OȒ�S̀�v���*#"O�mAv&H7�U9�L!&�f� "O,�{uLW	CR`��d�@�M|>Ց�"OX-�H$$�ؑ2jX�~X���"O��(0-�T6�3�Ԇn6�q�"O�*%ŕ-("�Y��?X��l�"OL�¢C�:�i�i+d�� s"O�s�	T��Z�Q�T]��Ɂ"O� *4�MȂ�p2-�+]�M�"O��[�kO	ib��U͒Hh��"O@�H�L��HF���́�&�@`Z�"O�IfCŇ#yn�QaL�
)D��T"OꑺB#�>"�܉*!Pu�h��"O,`�� AC9P�gh+^f��ه"O�xx"�]$_U�x�$L؇4Bz�"O��ǉȯ\�:R�+ɫ)�5�t"O�����F ORf�c�JK�8��""O��c����h�.X;6�S�"O�d#����h!D�+z&q�"OzdsT��>x�F����8W"O  S`@��/1��B�Ɓ�t�l�0"O��!��1.Ed
�kA(]j��"O��� )�DD+d�>[��)�"O�F$��&_�u�s�8��91"O8�+Ӈ��Zkz�y�cX�\L4���"OJ-[�OP�P�!���8B��"O(� �S-�YS���&h�	�t"O!`��_�蠍[�n�b���"Or��q鈋LlTȪÌN�}|�"O2��'W�
����>��Ad"OXXY��+U:�چ�]�^�,���"O�a�wH�1Q�P��-�"-��Ԃ�"OΨKAB��L}�x��-��!��æ"O}b�OA<ym��K�^�z!R(�2"Ot�2֎H%b=��b�=*5��p"O��a�jY6�
�jG�V!DR	�!"O�%[p-�'���$�Ws7*	!q"OJ����RR0���[�$X�c "Oڴ*���~1\%Ѡ��rO�0
�"Ob	�",)� aZ�Y7 �/�yb`�%z �mɁ��=zҍX!�y�H���0p�Q�4�����^��y�D�9L��G`������n�4�y��R��`����	��[׆���y���%/��d5�G��� ���7�y�$֜%R�J���5*���@E�g�B�)� l�Ĝ�1s���ggA�1�@ɳ�"O ((�Oo�MCtK�k��T��"O�-"PH�P�H �jZ��p�"*O�����V�B�:��a`��&�Y�'G�I3��G9B�*(��ΐ�/Ǻ��
�'�q�"��{�C���4I�	�'Ԧ<2WO� e��M╥ѻe\C
�'�r�S�V/g���F���T`�'	���͞o��xBg�Pb�'B@CF�	�)Y"��6G�M��:�'� ��49���{&����<��'�A �jB�?�hT���~��|c�'P�|p�J+w�\t��"E�u>P��'IP��L�"e� da<c��4��'�i3����kۮ!�vGY�X���'l�@� J!{��8�P!��T
		�'L>%a0̚RW��@Щ�:|���I	�'
"�H�*��/A�� סV�$F�ћ�'�R�@c�O-ظ��g ^��DUx�'��$`�(�DҤMC /Yja:�'���C�̫0@z��hX41�'](y��G���&��/��eY�'��Lka�.hl�[VK�e����'��C��Me���eg����4h�'�rM����%Sv8���0Q���'�칉�h^3��zŉ�x^�X1�'\�A�k�*�Ȭ��(M!s��l��'���Z��@���@�#�ęu.M��'��(�@�P5F�B�D
J�`�y��
 N̄��/m��(���V�p�(�0lB�F(��P/o��<��/�9+c���}�*�Ϗ(��C���Y�Fd� �YK$�Z��U�qQ\�=y��@�)���ۇB��@�	W����0�\���}� ��6�Р4(�H+`
O��a�P )BEȮm�ƙB�o�?�T}(u�A R�Ċfk(��c�U�R�|"�	|֙� !T�T>V�� ����0<�n�
�|�ڑ�<}b��h��E*D�Դ�%c�B�����Y0�N8��
L�_>�5	����!�"

3d�h�r����xJB鐷���.͡D� ���~��D�#jWPivL4,���QoB�")�t��ʒH<i�R��`�2��B(|ON ��^dA����[�D��ɻ
pKV�%����˃�&� �a����ݚ,(�q��Y�2��%�\15y�B�I./Ը8�D*b܌1c��S�z\�Bƅt�R�Z'l��ګ_8�|A�M)X��ĉE�#=��2��R����I�4"?���*�X,�%T��S>]1�-�
�&߆  s&�= ��գܡ��;2�	7`��sP��~�`=�	"��xà����U�g�]�o��I������?�lCw����)��us�DV�c�r��W���"��dhd"Y
	����k�;{M��x��O���=閬�1q�B���Y�-}��R��=l�8�d�����È�E�=� �\:G&�[�*�;8�Py$���*i�V��,`��:�h��^	����'K���	Ҵn�B�0Ŗ7ES��I +>q�N��ԎPfm{dE���3W�:b�@�!�?!�ɹk����-��-c0��^~4����4�F|�պ` ��r�k���d�/��1sCE���l��N�U,q�'��/4P�"!�F: �	I�Ჟ����?#<��N�Q_�M�s�# ���bZ�<	�[>��� R��<��ԕj�����(�i�\�Pm����i�J� �!��W+����ΰ0Dre�8N�I�%r��h��R�|vȕ�uW�˲�I���Լ!)l�r��9K#���.ǙX;a~�c̭��%	��[;t�Z9lʎ�� �3�˴}���'9(�����*�@�E��Z�.���{D�RR�,a�"'����O�\��U3p��Pb)OPq��_�L�!ҕK��hh��J��.���`[#��?�5
�HS���gW"a��PfFU?����=��O�찴E�Ovz7��T�JrK`b��&w$���`耡�y�l_tP��4@ČT��'�)���'$j�Z �&�4�d�b@H���C�Je�3Ʉ�e�2��(%q!��Ţ��(�FM0;��q���<��'��a�Rf�=�ax"Ț/Y.�@97DDX�ƹp��'�x2�/X��D�%��ظ���ՙ5 l12#d(<� B�àA�-o��c�	�,\I�	6"O��K$-V3�,�H�n��N4�A"O>��1�A[T�e��- �."��k�"O:���#��K�@I�C3O-�(��"O�ؐ�O\6����� {�.��\��a��Dm ݇��0F~�5(�j��$�IU:?~��D�$W�*��e�d,�5]�!+��Vzp1��'6����8lU8��m�;~�B�����(r�p7m�sڨ�?-H�턴:g��	e�6�����j&D�P���\��$�A��̬� ,�w�zՐ�(̀2������A���u	�=�4(�V�(-!���7NLS�K�TH��jX
,��D�v��d��"����ָ�����V8`�,�5FU1za|�ǉ�4���k�+D�z�
���n	�e�c�!?&���O���^�|*��XCo�oc>0P�I�<S����^l�Rm��u"��$^4NZ�=p�l�Z�<��I(jH�8p���XT�A\��8��&D�晙-O?�ɵZ e�/k8�p%�0��C�>_h�=�֩��HP�A�%��@Zlז(,�}��'���d��bf�ȥ�֠tDl0��Z�����O2z�$Q�s���d�s4�ЧP�̑2��J�?��0[v��s��:�ĎS��IsѣR�����6�o�x�aB	)�(�NiP���8<��}y�Z����RP�'���Sؖfwa|�KK�Qr�:6,�5+`�BDF���=i�ƅQ����a��O����{�������a�N6"O4U�j A+@�)�d�3�J%Z��d�ԍ�.�h�<T�6�ˇ`f09"rɓ0�(��$"Oa�;rz���9�pe��-�$X����#`'}r;�g}B  .�Q���,�.p3ݴ�y2�V���(���0�"���ݿ�M;���USf?|O��ҥ��1Y�ti`�/�nA��'n� C!e�&O�Q�I,�<ؑ��&U��r���[O�C�I�'i�9�����<Ӓ��3F�!&�c���HwÎ�a���LZ�(��\{d�a�3h�C䉒kNn�
�Eߩkn���Nw�X=����S\�OL�F��Or���.V�U��9*âƑsPw"O�hIU��� lq塑�J�d�	��'4|����Va|���b�8h9�Î�xq��)�LZ�0>���gи�ɐ{�A@d S��"|B�kڨv\:C�I5uX�i2�jȈsZ��1�D�D��WAB��B��p=	�o��_$�%{�5U�
�H���S8� ;���� J���C*h�^ ��M*6�	� !W"!��\�D�m EA͹f��1���"Cn��H4M8��)�P��Z�'F�9K��*^έ��cW4_Ixy�ȓL���\�C|���RO?!�4ل �Nt޽jD�߈���s�� ���(3,4"�` ��½�q*O�pf%ŊbDhT埱D�d�q4OV�愀�@Y�1s��(<Ox�+���%C���Ƣ^B�L]�F�'�*�
���ډhf#*y�����d��
�4
�̎�-4��t��!�^�b�!��oƸܒ��Y�N�+6�B	 ���׍ԓt�@a����ؒ��B�<���^�-�2(��oi)nX��=m��E�"j ~���.O?�
'tI�fLN: ��,Ѣ�єR�B��f �b"�+�V0)��4Pc>O�qqgQ���2h-<O�UY��F!l�Q���E���h���'�R,��%;jQ��Kb�����3ˆ:o���Ip�^�<��cG;CDL�E��z,ye��Q�'�����!#Q>�:�J��f@� ����	����7	;D��8���"p2��@�*.��&8D�Tʒƛ-��|����v��
d`:D����"@�բ���<SDxD�s 6D���P�Q�b�����L`A� +D�����LsPi0�hޫ/�Ȉ�*2D�D�gi�N힡bd��F���P2�0D�� ꠈ���x��ką~d��"O��@@�:X��l����	(88I�"O���@�l���ѯ��5"O��B,��'E<�����/����V"O.�"���$��ꐷHPiʥ"O����
X�ST���b�O��+V"OJ�jV��;Ba�f	ٲ1b�8��"O�H+��Q�`c���U������"OL�0Q�L$Vrxp�X�M����"Oֱ�`f�vQ eC���*8"O��A�LV)���uB6��Yf"OF`+AϞ���܁�AS5?t�yR'"Of����A-4�� hr�4H>i��"Or蓧	j���I��$jؾ q�"OB�z$/۹fV�i��ƣ�R�St"OH}���ѴN\h�lɱ:��Y�""O�x ��];<L*�De���Դi�"O.1��g��l&Ѐ$Va~rPY�"Op�� �	0�@u�#B�xMJ!۷"O������L#��ނ��u0�"OP�x�-�Ab��!7.��b"O��Cք#T]R�J�a���Җ"O�$h��=AT���ק����"O�-��� @��p ��2w(dP��KW�<x�m�� ]$��$�]"!3r,.dU�m�ǁ��:!򄅱$���%���6��u���!��U��X)��B��BT�sO�!�$������b`���
Mj�!��Z�㊭0��!z0��@g�6ce!�d)hj��KF�1QI�_!��HV��y�&j��~�ڶЇ�)rJ!򄉭@���i�C*M��!$����*��4!0�����Ov� i����铄G�X�S#�3Xvȉ2oE�(�4���(��'v��{Q.����?1�X�DA>AK��#�N�D#&�����O�3���3&�Dkt�r�p���K��d9�X�n�����M�3�a��/L�!ņɦ ^�k��kq�O� �J�b� &l�aPbO��)v�B�)�	  B�!~q��X��0|Z�LU#7u��$	~@URD�Ķ�\%R۴��dA�H�����Oj�>�#�6808��-�y�%�f�|���S�Q�R��Ҩ��Z��)ڧf���{3䌲r�`hphH�(.�	�����qn�	����ԙE��Z�r���$[���e�Opl���'a���r@Ϊ-��d�)Q�<��_�<��$*J(�<(%�tʰm!�MJw�<�p�&NeЅ�$'�"�3MZr�<�k�R~�-�Ƅ�5�P)��m�<�!��rp�|s�Ƌ/k �C�e�<1�FU�qO<$"�"�zy�0����h�<a��Ĥw�2ɚ��H2�H�H��M�<ق�Ɯl�6��'�]�mb�h�SK�<�w�կ@���ēN���q��M�<Qpc*ݕSБY/�iBv`
$�!���6L%��+,𕰃��)Y�!��~�JP �MM`�@G�\c�!�S�U]&}��U�bd=��LD�5�!�䈀d���ҬS�Q4�墳�}9!���6\7v٨�M�R0v�ib,X+$�!�U|^���ŋ�nI���Ũ�!�÷Y�Ɖ�Pb�;89��!GaȊ]!�05���1 �F
Q��.ޥW2XB�	�lN����l�.���oݭ]�tB�I^3%��E8*���A�b�'�<B�ɢC���l�Z`�-cEj
�KjB��"Q���eB]�)rl�)��H�a0jB�	�3���F�& �H�##HQ,gaB�Iy�(�%شEmDA �b��f�B�)� �١S�T;=�\i��5wf�* "O,,�ăQ)]�� ���0tY�Q��"O�}��a×�0��	&B`x@G"O���2���K~�ٺ4���+%��"O����ą95u�E��15��q2�"O���T`�/��Cf{�^D2"Ot-�0a�>wT��;�$�I#"OF58%,H�ew<M�w���c�NLˁ"O���0	5*
qc�
x��"O@)�%�_).\�Li #�$j�L,�'"O����d��7&4H!�T�f�Z ��"O�q��F�.�4�R���0E< J�"O|Y�'N�uf��# ]�K!Pр"O�2`A@=kP��C��͊Ne4	;�"OD�Q�P�|BH��5%�)kS>�""O��å�
/�}k��s��r�"O���0�ًBW�C�	U�!fPm��"On�Y�*ɺ4ppH�kC�e�%Z�"O�L�1�C�L��=s�� <��%"O܄����/K9v�[s���l� "O�0 ��1��!YP���T���r"O�4�Q��e�<ȪP��6x�� "Od�X�#ک\bu���="��[�"O$���͙p=���6s�t��'�D�2�إF�X�P�@�'Tl
	�'��qUiR�/i�0	#%��<c����'�ޅ37$�����a�_+ ��y�'��EbPΜ�e����l��a�'��j�I�#tU�3LGX���'�T	��.9N�}[�'A7���'ED�C��&2ɸ0�� �J��l��'��0H֤V�+�J(B����1�'5.`��-\;Z�|sf"F�Rza��'@<(�j�7yV��r��-�.���'�,ܩ�LA%�r�C<H{�I*�'M&�����f ���-	*?<���
�'��H����'ȸ�2�#2�vA�
�'�,	p%T@} ���σ+%����'���^$ip�p��N�Ј��
�'}�;��u#��)0cL-�@��'u�@0 �L1)g�5jg�G�#����'�TYG�
3Oȉ`�MQ�'m�P�'����� �9F��r@�k�v|�
�'�|��u@�+]��-J�Mլ^�{
�'Ȩ� *ͽ>ܞ�Q�I�^
�Y�'e�����>�aZGMR4J��'�B���G��ǆ| ���8����'�B��S��.||b!H�aB�}��(�'�v���	ǇJ
Z4Pq�O�{~����'/����4���A�oJ0��'��T	F�D����ԣm�d�	�'V"lZ�U*p�t������n��4x�'�,�%�0;Lђ9��A	�'40��S)�/3�>ۢJ�$?n�c�'^���UG�^�,c'��B�:�' i#�!B8J]�i�1�C�
�F�K�'��X�F/�/h�8YH��
��@z�'N���(~<}��ܚn�Ș�
�'�2�k�L��j�b��m�y3
�'"(D*K�%b���#�O�W�Bt��'Ҫa��k�<u�PX�X4U�}		�'�j�sa��ZS��Q��#Q�ҝ�'�|��,4Z��l��E-��'��-;bȝl=���ýC�d�c��� |L�d Ëv�6mC�� �f�:�"Oh���"J"Zj�bb��i�ɻa"O�9��7 
 �5m�� ��L�"Or�&`M32�Θj.���"O&	�1�0D��
�L��U򨌑 "O �t�H	N�i(�$ŵ1�����"O�쐧��z�a)˵$[���"O������t$��QH��qR���"O��0%N�Ro�,@��MYV|j�"Oܥ�w+ƃL�h $
�X�E"O ��H4J�#�R8Ui�"O�di�DX)1�u� �	��!��"O~� pA]�cV��GQ�4�zA�"O,�j�͟	 ���dd�4}*p"O6d�k�!Kz�I�M	|<Z2"O���IJ=b_�Ɂa�ɀ�V�چ"O��r���8:ʍX�*'���Sb"O0��'΂����i�=��T�u"O$���M֚e�q���S:.�@�"O"��0B���0�'ޛ:�)�"Oh�ѢMB�p5�H�G���%�Js"O��paH>I4-H�g[4]uح�#"O�Tiw��I\4�@�P̬�j"O�0�q
��o��qsF�o��9HS"O�� p�M�{��˙F�����"O|�!�w��0�� ӿU��y�1"O�Yh�!Y�j<�f`T�A;� �"O,p�&�:l�xVN]�'3��Ps"Od%{�G%�(��2F�-)f"O����� }�aRD�\�X�2 �"O���S��u�0��V��u����"O�����U��4S�
C�C}@�"Oj��gŦx�\(�hΑj���"O0��,��wq~aqG�3-��1P4"Oa���^�p`�E�{��	�"OV�FN�0Q�- SeJC��T �"O�aa�郂Pa&`�&��?VPX�"O(�
ԗa�����ހFg�52�"O���rד\G��a�cفb���'"O�8���Wa��QwE��܍J�"O���@ǗA� ��g��g�2|i�"O��B��Q�Z &	zQaS�m�>p�"Oa��g��@=M���"e��l
�"OrH!��TFD��Ȇ ��9I�"O�1����� a�����"G�f�2'"OJA�/E�&����D�W����"O~q��9~��2q��!�JB�"O"$�G%�s��4P�98Xh@��"O�+�`L?XEΐ �>>j�)"Ozt�S��I5�x@e�]� �b"O$dq�"S�J�!��i�E�v�"O�|⡭��;�r)��'f����"ODX��E�v�!xG�O]{�ղ�"OxQ��#>M�qВ@_�7���K�"O$����,p7�5#W�Ѓ	�;�"O�q�]�53��ү�(5~=`p"O��X'�X�;�����-F�	�8��"O��֨�s��]��!�^ A�"O�t���Z�1��aE��@��5�"O찊�a�:���X@� H�4���"O���oт�A9�`L3ƚx��"O�T�cC>}�)#���A�Q"O4�ї��R�T�	����%�~�3�"O8a��@�?p�Q�D��$�Cf"O� I�%V-3��"a��}�:��"Odᢱɚ�R@�l�7!D�x���"O|A���	9CйG�ˈ �)�7"O*��,�4	�Y��aX4e^`0�q"O��![�q�i��V�S>���D"O |�GA� ���a"��|C�Q�F"O�<�7蛁j�[��	�u6$��"OL������z'Ǜ�LT��"OjQQ��P�_�^) @�(?*T�"O|�93��?mk@\y0%Y�	�q"OF�hEL�'��ыF8 �j�P"O����6�:���^�jE�"O�X���:�i3�G�BѬt�"O��JPƍ@��xi�@�)��(`"Oα!"���M�H胠��,�α��"O�[u���$R���e��� �l��"Ou�2H��OI<5�<+Dr "ON ��bʐE�E�s� �4���� "Oe�a�G��^�£

��h�"O���lG�VE� � ,��$u���"O�:�	�a�����ËK�@���"O�P��[�|�80��-�"��f"O�D`Qk�%�(Ձ ��oи� "O���"I��ڐE�21�2�"O� �ea�0��a!#"N%1��ؑf"O��kVb��|z�+1AR(q؜I�"O2���#B,V�̝�Y�j�^��D"O�ɩB�6݈�[����{�E� "OxX�@�J���()#H���8v"O
(ʄ%��j� b�f�((�\�J@"OΥ�������Ӯ A\n9�1"O� s@jQ�A7�h!�O'�� �@"O�sń�Ev����Z� "On���(��`@S�\�Bs���"O0��V�hd}Qa��#M�:�K�"O�d4(]m٢�Ng}]hA�}�<�sǂ��
0��9$��b��y�<����3l�;�b]?"_n�#�u�<���� $��a��� �.\��ft�<)���(
���&�>iu�]�@�j�<іM��6�`]�T� 7,�
����g�<0G�P����D=tBnhᡉ�`�<�Q��6#���b���<P�hA7�Nf�<�#�i�)�7l�/PV�0��CG�<q"�ɒ5�9� V�?����z�<	v&���p�r�`�;$Z��v�<95��#r�T�W*5F��Fn�I�<�F�Y����A		;z��|i@�k�<a�\'�,��Ç 9P��p	f�Ah�<a�JL9�
�#�۬?P ��O�<�A�ü=�th�t���o;"��sFMo�<�#��J�,�v+�D��1ơHj�<��$�y\y���@S܉�.��li�tӂ��?�}����?��4s�Qc�㙑>L�z�'S2<*���)�i���OV����L>A�2�$A�-�&f���i�Q.�2�j�g�](d�0�&�E!�S�y���U������Gjj.���H+����Ollzu6����H��ɣ�Y�fˌ�K�vqC�a(D=
����)lOZY�Q�҃^�0���K$iM<�R��>Q�'�VeeӨ���=�O��D�i3�,Ar�r=h����#�!�'NZi�S�|Ӷ���O��+�4��6�Ǣgr������	eo�E���S9mY~(b4Fq؟,Q��V�Ig�W�%ptk��s�~E!1E:������L����5��Q*�a�b�����?�����?���ēT�	���ެZ!4��܊���؁Or5��IE�J��#c���pr����.WƟ�&��P�4�?9,O�	(%�h?� �xȅbC�����F4/�������ǟD��T�i>���H	:��a����ĉU�h��$ʭa�DI�R�;lO�����1YH�z��u�ij'!_$�l�b#+�?C����3��:Bw9�**�(�����<ۧ�� d��32Cø@�()�#��&xZ��Izy��'z��z�O^�U�e��C�E�ټu2�$J
�'�����3�N8y���'J�|�k&�+�M��4�?y�+����ܾx,6-�O�ʓ��	���z\&��!.vx2L���O���QPJ�O���1�I�3r�A%e�<Qsܬ	d Q}�O��5����� ��Q>A��L�[^�g�/i�&a��,�ɦH@���O֒�j�'n�u�p�֣0or����A�~�R ���Oޢ=�݇�x�B�S* �YX`�Ρ1M6������IX}��K���*�H^HNE�CN.��.����dyʟ��d�O���i�8}�E�T�/R��B�7rl3���~�	՟h+���|�S�,�V��@OO�:s���K�8���!j�<�6\�`�O�AD��O�!)'��)O�B�
$}Sd�P5������I���$U gK��%����c֪ ��NP��nJ#8y��Kw��=f���',.*!A�7VZ��)d�T=Y�Ў{��h�r$,*�?��S�az�ȓ]t4(�5t�=�����hC���Ms���?y����|r�4-/��Db�?C�}�]��)�)0-.J�(�'F���;q�bɋ��ޓˌ���4p;�E`�H[�O�}b	�z52u9��Q�W� ����H	N>t�m��/����O�%�<�I�� '��`���Ԛ�bQ�N.t3�*}��'ՆQ��^<g0�eS�L�~��؁Qm���'���4�N>�����0�O   �   �   ލp�F˸�x�rhK9�1�#l����_�)��ToڬrN�'|W�Ds��&�M3�i��P�E�d�F��FB*�@�J�O~6�I覑�	ߓc?F�KE�ַ1�v#p*�8s,Z�9lTA�'8�qEx��ϦIq4hF�w��Ձ��Ýo�,�b��<YAΓ0u��YH�T~�M�&a�l�"����|ج��)(_�f�O�jE�x�`�07M�8-��I� dh�
`�irr�����A'璩
�q��ƲLZX���h[j"�@����� f����X�'ߢ9{�h�2(k�J
>�
]�t"�*m�}j���B�I�"��+�E;�%	�B�	�LR6����4k�4T�$i��oj�C�I�n�F���F- �ѱ��:^��C�Ɉ���R��!+1Xc�6Q/�C�I�Vs��k��'M*���f��a��C䉃D~L��R�4}^�Q�D]�r��B�	��p�Q��ǘV����)zC�E�V$=y=L��dȫ^BC�	%X0�p�E�
2b����	u{�����!Ih����bEy�B���kT6pՆ]h6@��?y��&%A�X,G*�\�r�i�u�`)p!� JfJ�)Y#�M3�̘Ix(с��<!��Q�S`<4$����_�xO^3�LƷ2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          y  /  D  U  '   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=��J�E�TM�P������PŌP_`��7ju�r�d�O���<�'�?!�Ov�%ʢ���)�-#�E��-�����L9B8��	�}xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�z (PЩH��ɢ(�Zc���a&,O�$
�-ڼ1V�pU猤IV�u����B�ayR�BNj$����n ����ϻ%���OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O�����KO���O�<Fz�O�r]�pc�A�,�̨B��;W��)�1��jm4���?y���?)N>��T���GN��fg�h]$S�E�'*!���><`D��E|B|�f]�p�&��OnTh@�Ƀ ���S��;��L�Q����bi,�Oڤ��E?:���Aץ>k\�s�"O�����E�"��ƀ5h��×����'���e���M����M�@$S���ī�턙ZPyç	hBY�|�Iܟ �'����bĜ�$!DѦ@{u�@��G�Z��1DG�=�2��,�=��E|ҍ��NƤI��ןa�N��A��>(Ҹ���1(n�Q'�X� �	�i2��O�����'�@7�O�6��<��3�! �kUPub$�R�?k  ���,��䟨��\�b��&Z���T+h#�8���;n��B��@���P�h\�>ϐ	��$��>�RE�OD�G=���i'>��'Q��C�I�*�P��N�9��te�'����}����;��)��G#�e�R��-��`�)���HOJ��3g]�DF�YS��)
xѮ�3�ޏ;M�Y�'O^��'v�P����?����?ɉ��DT�p>�M��m���4	߂��'A��'�������(fZ�`�ʊ�u����ǓY\Q��rQ�:������/:j4�����	˟(�ɶW�t��ޟh��ϟ,ק� X����z5�|� , E(5۱矖n"��XSZ���d���g� ��)bH�/MªL��ЫFⴳO��2�X|R�
F�,��*##*�S�v��	$D�Bm���(w����t�@����&�'� Y[������dp�Ȕ��X�������aQ�LH<I�+�E��,����O�p����K?	�K웖fg���|��'�B�O��A�)��mIR��1�T��Ek�0�&p�ڴ�?!��?A*O�)�O��$�U\��
�F�t�q�1�W�Q\��5#װPm����'��Q�p�L�N�<M�&�J0��uv��'	��(Q׍�-~b����ҫR�4�3퉼"��h��X���Gwȕ��H�O����ɦ���xy��'�O�1`�5xq��h��Ձ����"OB��1�P�	cl����M ^V�<B+TI�	��MS����?�p������TG%R���
4.��B�$��?�M>I�S��򤙻G�4Z�'�� �ؔD�8!��ik�=�P��R�qЉ'e�!�d��U$pS'b۱'�If�w�!�X�x�-˗�V�_V$S�GE�Rѡ�D9<	ra��8=��,*�g� 5�H}`���Ȯi��>m���H� ^�4��c�0#6�d	���6�?	�°>����Z?VУ�MrcM���y"N��@5%�! �8�<��IR�yr$�@匰hGN2�~X���Q��yr� }_0:P�H�.�.0X��p<�7�	��R���q1� �F�*pd6�IK��#<ͧ�?�����kP���!�4Ӳ%s$��15!�d� ��أ9�:���`A!�D]�A��e"�-�+���C��G5d`!�	-q]��G�(�#� ��l)!��N�k�^IK#���$Y�f��(�����?U2�	�2�Н�3`e!���$}b��]�B�'Rɧ�'U�0a���@�r�I %c�Qv����d�E`Y���@��$�@L���.���H�*v�=�B�O1���M2V]�2�Uej�a�fIX��5��s���u��bt���1�]�i�=��ɽ%2���'W��eP��W�a�Z�pI�f6���IB��"|�'C�\t씙�eٖH���'�����ٚ���.�?�
�'.�TK���9���J�(L/��LY	�'p���̩A��nB�<��z�'G*�b��)��e���D�	B���q�~�'��Tc��i�#@�H��$�#��5Sd��9D�<���x��I-� s0�Ǘ(xX�2c�#�C䉗'�Nu�1��>�(����I#i�C�	���a�s@`�@�	�y�2B䉏=l��S�H,M�X5��� Q����ĐB�'J&qHt�X���b
*�ƨ��'O^9���4��d�O���h�[�D?PL$Xz2.¸2��Bڀň��K��幒�����ȓA�XSX7`d�1&�Q9p�@цȓ�8��g��*�� �Ƽ	A��ȓ,:TE�����ּ��LBR��p�OXPFz��D��$�Dq�E�A')1�@�È��	<1����ɟ�&���Z(qCD�gg͹ F0+�"Ox�[�&��Xb�uc��'5��0"O��Ѯ�4�t�hO�Np�0"O����G�N&��&*@!Y�T�"O�l!�OTe���N�i�d)w�DK�'�4���o#���v�D#)�D�86�� m��6�'�'l��Y��Ɂ�U8v� ���pf���Ш:D�p@'��(,S��s�#�z����4D�x�B�ң9M�mI'��=w_l� �1D�(xrN�T򔄁1`�*g����a1�� F�/�F�����k\r$�M4=�Q��F�;ڧ�(��"!�
m�z}������)��'r�֧� ���D�һ`JN8a'BA@"z�h0"O1
b���.3��K7@2C0|��"Ob}S���#V;�xQuOþz(�ŉ�"O84�M�!�Ti�##
V�1��'x�<�d��r\2e�1���n�Cw�O|?e�Tp���$�'�rX��:��*��˟,7��Z'�;D�di�lN�9���݉|�T!�
<D����
�Bgn.�Nb4D'D�h�ю�q9�܀0�x���g&D�,����W2�<�" Z��`"�*7}"�?�S��-$�H�Q�ݟ@��x�� �13����O*$
���OL��&�����H�F��'A�R0Y����y���1a�8���O�ay@�yReS�6��1�D.�E� �胅ܽ�y�J�%��pv��=>�R���@W:�y�^�Rĩ�b��/�r|s4�W���'�@"?"@�ß�1�)o>D�`FgK\��4�W�?qN>��S����U�3(H�ID��-p��eƚ7�!�_�yfh���6t'���d�k�!��^�2�� bSd@�x����i��	�!�ЀIЀ��!"�����$�!����h��`h�`�# $:�`TnH �d����9y��>a��㇧Y���BK#
6��u���?�����>�!��E��ى�V�2��� K�<����J�`�b�� �_�<���Ɔ!U}�X�$X&.�MG��r���YB<m��S�u:�p�㉧�(O�h�w��/�<��T�=k@-�"�O���Q�i>9�Il�'Gx���SU���#a�4R��j�'+lx��MA4.�RԐ�@H����'x.ЊvΈ��t��G�K8���'�R��I�
E�H`��Õ?C%��
�'����#�� -M8|�3�!SU�5�N�������3��� ���v�����( )���X���?aN>%?�!�C�}�� �h�3}�*��c�,D�aP��+r ���LǪh$�@�I,D��І�]�_4� B�)�v��|F�)D��0�B�z��/�aX�A�-*D�p��۴�<�Ui\�O`H���'�<��OV\6�' Ƚ��`����4#�)��a��O��O���<�`ac`Tyag��P������h�<��+�B9� �:@ht(�d�<Aң��� 〮L�v�֫D_�<1��H�t�Ќ���ސ:�<����Z(<���߂IA�|z���,u�*��K�'{��>a�X�O�I���a��a��� ~�L��@�O(��?�OH)4H�31�E
ìL�Y�m2"Or`����0^O�Q��Z�G����"O�]tcA	+ :=q�B�z4aG"O���,�h��E����.�>X�`�'�\�<��H�pO �hD�%?��Չ�A?��G�\���T�'_�X��0�׽p���j�DD9TZ92�+D�8�1�� ��A d��1�N��0G/D�@a׬A�@�eQ@|��Dg8D�lp��^_��`�u_�sT�H�k6D����٧s:(�%�O�ya���d�4}��-�S�'dX��h�^vRT" ӑD���OYS��O ��"�����1[�B����z�jL�1N��y�*PW�ƁV�"x�l��j� �y����#��q6k>:j��ֳ�y��;xI��`�#A��&�Z���'�y�+H"	�-p4�˳s�8�����'��"?���П p��^e��P��'//D)ȑ��?iM>��S���D�8�ƙ�1�!����W!�� ��)�Da㨼i�)�:���%"O�@��M&\��a�H,c�Bm;"OR�P	�<!Ш-��F�
!�p
O:�4	Q˞L��� H��mL���O�+G�Ӄ$YH��F��I���t|�=@���?��xt�	��'r <
����Q�������U9�n�qTeF�BXm�ȓ�Ρ	H�~;� ��[�PtdE�ȓu��E�F�	8 q$��s4z���	��(O��8�+�/.rP��E��y�h(�O��jt�i>��	ߟ(�'�ݰ��Z����Sc��'|\xpQ�'����׏�?.���U��3lk�i�
�'��=��O�/2&iCa�+jRT��'v�d�Iڸ
���6��f�" 	�'��а2*�T@.��L�32��PHH�����	H<��X[.ƣI* R��v��8l��K��?IK>%?��2���b�@"�Zq�����!�Q?V�*��Di5�=���5<R!���8�q���Al!�h�+�
.8!���G�@�SÐ�#X4�7�!�Dݐ9=�Yw
ܡCZl�ْZ��qO<�F~b�Y��?I��ς`�#�
��b]5�_�d��|"����	�7jެ�1*��`����m� e��C�W8��䅞3���؃+[/��C�I0����č�'`���G�;m�bC�I9���S�U"hohY�Ձ�W�B�I�5q
�����f�\R��(T6a@����a�@�}��[�c�"��D;4��B�i�~�2�'a}�AR�*_�D�R��D���B4���y�G���)�O}��w�O��yB)�97%L�2
��E�%r����yr�N�>�t�s�F7;x��Uϒ�p<)��	=܌�A��M�F�z8�s %@2��Z��#<�'�?����$^4V	�eJ��DU#�H����F�!�dȻd�TM0���8V�:�0T!�D�G2l�`#��'F��1G�iO!��.P�0(��0@����s@!�	����	Nx�Ɛ���R*�E���?���$¶"�& Xׂ��6d�`*"}BA�L'r�'$ɧ�'^-��j&*
�|�h� LWEy��ȓODP(��ݢ%���l�,���7��yIg�H�"��S ��4Wu,�ȓC���8��[�(�# .\�ȓ<*��%���;T ��r�֓.:���=A��I1W��DK$S�hq����7Fx�{��0ZӴ��	S���"|�'ɸ�`��:a4�X���C
�A��'0dl �!ZB;>���*�`y�
�'� PåG����
oE<�	�'6�5{Qo�!#T%	�L�/1�,��'d���"�`��5�Ć䳢�~�'�����i��y^$������K�P�GA[E�L�	៸��I�\�2���I�$�u�%�T�#*VC�;?*��{C�[u��cj�L�C�	�o7�=af׾c�H��b �/ �C�I"�r$d�#^� � ��ś<����$No�'t&L����O� А�`Ќ{���+�'{B�ي�4�"�d�O��#�����5!e�|$)��bЂ9��Gd�����El�� F'�)^	�@��-l�e�1�8ErL�e�-����
�� ģ͔a�(�=_��ȓe"%(À��uI���A�&Ѐ̤Ol�Dz�����9����1��~�D�v����R����şp'���
HR���l�tl����r4�tB�"O���%�V<"\Y� ��B����"O� 0��&F����a/�5|$t�"O�Uqcg	/S��qU�[�hnD��"O\0+S/�&(�q�o�M^H����PY�'��ɋ�7m.ly�l��j��]��$Qc�ds��'��'��Y�t�W���q����!�zԩWb<D�Ԙ�mB�nҔ�.�EnJ��7%:D��� 
��C&��S�U�F�R�3D����Ҿeꄡ����2�4�iS� 7����<WԨe�?X�Q����'�'G�Rٶ��3�������yub�qT�'�"�'oƔ��ط/ �0�s��*� ��'�n��pG�4�"���0u�(���'B�,ȵO�sG���$C��s�<E��'�αK"�JY�Ҩ��K)r���(ǓT�Q�,�ӬW;M\k� ӯi��f��@�'gE���d�O��2�2W�@��� LN�g h �O&W�Ȥ���OD����Z�g≥U�N�)���72z5e�N�yGF�"��P
P���	P�'4�ф�)�3��^��+E擹f�n,["5*�p��I|~�$(�?�'�HO �� ٨V.H�7DE=\�h�U"Oޱ�C�G�ZU£��f�� ���>Qs�i>U�	d}���2n��+�k���K7	^4j��ᢟ�8�	�P&��O%f�!v�6��Ҏ��l���+��V� �rk
�p���'��T{�
��?f�%R��[1A}��y�
[(c���  Y�G{f�b��'����D�l*�	Jce�#�b��aD��?Q��hO�b�x�C��Z����G�)��c�"D��Цo�$# �ɗ$B�e��!`�"�	��M+���d16�lx�O웦��h�����_
	�H�C�铧 �����<����?1�O�~��d�ϣm��US��� 4x4Q��O
v�ؤ���jW̉c�=,O�� C<�b��A� ���9���4��r&�hWo蒥a),O��� �'��\�(�e�X��Yh��H�R�%��H؞��-]���)sCG^t��� $��;���A�����������䌛nnu��Xy�T�X��i�'�?�J~b�4S��<�5͐6
��aJ�X.�0�'���+ �J���w�p���-�O��K�Te�[�Q�d�ѷX�B��U�3�ēGނ!`�Tt:X�!Dƨ�(�:�(�R!7O�8�TꐺD|l�;$�xB��!�?)���h�X6m�-G$��.�g��8���QC!�d�vNr�� �ʏF"Ĺ�7Ŗ'�xR�<ʓSi^��R��5|���QV�R.!��}���u����Ob��S���D�'�R�'��I���%Q�L�Ę������B(��&�H�!��L�g�I�O�R1ۄc�W��X�v㖲y��$��.Q }Vt�3�|i���xr��o�t��O�#.�(hEn��N�\�$/?i����SS�'y\m� `:}���dށU�ؤ��'v��R��/KP�T���;a��XQM�,R��4�L��>��%S ~��:��Պ&S���gh
'{� ��n�:���Od�ĵ<a��?��OP�x�Gl
Wv"�S�lM�!(Ta҂뛚M�
 !�w�`k��'�԰q!�
?7���5CӊoJQId��#�vp��mR�	���'�pؘ�A�f�� V��<r�2
���?����hO�c�8"L�W�đ���[�>�*�p�?D�XY`��&��X��{�V��qO
@nşL�'�l�C �~��4-Xᑀ��=�z��N�/)V@�"�'��	��(���|rq�A0)� Ib��Ú"��$��B�ʃ�T4�^�q@���way��4\[�=Ѐ�V�GE,��3c}Q����+�,���ܑ	���$]�5q��'!�	�m@�d��l�*e� ��¤Zs�t�p��I�]���#h�3V2ൂF3�HC�	��Zܺ�I<G�ԅ���3���V���ܖ'����[ir�����M��@-.�舘�D���)@G\�z�b�'���)�j�/u}*���4�r�-�@����C_�Z�$����˥O�r�!��
戟��z�k޷i��ӱ����TŞx����?9��h�x7-Qd����Ÿ]��%�1�с3G!�dC(��XC��
1�b8	Ta�+D�x��6ʓp�Nl�_*bn�C	I6:�!��?A	�&�$�  @�?