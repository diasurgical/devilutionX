MPQ    $�    h�  h                                                                                 WI=��
�.�]���Vm��/��H.r�BlQi&�/�-�F>eK��-��~����W�S,��.:j�9�����/���3���V�H��5��:�#m`�Y��[�x����$�x��Z)w17`S��l���;��
�/-�mۡo�kTKg��^L-P_Ob��4B�����H���>>F�ּa�E
,�'g�6�:�t>B�̱��N�o�6�$�#M�,^�"*��B�Ą���w��uSi�~��`�l8�<:~US�,����똟�O,ծS��p����J�?�C!��L�#j�
��&ƁY%��u��xc@}]���]�\��MOrz�+�� z�o#8z�v�/���a5I�p�x��O90��qH�#���Xbn�k�$�r|kY��U�1�M�WO�oX���D�P4���'+�����R��8����R�uZ����9��H�2��{5z^�>� �ܓJvI�bo���@�/��T��u�L�	�
%��\���Ჴ֦��������]ۈ�
*khA�i!��K�6�}]�u��� Ң�����6HR��kw��|c����B,E�Ӯ�A��!�z���^�l�����eK״$��l�(ʴ)������c��+NM(���N����`kv�*a���К�VC܉���n|P������O�8�¹0���d�d�|�b,�kz]@���_���3�XM��0٘�҂p=�r�\�%;����d��N/T��3ڨ4W��F�w�?�F�F'�iϙ�>^ԉJ�G�p�V��<�̙:�]R O:�����^ĎcLs^���p/E�H�DJň��U���2�L'�&{�f���x���E�Oi<Zp�\7'���g{6xbif�x�PT�(���w�*�Ƀl
�v_?";H�\���H��G OR"�G��xN!q�@B��_o����SϾX�e�r4'����v4|XWL$�PA��C]RP��dc��{��H�D8d7(��LDb�֒ �Tw��I��2���~ZI6v�X�E��*��n*I02z�_i��p���Wϒ�evd�|}��Ʀ��T5\%�ĩ���{��ژcn���l�W�:��<"TЀ��T����U!�P0r֮�_.F	�4�C{T��� �~��49��|�<�pS��.;��	vnk.�����c̆�{�����j�l��k:�GaЦ��%W˪��]��Yh�`|G�������ּSQ�,����~u�＾Xu;�Z�W�-�1q�出�tK�rSI�f�+��%��؛����A��@4�Ҝ����C5TG���T5���^n?��ކ�w{+V汇8��Vd�������!hn#�xx|���L�=JK�gbYL��?�~��#s����������zX�,Z,i,������X��S6�N��0\�I�[c�_�8�.�]l���Ĥ�F��yǷ^���,$W�"K��:T�|�]�o,�K�a����X�0D��2�=��k��K9���?n[���"'h#)��wV�7�H�^c�D�ze�e+O�C�Q�Kmλ�y��R2�W�T�L�GE��#�@r6�90���	�F
�v��L\�Y	8h�1��n~��k@<d����H�����Ztt.:��^�)}>vE?15��a��bKV�aZ,Y�f��F�J��0(#�Շ��K.��� 1�9�@lz˾�s�V�>��Ǯ���\���������L�LM΢�p�X��f�kN�z�q�t��� ��,�ӊ��"�-��<Z��/ܺ���m�*	�7��0l�)�{.�5��dbc�	���i����n����$؂Ŧ����Rŵ�ʒe������>%��k�<�nϿ�����r��krː�t�3�pE��d�R���u�ln�G� �W�ڪ�;/��fY���s��F'~�ɉ������\}�lZ�H�r��W���ȧ�\��*X�AA�a�hlݲj�6�d�(���H�Fy�T�F�-��1cXv�owdd>,��|M-ԡ0?V��HR�v��4��2�}*Jݕ��@��9��[��b���hǠz@Y	B;*���z����ب-�M�u�:x���ZGW��/T������!.���a�s~}�D�4�
*v�"�Dd��PW�EB3����>�@��{NS/�h����i�~x@7%���U���IP�b����4?K���S,��T���+�S 9^��UBb��S��i���JPv<d�/Ӻ�V8�Z�KjCs=�J5&�b�f���A���P���ά$�f�l(=h�>�D�.��ԁ�hz\���ѿ��� -�D� ����Dҍ_ ��,��Ɏf2�p�6U�OQ6�'z}C��;(����x=[>2F� 4�s����&�[�ǫ��T��4�4���r���.Pf��^��J��Z��a�ߌ�'�E�
�EN�ީ��\?��qU洁��t� S�~L�o����]lK ҧ&D	v�����z���!��:��ݯlr�	jY�ʂ+�_�U�Է�>C��@���bϠ�fExq�,zZ19-�e4��:����V(����=���t#m,�.��Nŋe����
�fU�����9B6D7��B���Z�u
��ҏfkU�<��_�x��P��R�D�R��%����.��6�
�������fW>A:&�qgdnW߼ߞ>�&q�,��X�{�!��2�ķt�*g��@C��Q���tP��(���*�GM��J�y��+������f��/�`���^��/V���#<�C�S��/I_�ee�-����t�
T`�L��?`�#�@�j�Y�(vC� ���3ٵ���Q�a`�6���vja8UW��J�v����!�RUl91� ��!&q>=�̵�_�������$]����(YB�B p����i*�����);��8ge�罦N�Ը�M�p.�ߝA� J��KDr;�t�����2����Ţ�p�A�i�2��y�����5��q&��QNK�A�.e_U�i$^P��믈&�� �s[���͟�K�*�U���U���������b��|��sz�s���#����M��? �c9�{����!��=:Ưٞ���@�zf� ^���\�bvi3�Km��^~L���"��ݭv4I㩪x!��GT|�"R�8jO�I�������{D=�ʚ�H��m�`�x8b	A�k�����96�>��$&��RdG��gE�16��Fty���L��N�3)���$���,y��*8��B�a��w\��Sb��٫�`��h88��:�S��ܦ�"�y�:��'�鮮>`p>������?���l�L���0&U�Y� u�3�~��،.}�:\�\Oe+�E�z 	j8��4�K
�i����Oap�<pCj��J^W�M�}H�V���6g�.E�F�$�'\|y��E1w bMz2�܊��������4ؠ�'��g��WRo�,�J��o���/����9���HTe��v�&^�8 :�e~��4n���=�j�xTo����	vH�%Tz���-�/-q��,��qp���Sۃ��*���$(��f�����u���$�x m{���g6�ޓ��^�k*@�ǔhɖ��� ��,��Ů����|p��5�q�����w�},���g��Onճg[z%Ѫ�^����&����Mx鉛���Ev�rqZ)��U �C�����GnW~#���Y���3�,����EWd��$b��Lz8h"�� ��S+	ڋ���pX�nr ��%�R����ж��N*�������*�̑�wl�F�����@��v{^��c�������<�:o�R�w��#{����cG�=���p�.�H�e#J@�	�0~�mg��]�&vƦ���vq�QuO�5��\r�x�b	�6s�i�/�T	C�?R�*���lE�_�)�;C�/�q�H<sB j4�"hm��S#�q방� ����f閮�PX;{�ˍ�a'd�����K4H�G��9�$"A�;]����7��sDs��7��	GE>b��� ��������8�~T�Iq�Xa�Y�%v#n���0��أz����	��2Pd&xd�����]�!a5g|��R���VB�s���)3�gm�R�:w�&���Л'���������!��0�kݮ��Fdw��i{o`�{�X���Y�:<-՛��&��Mj)N�����I=�V� ��u��;Z�fԘj��aV/�@|T��]]����;���Æ�A�Kچ�h��Sl�*��z~Pa���6��oɖRqɌ�h�B>}tf
rΧՊA���,޿��t���ꜯk��Nk���W�y5/ ��2I{�Sx�^i.��9U�2��+q�p���~V��<��c�nŊ��q��dϽL��\J�b4{��z�c��E�s���;�Mp X��HZ���zqP���U��G�6����0�ݐ2~{�_[	.��l�ߕ�?7�F�ʌy"2����X$(�P"��:/��|ЈHoǫ.K�G���JIX�R�0_�2�}[��F���C����iϦ/��h��ے��7�9�D�P� ��οnQy�m�4�������3;2�T.��G��~#�Nr��0Y��$��
_��'8�Y<`�h�p-��-e~6FE@��g���3�2���Q�tɶ���;p)غLE�8��	a'��-��<C},�V�2_�A�<JHF�����q���[`���@1��S@�����VEO�媋ԣ��Ah��zU�{�L�7�Ν�?�<>��ê����OC�Y|�)��Ӆ�c"D���p���`�6��m�Ά	��W��6�$Ξ.\��#�c���J��i5��4��$s����(8٭C���Q�vr��J�j���w8��ZPK��~���a!�&Gא�������Eh�6�T��1n�|�{ocȕ
K;6f��P�f4\4�Z�I�S��~���$t�׫�\�/FZ=Εr���A��4H�%�EҜ7���xh�
�j.	����c��ȡ�TFt�oޡ2���2{s��o�>�T|�o�<ދV�Q������1D�4-Ӗ2m��J�ˑ�{�D�Ʒ[�ħ�s]�h���@tLB��E�e[֑A똠:\�(������x�3�뷰�G��8�M;T��.�-�?.�X�a*u�}�=��
��-"��d	��W��3契�Rk�@<��i-F�F��l�i'.`x��J��"4���P����e��(���H?,���&.�vh9�ULU�/��n8y���)�%��<�8m/nU�Q&Z9�T��}�e�q�������A6�P��Χ�yfF��(� g�YC ���Ư�B�j\'3���C�P�-o�(�*$�,3�h��=Q]ǁ����c2(����/��j�b�}{,}����(5_�sW�>��. �<|s���ϡ}잢:a܏:40擶�W���^��_��e~�|�Ԫ������4�'���@d3
��șD��w1��%U������ ~G(�܊Q���K�c����v�a���@�A�,�K=�����j�)l��HjԠ�qĐa������QY��h�s�x�J�z�G�-lKT���خfUV#��2FC�J�%#�ʱ�>�N��C\|�Y>BfP��DhO���3DR�B41xZa���F�H��.kP>��$�xU�UP�eLR��R���苰w��./6Ƒi6��G}��@�W��Z&��d�$�z�>�.5q����K�Ŗ��2�Vt�gz�aC����3LP?�V(�d*M a��2Zy2���H�r�X����`����y��/�+����<2]���=�NqI�1pe �m����
/�gL��?�L�t�jJY(1b �����QP�`!� ���vgHS86��+���'�ص�gl�����!�zj=���Ю�ʃ4��T$��Q�zZ�#�Bi�� +Ԥ�/�y���)�gj7)v�82|���N�3Jb[
���*�|�����
|�DW�o���O{�l褵΢����m*���A���h��f�,�Űlư��?Ce:@��j��Q��p&]���~�[ _8�Hf;�&8�Đ�NT��ˉ��&���t�|� �z��͒�+��KK?ǭ�������o$�6<��������=� �����f�B������3�o����^Y�/�������v/6�x���oT��MR+�j*�t�1���N��{?�C�����H&`�r"b�~��W�z����>,H�r����b�'g�	6�J8t�H���nN����콄���,�zl*�x�B��n���w�8PS{N�4�`b�8S<F:tr����J�])���]�"��	��p����w"?|h�]LRl��@P�&YێHuc�Q�BhSA�X�|\�O��G+Ͽ3z{8��2���li��՟�a���p�{A�E����e�Hs�/�Ý�Xy��!��$���|��u��U�1�NM5-ܥ��������4��'a���[�R��������F�k����q*9�oH�N�qa�^O�� �����yﯙ��t�=����T
A�q	��g%Z�������Gʥrvs��!�a�~�*!���Nx�����s��u��s_�� �����H6�ĕ�~�kE)��u{����[�<,{���ł�ׁ���߷��昊bm?�Xsg�&����ו�b�G�,�i7���^��P�M�i4��ȸ�(�v�����S�C���w��n2'�-��)T�.S�梊��"�d��b"�z�v�<^Ư�.g�N)D��[��[�psi�r�C�%�r�2���Q�N%���s�ᨪ���pw缇F�bd��az�t� ^ʑ���Ӡ��v�<)Y�:�);R��ڔZ����{cBY�UB`p�8�H��sJ�1b�r}���"���b&q�B�:XۀL���}�O_Y]��\��(��ʂ6n�Ui���s�^���L*�=l���_uV;>H���XLH�a �6�"��.�q&AE��n����	�"X���˨�W'�J��5q4��!��<�z�ACƓ]ȱ��^��t��D�8�7^WQBfsbK7� Q������_��YJ�I���X��� b{n��!0��ۣ��%�f{����a�-d'����r�-5������9�q�N�]��O��M�:�ue��۝ж���J΂����!:��0E�\���vF�c�b��{�|���0���X��F_<�Y|��>��~�P8�,v'�Y矲1,��!^6�G+��a��a��䎨[������]ǲ���.������G\�#�^S�����&~+�45q50�M���灗���~t�*@rI&ϊI��g1�H.)�}F��r}F��P��U�5
�m]u��^d=R��CԸ�a�+��w�.�cVƋĔ*���!n���.�Խ]Lޠ�JAhbʉ���<�Q��s�Ķat�@�X��Z"�Uk"��f�O$+6�Y΋�~�����-}_�.i�?l( ���~8F��y}�וI�$Cq�"AE�:
G�|�Zob^�K�M͚=\X��g0z��2z	f�A����{����d�ئ��.h� �ۭ�7��4��D.М��[KQ�݋m{����3��HU�XPTi�G{�J#N�r��0�4?�
�/ܽ47Yw�h)ϔ��_�~���@{UO��>����:�<?�td�=��8g)3W#E�`��$��X0p���,��<�f��<]rJ���m��|��A�ߕeک15J�@��J��y'V�Qe#��$��ٮ��"o�Q�L5B�Θ4����*���O�pn��*��=l����Ӏ�"b���?�Z���m��r	���#����.�_��VVcV��<M�D���oR�$�æ����.�@F�&0�����E�ܲ���ګ��(+8��;ǐ��)��EC����.�on����co�P��;Q�[����f���s3��?�~��ݱ#p͒�k\���Z�sCrhD�0}�.,�� �����ϐ�lIh�W�j��U��鹞��<��Fo@f���h�RS��ƶom��>�1C|�3�׫�V��_��,/���4H�n2�j�J�!����\o��[|	��(h=�@��B1��@\=�|����#��+�>x\���ҩ�GM��T����յ.�:�a��}N�����
 %,"�"�dD'�W��3�R����@�X��Ѳ�����n1ibkVxv��ޚ��bP�Pn���5&Q��Z,7UC��U���l9��U���ݷ�_:=� �<ڋt/	�L44Z�Ɵ�D"��5��X�ť^�LAP��P'T΢�bf���(�$�t��$�rƊ��}�\��������-*B�6�r��BN�C�Px��b}��L�2��+��I3ȅ�����*}��]F(�k|�n��>�@ ��s�.�=�}�����<4˷��\��Ia��x��o���ꪎ��l������;4�
z���T�ݠ�Cآ�aZU��{�C�� �F�~B��7�C���-K6۽�epvxb� �-��%��X���C�%��l�kojO���o�����+ғ���xだ.�Gx��zP~?-GQ�I���IOV�q����z#���$�N{�h�~(����fK|���|���Dm�zB��\Z<7��`���y�kK���8x��P���R�����W�j��.�V��eb�?�(��W4�&���d�i���>�V�qV0T�A^�:/�±2�^$t?�)g�:Cߴ���YcP�6X(�o�*�Aݴ:9ym�W��J3�R&�S
+`� Ӕ�/Lo���a�<R@�>� �׮I�^e�?1�D>�q�

��L)r?�R�{�j��(젱  �Ɯ�w�
Q��U`�m���аv�F8��'�-�l�ֳi��KMlo1���!ܣv=}BB��o�����|}�$�ؤ����B� �0�J���_,�Bt�)��8���ݝN9���냦�9ߓ
c��e��E�_D����j/���%�'�y��˞�~���zz���C�C���ܨ�~���c��^��7�CeK��������Q�&��`�v��[;⽷�Lq����Y��,��5Dс����
�|�n<z�S�z�Ԇ��H��~�����4��,�r~=�!��P�v�If��>|��د83س#��Q�^4���Y�=�1q)v*Cѩ`��Œ �T�R�=�jJ��l63��o{:�G�P}&��`��b�ۿ�d��R"��ou�>�5��*�B��}�Sg;��6ozt��Ĉ��N��1�G�D�Tw�,�j�*.l$B�K�Zj�w���S��࢏<�`z�8n�:�3��~���P�pNT�g�d%�p�}y�)=~?�=���L�@��۫f&
ӵY6=Eu���I�3)�\P��OCn�+�Y�z֛�8?��c��MŰ��a�@py�:�@�j�H.V���$����fy$3�/|<�h����1-?ZM�G���N��u���z�4N�'����V�R%3�iC��/
����ȝ���9<�dH�*��l'^�n� �ﺓ����*墾O���� T�P�	��	,�V%����޲%:*ʀثT����'��yB�*|��蚕������u���! �]О��e6Y�W�9��k`2�Ǌ�y��ےԖ�w,鱮��h�2�T��<������s�3�*�a��ׅaγ]���i���P�Ũ��;M�{r�������v�bfm��ŉC-����n�Z�T�?��j�)g5�AU�Օ �d<�b�jsz��w���V�ċIG[�A9��Zp�	�r�%���mOT��E�N ����쥨e2��Xwb�`Fx [��H���^�E�X)��A<D�H:ec�R�)�����/��c=������p`b%HJ6��慲��e��+,&l:;���܀�����O�(�L�\�ʹ���6i�iwa����y,�5g�*|�ql�B _��;9(��'8�H�� �X["^@�	-qa��V&����&�d�4X�@���'Z���e��4�MO�)_s�XA��K]��������O)D��;7��=��b�� 8{�4����(�4`I�UX����n�n;�0c����s��������d�G������m�5�J���������)G�����v�H�J:-W��m���O����s�g��!uǵ0�S�FUFp8�{���q���s���<c����v�P��s�G�F�Ԥ�����\f���:�\�����ב2�v&���]�ʦ�
Bw1�D��_Ց�� FS�E߯	�~Ǉ�oS
��H(��B:F帥t�e~r��Ԋ���̢A��~��x~��RV�I�ŀ#���M?i5�1fѨ�#���z^_l^��Qf��;�+��Ƈ��V�O�e�/�5hn�衉�н�x�L���J���b�8i��
��Hs������Հ�/X؁XZ�h�0��NN��� �6�����~@�z����_Q�.DL�lc��u�F�`�y؆���|$^.�"���:�0|F?�o�0�K�s{����XET70�6\2��\�\ȁ�ːS_�ަ���hT��ȯ7�p�ToDi��6ő�DQ/�m6b�ʱ��ÖG��tT���G�N#��rG}�0��xZe�
U���O@Y�nAh�MT��g~�H�@6��aR���ޡ3w�t�i���U�)��Ep�3�?����R����,
��7���7EDJ���a@z�&����@�B1p�@=Y��~,�V�� �o�
�4�x���\����L�l�Γ�������Ī�q��	�x���_���{\�"��x��7!�����,\Nm���	6c�����8.���c7,[�@ַ���̪6$�e���}�c����v�A�5��z� g���Lϐ���ǲ���/��P��ؽ?��$�Eª�)��FR$n�F81x{�*d;lt��%�f����x1���~�)r��b��M�\��Z39�rC�~�k�ϧ�C���U�R���F"^h��\j$o�%�����o�Fj9�W=������o�z>���|�?k�r�V�s:�Y�]���4c9O2c�Jn����0	
X[w|��);h�D'@�=JB���}T��C۠p�(�ʶ��`x����G�C5���T4$��c�.�<~a��}	�l ��
���"���dy�WS�73�%�$�@�P����<�Rͦ�wi��`x�^��2Ŏ��P)���:�B�C��z¦,r��\�Z�-9o��Us+T䤢��ڢ��W�<��/��Gb9Z�Jt�*�����DW�9�A��P�l�Ν�Gf��w(CH�Y������e����\]t6�«~-)-��E�Q�"���j��Y(����2�[S�=�HȠD��s�u}����U(k��i�>C�1 e��s�{�ϗR�X�z�o[4f������_����r ��ihg�X!��]Ug�6$I
ճR��2��uȢ�PUw�@�~UP $@~=~���u؎=�KQ�ߧ�%�vS��[�w���7P�K",����l�s~jʗւ�����ڷƷ��ӻ��S��yx�9z���-"wDɄ~���W�V t��\.���s#�f��aaNV�r��P��fFc����h�j�zD���B*�Z����W��7X�kF������x��KP߭R�5�ά���=��g�.���G����v��2_�W�h?&a�d̼�\�>��Oq�w���U����2z�"tz��g���C��<��˺P���(�*C1�ݏbhy��k�~���0О��`<I�ӯy]/���s4c<�nS�ٙ�ƀ�Ip��e�y�)��� 
�y�L@b�?1��v<rj Ԟ(�� 1N����RʭQ�7^`W9
���vew8��ݫ4Ni�7�֎=��l
U5��Y!7�b=8������y3��W�$3���G�x2B�f ����e���Y����)�f88+��=+N�R��P��t��0���:��<RDC&��e������P��7��a����z�� T�J&����FtLآ�d��4���0e�uW!CΎ�R &e�1�[V�K�>S���������������B ���|���z�C�U	��c�����y���t<Ӱ�vĈ祍���=���OFg�5f��a�����|v3��v9u^q��>���jv%p��}%�MX�T�j<RpSj������q�{5��ʫtň���`4��bzYA��A���j�
E�>����(+��;��Gg�z76J�t*��eN�}���8e�p,�zV*��Bs�ل�H�w-dS�o��5`��u8�p:j��C��ۚ�_��Ю��(po���D#?��=���L�4u�v'V&Y�u٠:��sI
v�q\�� O�T+��z1�~8����rb�/ŋ��a!��p���;���^��H�M����Nn��@f$n�|�N�����1���M��O���$��J���4���'����qoR��B$	"�J���aȝ���9w�H%�S�gU^1 k@͓�VJ�P��*n����T@��P&	�Y�%��g��fB����[^q���W���t��*וl�U�������i��u���m� >1O���6�����ӑk{[���Ö��&��S�,�'���ɪ���f�����X|�a��.$� �X�W6�.��X��,�z�y�LM����:���^�bv�
Kk��ІX8CHr�m�n贾���*	9�$�ӹ�'$�P>�d2�b�zɟ��D}�����D�Nڜ6�ѵp���r��%����ZЇ��N���)� f�3HwݹEFS��Ut�ܪXT^�Y��ZQ�B�s<_e�:��R��;�Я+�ʲvc8/D��p�H.��J�Z����������M&g�������	��5OU/�+�\#Pf�3�j6d :i�5S�<������R*W1�l��_�w;4(P��7:Hm�
 ���"ٝ��auq�������g_����Xl|����'Ց�@լ4�(ьġ0��A�Pd]>����}�)�*��D$�7���8�b� �Ä�O�W�ĭ�I"{dX2����n�6�0�ͣ�aY�\�|�Ò�ז�d]ˢ���u(D5H���~��g�b���Z�����Cgq:�X��(x����@=хB��!�ق0{îzӯFu�����{����50�N��1%<����7�^�Z�Ҝb��O�i��%������}j��W���В_�������/]}��Eu��&I���\�'��y�S������C~ᩚ���y� �C�#ɝu�s�t���r?���D��݊��~�ٛs�YԨ;�>�J��H#5�ja����$�'^Z���J���c5B+��]�$fV|3D��NT�W|n��������GL�,J7�Mb��8�+l˗��s�n��LJ7�~?�X�,ZS7�����Ÿ�=c6֙T�A."�5�����_�N@.1/l� ��n�F��`y3aQ���t$y�"7&Z:�F�|��{o�#�Kù����X k0��2p�?�]��7����uHZ��@$7hX���b7|��:�D�?��э-��XQ�tLm�(���O��>��YIT�=�G��#�{�r�0�#�u��
�hW���Y�%Bh_�k��#s~G�@��ʳ ��4���|����t�s!����)���E+��Z��N���͘G,E^��/�2M�JY��3��A�
�7��41�ډ@�8��y�zVVH��7�%���j��7Ғ���vLk��ΎP:PkYm�}��"�f�������ç��Bu�v�"}���k����ʌm�(�	q\WY�'�
�.m�����cR"󿻏N�����:A$D񢦂�zپ~���y��\���������P�(��+����|����W�S����tIE� M�>C���Qn���������;�+�����fŹb��C�$��~~���5���,�\��Z��rNA����d{Q�xҭv^���h�Q�j�8TtU��'��r�Fe�޲�#���Ėooc�Y>��p|9���BV�4����b��4~�72�״JI-��,�I��N[r ��h��S@ŋB'�0����򟊠��4¶�Cx�����GC��s�>To����R�.�^na;9}ă��
Tm"|0Rd��W�k$3���c��@mh/��V�r�́��i�Ex�	M���w���P�-�U�+���U�",�E��T����9ʜ�U.Y�俇��U+����<P�/?�FB�ZJ�U/�����Nե+MAư�PU�Θ�(fW5|(��|�����<�@y��L�\�Dx޽��a�!-��J�l�������b���r㵊�29�:���!Ȼ՗��8}�_h�xk(���de<>�k  ��s��'�3���@9n4�o��������O��!;��J��D_�����Ѭ�14>
0����ԫ���`��l�UR6�5� ���~8Yb����I�\Kl5ʧv.���1O���#���tݛ��lޛujEò���E�A�o�auA��Dg�.�4��[x�#�zFKv-��ɿ����V<��C�{�#�d�#�N1�,�� H�*��fAjәU��%I�D�v2B��
Z�$���n���V�kATg�5�6x�7�P��~R�l�������Hч.��Ƣ����>��M�W*&<yjdZLC�K1�>}Gq�����pcq}'2UxQt�.�gKC����D^RPp�'(z\*�ie�j��y�Ԉ�<�.V�	eV`������/BV��N'�<ȼ��t���IIˊ�eQE�D���|�
�lL{�h?�3Uq��j[�1(b~� L�B���-Q�`�$S��nAvx��8A�W�O�$b���i1F>
�l�����@!�V/=�K�!�����2�Z$I�'U_��m5Bz� \�T؀�)�UT֍��u)'
*8�WP����N������vO߉u5��/���xD޽��`%��`�w�Ij����t�2���������(���h���O�]iʰ��Q�-r	e��U���� ��s�&nH����[qH᷹y����A�V~d���m�7� �N�|�z���0������~(^�t[���J�g�.�?D��E=�5�يR��xf�h�����Ni�3�z��@�^�gR��)�g��v ���j|�� T���R�j�mW��о��m{0�#����y��`O!�b��n��"���u��4>�tEփm.���u�	g1c|6%��te�1̸h�N�+�����ʈ�,媧*$�&BNq7��F�w�)]S���EM`���8�-:印�sS���x���z0V��Vp*���_)�?yxjh��LI���}& ѯY��~u�ZU���&�P$\�(Oy[ +��z��E8�+��d�'~�f,a\�p�p��62͆�ҭH�������:c$�<T|r+�{EU1���Mf�)���J�k�&�44��B'2#t���R�G����e$u��\��a�9�PKH�o��br^`�� &�C��ގ� �a�i��V5YT�9��� {	�I�%@�4�ڮ���6��6!���oZ�*2������>2����udjA�e �$��kT68���k���ǀZZ�`����j,L�����H��u=�!V�(#3��3!����װ<׻ԧ�S������J�J�G�Ԛ���Mo��u���'�v���Ɔ��ACc|A��+hnñR�ʕ2Ũ��m.����|�dM@b�{�z�GT���V����?���S���~3pĩ�r�%�Xs����"lN�w�]��۹�8�?wX�6F.����-��E9"^������J<z�:[6�Rg[t�ty�e�|c3��f�vp��HI*J,4����Y�%�Sx�&b.@�KT��}���jO�'��*�\^*��ϒ6_ufi-*
���F���+�F*2�`l1��_F��;/H���V�H(ޕ ���"TC�տ�qױP���K��RT�X'���_�'P�-���44$��_�< AT��]��l��;��ey_�D_�e7/`�3��b\�Q �o�j�����k���I]�X� ���+n��0�뼣�o/�׏Ξ����d�n���?�:5���0w�����~�� ���>I�:�yb��a;���һ���E�!�D0���u��F����'{ۉ��g�:�)�|��n�<����zF��{֜}D~��в����������R mr3��MMF��PJ��]XZ����Gg�%��k�O�T�@S�E4��#�~�����\BF5�>�W��
$�.��t�;r�a���������֛n���}7��ɰ�Y[�Cr	5���Z�࿦^U*+���ʸO�+�;=����VW7<���L��� n
�?�i�P��L/��J�Fb�v��f���"�ts�s§9o@X��Z�]����X� zc6�i\Μ�#��\��_G�U.�5�l٠_ī�F�v�y�[�z�$��"�ƾ:���|�u�o36�K�l�N �X��0��2�k�8�r\Ɛ��vUߦ�t�hʳ���5/7��@�D� ǜlv���Q��m�2� Y��y�
�T
	GLV�#�B�r���0E�M��:
K5����Y(�h������~��k@��^�j��5�W����t5�����4)D�E旜�u����1�J�,�K�m�,�-u�J�#0�E��\Z��Qf���1�Ү@s8n�t�V�����D�@8��ncK�ڜ���L"5ΉS��(!���Ng����»Np�����C�qN�"s%,�p:�1�ĺ"Y�ma��	�u�3S�^C.�y���^�cm8��6i�՘#� _ $ߜf�}��}�qC��w���ښ֮k�c5[��ꖫ�fk�9G����v%���ME�_��y}��|5�n��g� �ȁɍ;��z�f���F�i����~y	o��A%�Ö�\x<Z)$Ur�4��.���ăVV�!���Sh��j�O���O����F`"s����u��.(o�-%>s�|t�7Ԩ�oV}��;���4�(2Y��J$㧌g�@i�[m�ժ�JqhnR$@���B������-�����<g�x���#U`G�bN��T�l���(.���a���}0R6I}
��"W��d�}$W�E�3����\�@(�f��t2���\44i�xGN����Ǝsv�P����p���-�0��,��/��h�B�9%��U���ڌ$���?���t<�E�/���=�Z����nh�ѥ���?���Ao�P�WQΓf�� (���������.�\�5�޸����-[�󼇂N���Ի�)��30�Y�2����V��ֆ��i�}�å�WU(�_�_�>�D� ۏ�s"��ύ;h��T�{#u4��S��+K�Z����2�<�s�h�u��f���ߓn��,d�
��ȅ�H��9��"BU-m[��5� Z��~3T�H4��iZK��|��v	᫴ѭ���!�����Vеl��Tj�{�r@�|�x��Rm���≔Π_�*x�V�z��#-�"u�����	V����6R#�i��N���/M���L�f<�;�������D��B #�Z����2�h�muRk<F����xA��Pv_Ry���|��1���Z�.�b����p&D�h��W��T&��d��μ�%�>x��qgf�rV%�-����205�t��0g�mC�Mے�*P+��(:/�*9©�E�y~���J��L��dB�`�:��噚/����):i<+���2PI&�+e��_����W
�ՍL�4�?g��l��j�e(� g��|Q< �`�0�����v��8�畫j�'� �DE�y��l@"F��!���=� O�<�o�!�Z�$�GW�@���B��) �؛����n}��Q )b�8n����:NJ��N�h���V�� �gD!��|�Dyu}�[Х���4X�Ȥ!����}��Zl�YWq�Kq˻ޑ����J����W��m�e�+q�ÍW>+�Ҵ&ɨ��m[�+�4�[��ϸ�|m\�v$���,ђ9��	��|y�zwF�o�7�����o2��*���"Z]��B���=��e����G�f�
1�O���	v�3)@B�lh�^�~��
���gv*٩qv���g9TiKR5Bj�/ì΢����{+��a�c�4�e`j�[bp�HdK4�۴�@D5>�wg��ϐ�sw$�n�g�k�6 �t�զ�S�N����X3Ɲ���, ��*��B)4�e%wc�S����i`Ne8�h�:`,��N�{�I�A�1���uo$p�	,�zO�?�a�C�L>}3��~�&��YG�uO44ǟ?S"��\YO�C+��z���8p���X�8�A�"a�&mpJ��1�`�7�H_�z�/z�D��Tp$�|(��v�o1>�?M!X(�e�沮�fi�4�A&'͊��,R6���[���W�*�<qW9�<H[B��]9k^�� �A�솻#���y���3Tvw����	=Z#%�ą�&m#����ʬ�������j�*��B��)*���_[u?ېKf� t8����%6j��jlk�����<�;Ͼ�Gb",����MC�C�����Cw�N�����SI�V�H�N�W�>2���b"��oMJq�鰽2��|ovͺ�!n:���C~��c�^n���Nz`h�� E�R,����zdh�b4�z�(���'�:a��R�ژGg�pߩ�r���%]�S�Z�н�4N*S����-�S�?w�64F	���-��9^�!��ia�����<��`:��RB$]�FX{� j�c.���{�p��WHd�J���w�2���y��N�&]�L��="�8���/n,OKW�|I�\�$t�i36Z�i�>���2�ʑ��v�*��ll�~_�H2;*�r�8��H�E �~ "��՚+�q¼�':��]�um�X����� '˒���(4o?ь��3A�[�]��W��;�}�7�)jD�)7�M .*!b�x+ =;$������8��a�I��>Xhy��R�nL�0�BP��-�R���y��M�d�2�0F�P�5���K�9�]E�ںJ��M[���9K�:>�!�����"�v�6,Ѕ���!&^�0�+
�pM�F+U=N�a{�xk��Ѧ ��2�;<4��u�^��Л�����E�㲝���??�)��M�x��m�[�����vz�]3Ҝ��;.�چ��=s��TS����z�~��� n�݋|�9���S#S�鰮t��ir5`.���4�S}F��0�ijH�c�:�zx�t�傾�5v<h�Y�f�Z�)^P��� =��و�+��d�o�V2[�m�i�nG(��0�g�LJQJ-&Ib{E����*���Ss����������X)�lZ������u����6�Y ���E��7}6�_�.�Z�laT�F�F�1�y�u˕5V1$�%A"-��:v�|�@�o�hjK�����ehXv��0��2fw��ḿ�2r�$��Pa٦��?h�/��)Q7rom�f D▜���Q@��mg6����4%y�TU��G�ɫ#�)rXp�0 '��`�
�!�nc<Yc��h�����g�~���@g׳6�*(�2(�Zt�����l)�E�?WԐ<$�Dz5�,�X|y��(�bJk��x�w��-���/1!�@X�o�V�QZ��[���{¶���=�`L���΄�G��ib����\<�!v) ��0	�l�!"��E�+S��Lr��.m<�	�;������.#m��B��c�n���b �����[��$zhb�x#)�t�"�,-m�����|�|���Vܞ���a!���pA���T��Np�)���s�E��a�ה��n�e9Bu��<�(;����T�f{�|��H��Z�g~t�ױ���~!�\Z^Z�I�r��V�~���J�����c��w5h�j���*5�����Ȩ�F[X��h�_�>����oY��>N_|�r��C"�Vx��j����?4�� 2���J��U�����!,[h���:�|h)	�@���B3������h��AΡBe���GxH<��>�9G9�j)�T��4P�.�ca�[�}:��Q��
_"2�yd00+W$?f3�F%�)�@����M����7��iN��x���ʺ���m#PZ�
ËG:!\z��,#���-���9���U������K���l1<��/u:8�qZ <��g��쵄�D���A<M�P���ΎZ�f(ts�����j7���	i��\.FD޳�F��-�@��h=��(tү�3d�Ϋ��H�2�fJ�n� ��Wy��}eG�2W(<Fc�Z�U>T>G ���s=P��{���ܶ-p47>��װ1��<��ΔWi���?����~�	��.+ �'��
�Ax�@*
��ˉ���<U��/V� �$v~.o����ؿ.�K���'�v���مHT{��_�\�%�!�lLj;z/�MYķ0���P�������d��~x��z<��-��e�5�ص13V
#���y7#��kN�а�j�T�` "f7�ߙ诵��D٨
B�o�Z��Q�m���7k7X%��g�x��P0��R�{3fx�C�o�~G.�?��X��+. ����W �1&�Ld�n��:i>s6
q�&�-�����M2?t+��g���C��Ē��AP��(U@*�:�� ��yY��O5�ڊ���?`m��� Z/8���m�<>����:]�;~I��e�Ni�z0x�r�
v�?L�ͯ?�~gXHjn8(��� ��|l5���Qwį`(\��͌�v.�N8�1���qsX���y��H/l۸R��#!H�h=i�p�W�p����8�$�{�B��
��B0�� �r�ض&��K����ۚ)�t�8	����,N��	�ڃ��`��By��1MbDM��V�)�2k�<���js��c:]��2~��˶tBWv��J°��E�#�e��E˩���M���&$)r�b�0[�.%��&m�ķ^�U����%�����ĥ|)g�z��%��O�r��Ǵ��j)��_z���O�8щ��==\-�� ����f�̢���6�Ģ�3Dr�篩^��ĜE����v�~�̢*�~vTR�ǋjq?�X뚟U_�{&mpʼc��P`�5�b��?�u�>(��s>�E�9R3�.E���g'�j6�!�t�p��}�N�甁���@�,k*z�BC�F�w��S�����B`	I(8��k:��]�)O���W��P	���r�p�xZ㕕~?okH�:Ly� �GZu&�N�Y�6�u
.� ����j���\<��O���+��zBAt8+�7��F_�*aҐ�p���,�p�o��H��J������h��$�|�D$�q�&1�<�M��J�,W��a���ANz4:�='h���$R�ܙU_蛾|��=��+9(G�H�4��X@^Ċ ��\�O��SѾ�����A�T���"	��%� [�A ���-��"@Y��(��e�Z*�G�����[I��g�ul��� l���36�$��%ik̖A�v�k��Ԃ�,�������ី����t�^���������MJ���a�I�G���/��}�!��\�M%�늃�/��v�¡|uз�C�����&ny�@&��G�����^�ՁWNd�P�b�RzZ�ͼc���c��5�Pڭ�U�p�p�Ʌr��%8^��YH'�X\�N�*�:N��Q�n�GwN�=F�Wׄ L�{Z^�UK����s��<��c:Q�jR���\1���1c)�g�ZFpLI�H�>J"��R���⡨�E�&X���G���Ҧ�J:VOƦW��\�>�sK6U3i�rx�m�}�H!!�*莐l�_|t;%�튓��H�S !]"J�z�u��qM�\��D����r����X��6�/Z�'F����4�4�zO��)yA
�]oU��!w��;��dD�W`7e[@)�BbY� �&���_9�y�ޭ���I�
X�0���n��.0O����S�͒��T���KHd.�洇�9�n5y�6�f���ء0ڕ6��V_��4m:���Y[n�= tұ�q��R�!aТ0L��k:�F���	��{�l�]����ao�mI�<��Ⱦp�\�om��>I��V��ڢ�x�8�H���N��H@(�%�Èj������/]j����h��g��5�mJ)��C�S�)���Y~rt�[�x�4̳ɮ[��Dt��r�~d�c�.̎&~�O�dN�#ި5G,����9%Z5Q�sє�����~^Kh��[�/���+>ԇ�#SV���Q,��(:n ����邽�K�LeͥJ�%�bV4H��jȗXϪs����]�\��.yXD^�Z��~�,.�:��VS,6�i@�R���f2 ��_=��.���lOA}���_F��yD�����$�b�"�g�:Q��|2,�oi��K�K͚�[X1�^0t2�p��Z��(���N�K�ϦQuh@��4<{7���[��DU�������G@Q�Fm"=��6����qT��T�[G�]�#�0�r�V�0��2�I�
A.K�I��Y�=h0����9�~Xο@"E3�Q�p�_��]7c��tkP|��	�)�DVE\ԫ��ҿ��^�,��~�M$�#%�Jj�.M˒���&�r����1\#�@���j8{Vg�8*�vBF�d���I��x.TL<W��aC��j�(/��׿y�q�dN���#��g��")����Fd�g}'�֐m��	"�*�f�.~����;�c�ī�,|��
p̖�$T��s��������6���]k��v�����wͫ��s���˸��ԐD����"�E�}���Q[𲘪n�Z��	�����;����N�fV7"������ކ~oiܱF�>�9�	\:\(Z��r�̩�W]�5�ӃLGҾ��29Zh)��j���2�Ř��C��FV�������A�Qo�Ā>)h~|���ޏ�Vs7~��.��*W4υ!2O��Jڮ���5�v��[cl���(h�߱@6(B�����@���tѠ��
���sjx�2�Yg[G�u�5�T �����-.�gaL-}���l1�
�
z"��dk&W�X�3Ǔ�t�@�o��I(
��X1i�}Sx}7����8�)��Pַæ����r��5�,^�'���U��9�ZU_������Ƅ��Gw><�/�=3Z�Z[��`�6��@�Rץ���AwKdP&��ΉӴfh��(/7�����������3\�v�ޮ�rz�-��1��nT��kҊ�$��/iG�WB2JUr�)�F�IV�_�}@�mv�(�L9�U��>�W� Q�]sX,�σ�.��3���W_4ү���U���K^n�r0�^ꎪՏ��D6����"$�
A�o����~���U�6�j�  �l�~)���H��z"K��9��gfv�`�G$���������w��̑Tl/��j�Ђ(���2n���WR�?U��ըVx.fz�n�-�N��pC��P�tV���T
��� �#*��'qN�!{��i���f2?��f.��V:D��bB�JZ�����tq��uk2��F��x���PK�YRo3A�F�~��Z.�<>Ƴ3@��U����W���&��d�!�o�>n��q�j�蛼�!5~c2��tf�9g�AC�Sj�UՙP�+^(p�]*/Ӗ��AFy����?����]h`(���:x/��v�߿/<yg��E��d�I��e����������
Q��L,�1?�u7bLjl�(��� �f#��	���Q���`ç~��K�v��8r�^��Ӊ������:lvo���	!�R�=$�v�r5�e�a��7�$�ے&d��'B��� ��)�ѝ���p���E)�Y�8��}����N UĻp�-=]�����a�l=%D�D�Q�i�qYoΪQ�Wl��cw�>:���-���˱*����؎kT�7���e\a�����h�Ȗ	&�v���[�Qӷ*�4�H[���o$��잭q��H����|Du�zmɈ��P�ԭ��O���e@���U2����S��~��=7���;#�}�TfԮp�����V3_�	�b>^{最G1�8��vd��'��9��T9�zR�yajLˬ�(���Ca{!�������^`��hbf� ��yK��vÝ>���֔���2N��g��6�ytt\�̉8sN}�S�������,6�*�B���w�:#S封�V֜`�L�8�>%:V�F������w�����+��p[-���?���:L�E¤�UE&�iY��vu�G>;I�5�z�\w76OJ/�+�;z���8��RP�N����a�p��"�'����_�H���e��:�z�C�$Z��|C��lUy1�yM����Gi���=��Se4ub�'����R���`�趻��M޽��N9c�H�G�S��^q�h W���"7��>k�����DT�R��Sb	�ځ%q\��\�$��
M�ǵ({���r��`��*CÙ�A�[�#�U�u�@��: ��{��`}6 �c���Vk�?��_��f�Խ�,b�|QL�����R��yv�DТz���>׌��DFH�6�{���� �e�M ���&x��ʅ�v���ל�r�[C�Z��Y�OnTh/�{��G��榹�X�<�ed��	b�z5����ܯ]�C�0���l1����p
6r}�p%e��V���1�N�����u��Xw�3SF����A���^��)��3�.�<���:�b�R�?�����6��c$��wXNp�H��?J�,��-��
��$\E&S�z�\p��'N�e&�OA�2�K\yR����6P4�i>�/�(�  ���l*Ø@l�\�_N; h��t�HY� '�A"����Pu�q�B1�]�>��ӛ�+�PXX���J�'�>����4��!�0���Ae�]*�Z�<���s�x��D�7 �X$�`bmY_ �2������媭{��I�iX��~���n$E0
Pc�7Z��H���/Vb��6d�J���ݻ54�.ā"��S��pB�F<8���/��:��@���Xd��,���	H!�b@0�1�fG�Fፖ���{,���ؿ���� ��<j:�kn���D�F���2��;8�S��o|��h��C�����~�b�����l�q]�!|�1��8�̆ң��w?���S)���p��~MuG��ʿw�/��	�1�_X_t#m/r+���>�����I���\�_R���!��5���M!����5,�/��v��Y^F7!��y��O\K+.� V���/���Jn�Z�P�߽�P�L�i�J#E�b1CؤUZ�� zs�B�¸���j�X_��Z=w�`�u�t����6έ+�!M�;��_�d�.�Pl�A��|�\F�py�
F����$忳"#h�:,Ɯ|m7�o.kK�Ț_P�X�#0_�2\����V�#?&�Z,�Fc¦�%Ih����Oo�7h|R6�D��=�����Q�!Om݃*�Q`�*��/�|T�.�G�#�WFr]�0v�K�R�
�Z߽$��Y�B�h˦;��+:~���@ݡs�l� �P���P���tڊ���_)U�-E�������:���9 7,1Ӕ>B���J�Y�>3�X��#���g1�{V@D�
�e��V�Q��5���>����������L�!H�z�� \Y[׬Cϧ�Rc+�L'�����fY}�b�"����Z���库��m�_�	]�pŵe��.ٳ��ړc�:俧�b�fs��ы�$�_�n��*8���`;��}��r⥚g�����ϗ�l����J�#�C��_�
���Ee<7�*��Mz�n�oQ���Ȳ(k;�G��wiEf1�פ�rU��+>~jI}������b\U~�Z��sr��,���B�Йo��Y��}���hD�oj�:����� T���ܷFQ$=����0��oO�>�|%�Q�y�VnxE� �ɥN��4�h*2�1J��a��i[^x����sh��n@1�B6~�b��PQ�wu`���M*Mx�l�t �G/R`ߠOT[hͬjʹ.z&�a���}������
2"��ad��WZ��3� ���!�@Y%&L �|����i�z�x����
\���P�����}�����,���c�`���96fgUPK�+\��A�o�"��<<�/�@.(9Z�6C�3�"6��:���v�A�iuP��΄l�f�V�(��қA��bƬp��10\d�pީ_�]D-�:Ǽؔ���ۏ�e����M㡆�2�cZ��0�'Z{��J`}�>��(rsg�P��>
� ^�ss(���Y����$�,�B4mAѶ�s�k}�N��A�ٴ�����-�d���+
�@�ȶ���4PS��7U�[���n +�2~$Y2�5�K�iD����v��ƴ��*~ٶ����]W݇":lJ|cj1�\�1-�-�L�ͫ���H��e���ĲxI�Ez2eu-i�ɫ����b�V l$�E�g��#E��i�N������1�'�f-�ܙ��J�P�D[B�h�Z^�?����>�
k-�S��j�xrj�PfsR�
Oq��������.�YG��l������Z�WՏ&��odFA鼷�K>i�=qx�ύ�n��Kq�r$2�+�t�Og�LkC�̒��1P\��(�D*��?��	y�g���jp�f�u�.`�{�6:�/.�!��2;<�5+��E����I7lye=����E�hh�
,�SLg`G?8v]`j�t�(N�7 �<ir
��v/Q�l`^���*4v���8-%髻��Nn4��@�*lFt���v!�;"=��`̍�a���#�V�$5֞��N� �B�O H����4��A~��dO )_8?J��=�N[O��*�H�\�u���BJ�MDJ\��L�e�����`|�rz�`t&�Z/�
I��Qs�ˬ 8�I�J�)�ڲ �e7,?A�(�{��7z&ډ���p�[ݔ���S��#��-��� ����ѣ�C�:3�|_�Yz���qI��P���v�`w��;l��S���n����e=���vjF���fϰ��`$+�:\	3z�	�ݞ>^V�����q��*�v1>��[�����TT�^RxL�j'5g�΅ǟ�H�{}-�r)e�`���b���Q������3�>�@6��8��@�^�gE�6��tQ���$Nx#�i����+�,Q��*�<B�<��pw4�US�����v`p�8��:��;��ʉ��I���������Np���ˁ�?e��Գ�L���}qM&�LuYX��u��iV�~���U \�֍O�+���z�S#8�~m�A����ҧ�aH�.pw��"�%$�H�T^�������b�$�Q�|�ݒ�gEh1O�EMR���b�r�W�O��w�4�"	'����IRG�i��1��ؤ�Ȟ��̀�9��	H,z&�Nk^�.� ��=?��J�q���B�{TG�/�뤧	NKq%,ؑ�w汲axʢ۾���^{h�[
o*�^5���j�>� �Њ�u���ʔ E3��G6{����l�k	�lL����;���A,�@��w[�T{��	���3]��Q��U�q���'�';��?�z�3��6_H������A�Mۆ9�a�a�e:wv�2�2�(�-�C��v�ԡJn/僬�6�1g���c#����d��b
z'��ٴ��X��+���c	m�x�p0j�r�[%���τIЎ'_N�������HR�jpwD�tF�3��|RFܱ�J^�$�z�|��m<�3�:G\�R�>8��Ĺ��l�c*���vp��nH��Jq ���Ean���&N�����H�i���2�O��f�\Jӯ�:��6K	�i�;����e��*�� l_��;��I�HI+ B��"@!�+Jqò9��U��>���l�X���e��'<����<4 QH��Ό�S�A��]�vr�W\����qJ�DKD+7��h�zb�y� n^r�օ��o삭V��II]X9C���U�n]o�0��R���-�
״�c�dd=@檕��S�5���Ĝ�.�κ��Kn=��d�\��*�:O?����1�sȦҧ������!��0����at�F<ZCM({G�S�ަ�E���t<zC�ff,�%<��L��lΚ��%�.���7i�8e�>l��U�9D��%ª�s�]��c�lU��
��1�#ŵ�@�SDƿ�뱯~(���Ѩs�#�*^ �d,����t>h�r������٩����Zv��tJ��D8��3{�/X[5g��
k��+��^A&��H��
��+I������VÆ=��
x�^��n������<u�L�%�J��mbrX�R_���R�s~���� �%n�Xz�JZ�R��������U6���{l�܇uV��_3:d.f��l�ak��F�"�y���fGK$ =�"��J:��|�bo���K������bX�XK07��2�Y�夝Á^u.��)�A���h�bF�j��7�2���D�E��X��gQQ m���lF]����
�T{}G��#ޞ5ri��01�(�{v
7������Y��hf���=~Q�@�����p�n���JZ�N-t������)�E�����كҵ���R�,l@��V|�U�J ������B,�G.�bD�1��K@�v��`�'V$b�S �����Z��~9���7LrT�uFO��^����&��'Z(�J���+�]��"���\��������zm�=�	��`v���.4"�s��c��D�"֎A�|�0�$K���i��م���]�H���B��,�B���O2i�2�d��N���,[��lJ�zfҒ��E@��e����{>n���S���m�;�8��Cf+��28��+��~eI���~�ͯ��\p��Zz�re�͎\�kqÃ��(�t
&��qh_��j��t�;/`�yKFL�8�y]��o�OK�o�ی>�]|`�B���Vi��{��	"4l;2E�2J����S�8�-[Y�ŪK8_hZ��@L�B���=�Q�M��� ��� �xy�i��vG�NM�,�T�o���.u�a �}k#���w
}y�"��d��W���3����*N�@�lA�>����ni��Ex�����b���P�;~�ܵ��h�/`,����$�9��U�I�F�Q⼵���H<wR�/F�)gZ�.���=�q� �[Y�A��P\�4�%Tf/(���1���E
Ƈ�7{�\�7+ޤ�(a]-G� ��������@�sl������2 ��}��B���U�s}����F(��K�.>e�= ��ts�D��y���z1J�g4������c�]����T�ت��&� }�� �d-
���q�&�OB4��76U�@���v �[%~�Z�����?�K�F�yH�vu`Ŵ��̘���+�mb��BӃleD�j�|Ղ�k��h�&�h	Γ�Y����6�K �xdc-z�{S-D����e�؆+@V�G��
��"n�#`;���Nx# �>��1[�f(m5���̡�D*��B�Z9o��ʏ�/�k(N����x-G�P���Re��W���y6�O��.ߖ��i̙�\M�Թ�W�&�d�żR8�>d�Aq��T�^a���Ut �2�ht�'gR,MC���
P�(�C�*%d�ݱ�y
Kˈ ��ڞ��T`��m�QZ�/�Ǹ��Ŷ<�#�{�w��I���e���������`
�L�Y�?Ӗ�X�j"(s(	�a �2��87�t_�Q(qV`��	޾)�v?��8��7�ִ�r�ְ�Ge�l�<���}*!YEO=�/̨���[0R�y��$p�\R���BAޱ Rw��ڼ��?9�)N�)8�?����N��Y:1	�ca�𰇮��b��}GD�q�G��'N�D6뤍7�ۤ�����E����#˧�|h� ���D����ed|�ô�����&5j �\�[��G� >��f��h�<&���iB���d����|z��zc�Ғw�f�#��ǅZa�[΃�������tYl=��ٱ�U��f�� ���u���3�r�XF�^1�����n�vX���0ůETo��R�>�jw�	��&mQ{5v���!� ��`��b\�h�>[��;�����>��H�J���_n�:Ckg���6l�	t�b�̿�Nsqf�Ĩ	�q�5,l{�*��PB�����w��S��s�'�`:�8+��:L�<���5�|��b �c���<�pф���'d?�G��L�L*�!���&���Y��1u;�XqKY+e0d�\핹O�\�+��zSK8\c6�(=D�[ŭ��a��Wp��.�K����HK���V�0Mw���E$�&�|yZ��bU�1�
3M���}����H��Ҽ�4��'9i2{�vR�+2�K��e�C���p�9٨KH�̥�I�^'�E ��q�Xg�uc�L/��}�&T�9���	���%�s��F��ׯ�}!������7�VF#*�q��Y��KL�u�ޯ7ע ���}N�6�w��VRk�j��X���~��3�I,S?Įr��ᯌU��E�����:���0*����¤}�:`)Xp:��&��^��[�6M�x�露�� �v��u�Kc��hFC��O��n
���n�̦*�,�����ղ�adԯxb�Uz�n]�������&�ھ��3J�pK�Nrsߥ%��6�
��)=N����K���<4�Րw���Fu�݄��!�L|�^��:���e���<�]:�u�R���2)��lX�c���-��p}�H�/J�����陀��Z�Q&I��#k�$1I�^DO7U���\�M��We6F��i�Ϟ���o6.S��B*y�lXGl_M;�;����H��j ]�"�^��?�q�Bv���#���"��V�X���ˀ�+'���b��4[�f�Z�.A��]�7��r4��injL��D��76Dq�b#�� )����Hd��g�1yI���X�b��A/n��Q0���m���>����w�9 0d��n�L�J�5�Vkķ4��Iw��&�T��e'��%��:� ����iЎL��"�߅dץ!�W0�9�\��F�F�:�r{bu���D��p�S��Z<���a~��S����ǆ�1S�	N����(��9O�9?�����3jT�b\[]����Hnf��ߕ~2���-�S_��f�~�>���I�J�%� ɿ��� tY�r!�O��7}�?❿ 3/�U�����fs4��9���!5�_��E���p�^<5G�l6h�ů�+d�ӇAV�*F�*����tn��9���kL��J�Qb��Ȥ��Z�)Āsyl��n���=mX�SOZ�q�-����"Ÿ'�N6�Y��c����eq>�_�/�.A.�l �0Ĳ;F�]�yU��!-�$�F"ɫ:�E_|��o:s�K��Q��vXb��0RO2R�������˪��G�<囦b�Rhq^)ۅ5*7^	h�=ND���s����$Q�8�mSq������ �`�^�TA�GS؎#�ar��f0���9
��ڒCYO�hD4��oF~i�N@S����.�&*ޞ�S�[t<M����)��E�k�����0ļ�,���t���J{ȝ~����L+���=A�1�u@z�[�Vxe=����������Y��)�&L8�p��r;��ܬyo[�H
S����=��$��X�":O�����~x��m�;	����V�����.�z@�.x�c�Ϳ��u���G�	$�ւ�d_W��T����A�hK��#܊���;����2� �r��a[�����E�᠀g���<n��Y����(�;)T�m��f��r�mW��$u~`i��W���j��\�"wZ��r@kô��iσ�����T�c�bhz@�j��q�t��v*L���FGp���X�*��f]oE�>�}|�˧ԯ��VdZȉ֯���͵4 �T2�p30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��} ��UWP�Hh1�;�f��l݇�Jߚl�.�u?W�������Jd�WT�VEk_+�o�y�wϢ�w�Yc$�����^�l]b���
_��Dd�3ٱ���k	�9%]���^Al����}���V<�
=��s�'KK9�#�~v����B�I<���[�z��!������c��D�P �=�����:����e��$^�]�]��.�(� ݿ�E�o�hO��z�Sp[�(�혾��K�Ǿ)J;ǜ�zH��z: >ߌd����+|�"�<�H��l�
�M�tc��X,�D��e�b)��n+yL(�f7X2E�3�.�/���1��7��؈MsQ������{�+'|�.��C��@�7_����i�)j��{�!� ۷͖ٳ���U�!�0��\���� rbExy��⵭��T�cUc� �'�a6&~lx/~"\�&���+.G�����k/�~��<�Q�]���/�UZ4Dn��&]�\ֲ	0���+e<�6�p����ꓭh����@��#c	��N�
N�p��Z�(��xmW�wyM��({Cn$�]x�I���b
�^_�Izmh� 5X��.��,���$J�K6��\����ᡊ�J,+%��� ��^�����Brn����WwJaÍ���>\�D����Kq�Ţ���c���"��Y�P(�=�q�#�2n��M�I��6
���d��!N_W�q\[���#AC �+�n�K�PDL�������㳙���/t�]X5Q�����K;�?Ч�4���\X�%>��f�$X�9�}���u�I�����I�e��%1���X���ь �v�����]����iC����F�c���{ֿ-�����N�f!Q�\������8�qe�ϱ	}���DT}u�Rf`a~�O�R�a���tI��.>*[�y��t��Tq#f�K��Wxy	����Fa��)����86P�Y}X���ݍ�s�g���zB����R��C��70,�ԍ�h�R��_��I^��g�Ѻ��fH��N��,z �%6�t!u�K�!g�A�l�١�9���/�A�G\s��t��~u;�Kp壓��[.�/�V�Aפ��Io[C���$�z�k4f��8X��W��5��(t���۹�nl\�4W�m$d�,���X�c6Z��(��MeT��+�u��;'�;�:���!�(��+t�(|�d�pFV̢-���ʹ��JS~L �� ���#J�#��A�C,�,�*���S�ӟ��]�� ����mkVQ���^��N<G+#'���b`}������K�V�=o;�WOhVp ��O���f�Q��y�qk�(�6��)2���K�}�뇾�č�C�qռ��B��
����
�Z���}�K`BbOBlN��bWw���D5S
�T�oQ�'�X�p��dÈ��KW|7�\
�֩�+m�Lv�1%fm�"d���	5�u�1O���	x��jOg%E1dIv�Ҷ�VW�^
�j|��f��h�������SP�3/��;/�r�[-�G5�]���k���X&e<a#@�=��4���	��rD�7S�?�x	N����	o���$D��ߞ@�3�r4!�Ť���c�#ӳ��rT[�?ο����`��Ր�P�Q�¡WZ�6T��q���^Ck�=�+&��v��LY��_���rkw$��ʇ
sc�1t��n&\~x䦀8��[WN�F�T��!��ps����Un�p����AM8�g�A�r�����t�y�q�����f��IM� ���RAKkˇJ'j�q����ߚ�?�S������)4�1U�Z'?#�,'��yh(��T���²M�4${a٭<����v���ˎs��ǯ��!F�x=�f��R�x�̳D�J�㎿J�s�������؄�+F��h��q`�p�-��|짽����v��R�1Ŀr��z���dyB;�q#����c1'zݺ��<��_�`���L��B�a6�f��T�� �����!<*�7z�H;�]	�kS� N�OiMe*�k-��^A��.����b��^��W �iD)<�Ԯ�;Ư���|�C�A�DQ�����������H'�:fPs�񿆃C������w�6T�/�P"^��tPa6u�G��_A;+��޸ދ�1��ۯ⧨������c81�k.x�+���_DP���[��s!��%$�x������.I��ň.���:-�w1�����$��)up��^��J�觭��W�I���O"�4�������k�^�[�C�3�p���=xw�*�<Yd�٫L>0!* ���˼h�����	�EL� ^ �{J�Z��s�	�������J��nW��V��&_������Xw��~$�üHl��!��Ha_�ϵd"h�2�~��9���>ulڅH+�Q��K�n�2ƅ/\'!}�9_�e~I�P���?W�a���Ɖ�3��N���Mx��� R���x�����łe>��$q�L�к�.�q; #�E�q�[Kt8�szu�[�&�|"��Zj�~�{���kǏ��Hk��z��ߟ"����+O��o@M�L�����̠i��{X?j�e��b�2ԡ	Syߚ�f*Eݖ?.����$�>��]�s�9��x>�{�3�|m.��9V�n@tf_b	j��[�)�5�{�l� .am�I�ߌ�*KUV����d��+���U��y^?�h���gn�Uy�)�^X'�Y*&k�/q�.�y����G���L~�Q}<���]���/�i4� ���9��oI%	�����@<�������Aح�QV�l������	:��N~��ۣ
Z����k���Qږ@P{V�H���#����f���O�<WohܛR5�=l���i�KKy����~�8`�H��<(����J��0+8W�Vc�1��������O��C��J�����\�����b�~���5+=�	������~(�qP�\2AR����I��f6�� 
l����_j�7qυ_���HC3["���Ku|,Lh��C�|��$���/G8�Xhg��U� K.SB�������\*F#%�1bf�İX���}����'?I�����x�t%�=�+����x�	����M����fɝ��G}�c��h�u^-R�5��	ԜKQ�]�� ��mZ�����g���Z���}}ȅ�fe��bdG��g_s�D�2Ԣ*�.s��2����f��K��bx�~��z��O�Ja*��� ?8�o����<�����:������h �R�3�q���8u�(�$�an�R���_��^��1g�X;�D̮�˳a�%,�ڠ��2tM�I��x�g�Gl� ��K����A��F��t�0�X��>O�D/�"�AJ󭆕�d�J;z�ʗ���ΚQ�����IGZ��(���n:a�c��H�m�+,+O��Z6-E(�M��`��@X	���ZMcI
���M�py���ʹ��^��V]&Pe���~r�i�����3�� �\��ڜ��S������!G��`��S��l�j�h�������n1M�7�6zP�����/��'+K{��v�[Ã1��Dǩ6�&�a�H��gfv+�nip1#􅃢�o�@f������]��4���ؐ��!�1�P"�0'�������ٍd],�!"�"R/{�\.G�f7h3�Q���gO�OC��rs��WDܻ eG�@7M�~<�zI�: ?��۔f��
��D~���IO���^$��&�U*���ы��1V*�Z��_wbS.�����:[���9؃��װT���Po���ÙG�;�Sq�p��=�9���E�Ŧ)	b�6���9>�e�]a��ta(RM�
3��i�9�Њu3痂ȓ�;����z�  5�RLx��,zd}��P��ˈ��#��Z~��B�J0® yC��:����U|Qd�>4�"g>�q�g�yJ�C����K��:��TS4�T�ޒ�)��W[7��W`M��qSu$��"ԥ�:dtj-<�n�#�`K��U+�f3\Q�tX�P0=�J��-����K������yC�ӈ�����L#�����k���+��5p}�����Q�Yq�f�ͱᐓ���b��+��B�1���7�ޢn\�����u�?_&�?��B�2oU��xټw�n��ZS�奀�(�uw��d�[i�uջ��@�&�e)�l*��A���VÚ�J���Z�F'�Q��"�+]���y;Z:�g��(�G���h���Wޏ=��l�vP�	�3ir.�eS�2(��Z�B���-����ؿ"�@]��rE���E,�F*{#}GV�\]���e����
�,���P�G�,2Z�ԁ���q�=�^� *=�
�&�;�	��S����a�ka�b���0s�&t^]&F���+8+�nW�g��>�a!�s.G9���Z�Z�q��%M�����}�\�Y��H�@�q�	E��d��`QM ٨-Z�+��_<'Ԅ��;|w��z�?1��kx�OZ+4|�lU�v'��,�|yR=0���:c;�\'�4����(��.j��m��]8����I6�Fl\��PR��v�6�*��2����s�z<�����rG����h����`~#!-�������JC���	����1�zy����&B%��#���ͥ(z��5��s�����9f��5B�����T0������a����^�U9� x8\i�m�*��)A<�h. �E�=t�H�WJi���~�c;�ģ�/�C9�D��}�|.`�[^V��'}dbP]����0CA�t�l���a��T�pi��m^f�,PK��u���"�A�#A���;�������Q���ք����xH.��pn���T��[D����%Nӗ�+�����lIɒňX��Ѥ�{�!�m^~��B���Yu�	^���{у�X�~�"�"�Y���q��^��AC�&lp'������#Y�@��r�W0�TI��:��z�%�Ƹ���� �D}1J<L'�+����1�@�t�x�5J�w�Wq�VR�_����v&�ll�w�V�$|[g�f��lz����^_�hd�jv���	��9�1�+�kl��U>"�R/0���o��'K"9��~���ݠ�j2�UXP�s�M��} �@b���~ <}�����-Ҙ�,e(��$���:�t.{ �C?EA  ��N����z_��[1ǻ�u$`�6]�h=ž�����H^1zח���a�+��O�Y��v�&�n#2�J�n �Xir���Hb��mԋYy	wrf�~�E�%�.��g���o�~D��U1�sn���{<_w|��k.��� v@�6�_������)'&r{%b� �'�3�͌ �U�HҖ��#�y�ƭ������y��RƫÑ�,U��QP�'Ѐ�&;oG/�|�#u�ⲐG��������<�=�]�Oc/8��4A�������>	��ʐ�<ý��-�]�E_ޭe �V���<	�o�N(�0ۍZ�rf���
�t&q�*l�{�N��D��ƶ��ڵ�����Gh�z 5������)���?�O5<�hV�����(��ទJ��|+b�"��"����b������y�,�o�iJ�����3m\|���m��h+��_��q[������M(:�fq�?2��j�%I���6gqs�rW�q�_�:�q9�j�C1�+t�K��L�x��-v��/i,�/�XRr�PK��~Ф0O��k�\T��%D�fb$�X�'�}�})�_I�����y��ܷ%����F���G�3�������t��j8�>ı#�cPnB�^f-|�:�շ~ժQ��ːJ��ׂk��:�����up��TE}r�ef���ǌ���>�gGT�Q�*I��X�´Q:f���K���xV�����9��aT����)�83����D��P���C��*������.�RK';��ͮ��R�ƍ��R@=�_�v^�T�g.��6��K�e�,W=(ˢ��t7w3���g4�-l�Vع�U����IAe�[�H�t	ޘ;����堽����k/���A����?}�K��t��B��hi΄ﵳ!=l�����p(�Kaɘ���!�1�Vm�g�,U4{�5�6��(�z�M�2-����E����csy���e�[������R����EP�	���U瓧�l��3e��F���Ͻ��z��!1��`�7��bUj�^
� ���&�nkZM?�6d`&������z��*g{k��@�݃��q�6؀���H�;|g�y�X�1M}��J����)���=]�#��9��<N�[*".���X�B��w�9}]��O"e@B/esP.q��7�hA���v�V~O�A��L8����D�؅eqNI7���<�gi�$�\��b�$�ҴDh	h�s�a�L(Z�M�?������V�����b}���d�J��[���O ��������+��zx�q)����p~�=�������,�{���h���ǈY�v R7`�3ęţ������lW%�eF�Sl� �S�R@����d�E:�k��a��M�̟ ��77r�D0��y�i:? ��?�"Q8�n>��̙����g·*y����Fl~Kz�)_�S�jTK���Q�҉lO�7UJ`7bb�S�=���V#��VTd�U-���nN�G`5i��s����QU�0�:��t�-!���I�E��0���!DE����w��V�M���LkL �PO5��A��>��Y[���,�����9��
H�l�A�_�>��L�nF
�������%�&)@:��kH2F�˻G��!j1nr%�S�0ǀ�os�5W�N�i
F��p~P@��XO4̖�)��@� �K�4b����ZJ�S���F"�)�U����Z���g˟Of�m�o�G��V�n"N;m�4"ks�ΣV|�C�V2oC?�t�����A� �I6I���
��|>�.!���`����q��7�3I�S�{�I�V�Ҟ�#a��$h��օl�CZ���FZ��0��#�~��#r0'���uJ94�6�� =9>#>i0�y�U-D�3��!Rt����k�it�k-����"D���P�w_:XU������M�y�g]q;���#�D�����%0ܚB-)R��h���堂r~��e��%k�v2��U��>����u��|W�=n?�X\�ϻԋ�[B�6�>	q�#4�P�2oS����9cp����X�|ݵ�ܜ�I�e����hC���۽�#S*��}��Ϭ����eb�e9&:*iJw7�&6�Ot?�h����i�T��W���y��#q�LӻPm�p?&n�D�t�u��Ѝ��/���| L��[���C�<�%bO���S*��^p��<�j;����Y��D����������&��q 5Wy������hkxf��E�Ѳ ؂�[���< �x�%6�V	񎜢Z�T�;�F_�v�s�S�ݟ!�c��%O�j
(��RZ �׿v�lB^�������+ۓ���:����ʑ8��@���2B�F���Y���F�E�%�Ҳ�S�o�"V��E�z�S��r�E[M9�\ۿl`20�d�. _n�?�Th
�	|�5[/��nԭ�q(l؁�5!�v*�wh��������2�Y�X��۝��6��5$����վɱ_P������\�S'�n�׬�s8B��[=�V�ɢ��X a������Ӫ�O|�]�q������gv.�PT��U.%c��&�:d�V�&����;�v3/[�r���힧�w��S�q�9���H��$� ��V���������"�b9�%�ˤP*d;GQ��A��bxv�o�k�nT��wm��mX*�����L�<�-��tC��8�����wBϷ|���Ͳ�Q�Q���H��c_)�y9�.����ڈX?rQZ�ݖ�c�#��{� �q+p~,XJ�vi��U�{�i��hO8��T�l+	06�1��}�zL<��Q��\F_=�8a`�]����R!4) .��H�sǷ��'<ʲ~��g{��ȼ�|�`�\ڒ�oQ���w�R6C�l��l��g��+ݥ��Y1c�[p/<Q�X�NzRP4���f~�Oo]!�F�w��Q����j����5��
M0�)`ݔ>F*��+v�X��$w�-�2��Aif0���h ]v�^#��c�m���!M�p8Ň��2�:֑�j��V۷�<m�7�2]�?_��>�`vG���{�4�r�_�8Q૟L`T�@u�=IG�l�L1Z"���3��q"!&�F���)T�h�����*���O��s��L�!Uc�f�*����r顯�Rz��îMP�=K�4y�2_�kѩ�A����>+rMj�}��ՖD�T4��5;-�P��Օ���$sb	�Cgs�9��wE|��˦H��qn0��yb�A����t�������x��ƕ�Nz�'$�z�@@ �Љc�J�&弹t�a�h\Nܭ�-�=�Yw,��z%V��1[�?����c�rd[�����B�(B�,G�7pщ� \c=���z��ܓtN�=�4~�"�p��c��q�?�a���l�S����=d"Dg���IÑA�'|�4,/�´�RC{��$���E�������݇i��I��?��^��}($a�cɈ�ζ��l��}~�ߚ��Q�6�^Ó��Br�S���̑�l~�82cw�q��'n����H��yF�Y�.��PF��-��Z����m���P�>!���)j�$ɋg,2@�)ć�d��j�)w�gv�`���� ���2��ԗ�dfD�*���O��u���s�1c%�d&��P���Y.8�ܚv�xmu1�y��P�����3��G�|Y�t�å�+��x�^��3o}�48�
�W��W.`��,��%@0F��i�3�c��һ�,L�D#��ǐFN�!@Omeٍ�ao�10+��Vg{كZ"v��f��ߜ�ޞ�a�LrhU@Ě�w��bh�-�:KI���dO�	�J8p쪞o9d�)xQ����K � �����7���=e��N/k���-|��d-�Rғ���j��X���NP�N;ё3�U�`
1�&1��$,I_��a� ������۬[��u=8�};H�M"{���:�����7�����uO%�:A,�G��9F��OW$"�#o�|g�[�C�f�r�\���}KnOԮ�Ta�*���M�A�~)�8.����\���旮��Gͥﴶ�
)ԺR)p��nxw��4z��;�ԑ��Զ�9��hȸ�����6KO،�?0��c�
�U3qvl�����Ǩ�:�5����D�?/�jZ=�K�E���m����Я[���7��h͟8bסj�:��|��>��<�;��·�fI���n	�tH�䌑&��R����^s�i:<
V��5���vw�,�>�����Վ�fO�������Y5��C<02 ���L'�����,Y4Ɵ�Ǹ�������J�]����#cZ�g$��(�Js��W8j�V��_a������R�w�$���M��lAd��QI:_��d+����&����9	:
��Yl�Q����������ƶkD'r?�9ФM~ڛ��=����> �n0ƺ�i�ҙ�G;���xW ��I���1Y� �weo(6$�
q�A�h.b� �Q�E��ѲL��I�z�7�[X���|+����/"<(ǀ�H|��z������h-�+�<� ���2�����̱��G%�X��L���b�Ң�R�(y�b4f߆E��.���V������<�=s5���IG�{�Vv|�I.ޅ���o@�)_�҈�/�)��{��� ?c~�z��:��U����xZ�@խT�mF��yo�u�i�ø��U�~8L'�o�&�6V/b9��b����G9G���T����<p�]Z�v/�|4����
a���V�	Up�wT�<�Z��=��I���W���w��2�{	�E NX!�T�ZV_��\p�����qkW{�6=��1�ǭDf� ��q��-!�h�c5�G��"ݽ��V�6�3�/x�1۝��g�2�J���+�z��=��S�n򸎦M����	#�JE������\�n�T���/�������6��=z�(a��q��$2����1/�Iir�6��{xn���_�5�q@d¶QIC䙶�Ҫ�Kf+�L�8�t��:�p�J/��XǇ�&�Kc��$z��˄\{�%"��fIs�X�S�}}"-ꈘ�I~ ��e��|�%�V꼌 ��J���uw�tW<���ϲ y���ĸ�{c7�m_8�-#�(��<h�-hQ�4�q,��U���n�I���m?~�S}ٗfD�uǳ>5�E�r���&*��w��'G���4f��K�H�x]���r.�� #�a��I��V�8���=+�C����m��C3�^4��9�R��/���p��y�r��5�R'M�_m�^��g�p��U�,�3���,^�wˉ��t�Zl�� g��.l+y���Ĭ��7�Al\��FtИ����2�W�?^�/�%A�]�&r%Sݙ�\K���6��%�H�ຒe�|��(X��?��R���bEmܷ,|1)�<�%6���(���MfkS����i�܂�WGc��:��׻�5/ǔ��ƓB��G��P$�ς���G�s��3LsW������Dnh��n!x6`��c�i<�j�&e��m5�ƃ�n�"M�U�6�0-���۩�x{���{2G��E�"e��Uf06�h		vH�P�g�5��1��僓��a_�C��$��]�O#� ���M�v��?"�s������꼭�*�m]�P"L�J/,�m.�7Y�)�bm�҂<O3:����2�~Z�D��~e?a7>��<@�k
�B��ו�қ��D/�#�;����D��3S��Џ�<>��|V�x�ぶ"b$[�����K ֞���9���g���4R�V�n�?V�D�Ip�u=�!��<49��5���l7v�5�N���R~?V3+�&Ū�#����3������d� ]�RNv���d�fO!��|c���/@���q�������;0�+y�~:&|G�xbQ�թ>%��3�w��?g��Cy�
�-��KA�e���S%(T���7���v�sx*7<[�`���e�Sf���3<��
�d���-���n5�o`�m������WwQ�!ͺ�G���?-(�d�0���e��p�c���/���9�t���Spk3O�[�5A4�3�� }Y�;�S���5�� 2�N퇹�}���!�n��#�g����C&]��p%2�@���+����n�j�S�3��"]�Iw��6i����\Z@�X���/̽$���������V�wf(Z�[��b��"�H|T��Z��Ng���fE��o-T��6�"����<�W4)cӵ��|�Y����Oo��xt����� YI��Q
�o�|��!�5>��J�ָ��7�4CI�BՎb�ue��yۼ#�p.$���̻ͻj�}��A�,0����%}p#���� u�߿4&�1�'�<>
�0k��UԵzº��!yB �ط�k���r�������WΉ�����tX��`���tj��nߑ;��C����*�U׃S@�!C)�gmh$/���9lre���,ء��:�v��BUN�>T�⟾�E��,1�$O�*�vB��q��R>Pʽ#[qoP�#o����~'9
��j�@�V��Nޜ�e����N�Jr:���*Sj���*�+�QӌR�e@�*P��7��6>��?@���*�J�W��$���
�L��m��(?�%sDX8Б�i�дu��R�گ XLč��P����3h����_�J7b�1 �^W�b�yj�|�j?����C6$��[�������� � �^"	�K�Xx��mE؋�Gۘ�bj��� ��%�.ƒ�0R�� Z�e�;����}��:\���	�b���U(	�ZGa��5�lI��Q������҇��F�/�'�O��8�����kBj��˘&YE�FL�%;���io7�&�B����S�İҾ*?[Ԩ�\B X�����s fI�?�J7h���	#z�[�5��KF1�#6 l�Μ5(�vׯhY0֍������Y\��"���]:�5+�����R�y��(�W�0�b�x'�Ή��̉s=9I7=OM PnUU��aSf4�%7���/�C�����=w�Y6�v�'��w}Z鋣�.r���ٖ:��í���Hf6vz�.[�����R<��}<�U�qWU��^w�H:�2��P�'~�]iJ���Ј������b�Л�2��*Ɖ�n�H��b_j�o��n�Epw�+O��<*���Q<�3��_�H��;�w�$�|���Ơh��Qu/rq�*/�)~q)����L�!��?@tSQas햎<�#����`�+��8,��T޽��|��p���7�8�\Y��S�+�Jc����}
S*<����FFS8(�]2����z)yK��w�s�ϸ�D�ʙ<��.�l�o��ߥĉ`D�ʒ��L��Y:,C�Y)췾*��߲����1�� pV�_3�z9������§�~p��]�h�F�>�x�����������
�(���m���&Fq"+��[X��w�9��y2A��1O�g����Ȏ�m���+�7���.
b2cvi�/�\#����m��<2D�?&�>T~pGoV��,�T�_���?B����T�b	ud>G�+L������C�B/!-���m�TI�D�va�汶��Tao�(�1!Tp!\O�f�h�Ar����ٜ����ݮ����-{)�;��u�L��;��B%���*�M��1A0�՝^8;�L��	-�@�\[�U�GbP,C??�@�L�^�㧍����'����0�ub0�Q�?��t���T��4ݠ彯�����`��7@G���j|1J�fi����a�>�Nc8�-3��e4w9}ɉ��$εh�[˥�ڜ3ncs�
d��l(h3�-ʘ(I6xG���p�te�dc�l��SbZ�,�lt)}=���~�G�p��̕wl\�!�a�.*ʳ2F��=��_ye�km�QJx`�o�w�{#�/��{�Y�{��8$�Z!EMU"�\i����磏�GZ����$(�G�/�;���}��0�~�f����b�Q�6��$�Z�B���|�*���~+�c�����>ۯ�����y�0G˵�XPr�i.k܁�F������w������j�i���q�2�֌P0�k\j��w�2=v�\Y[ ^U�27x�� �CD�����,�����i&�j����ї��GY5��n�?��14�]p��?Gd�zU�G�a6Y.��p�+Z����3���4�n�枹��~J����6���@�D���@3�T� 0�sV�DJ�s�H�Nr��@�$~e�;���d1iu�ʷ�{ k)E��MG��cW��Ei�<Gbh����bzP��#X�4�"K0���th��ӳ���Y�a�9���xx����HՂ�����􉙨���f�en��Nv�\�"]���x��ݓ�ab���ߧȜ� �N���3ϻ�`\9��ڨN-I4���+� ���>���H�u��d����ͬ��:���O�~v)� �`uV~�:(��G���FZ�kOި�Њ!R���g�f�Je&���h\�g[}��O[�T�rd�.��hM)����e\� 3����mH��˶�z �38)w*jn_֧���hz.��9�<BP�� ���x��ްQ���뇱���*yn�m�5Uz��+S������h�$�5IS�ˉ|���j���K�ck��P�r�e�"���y���P8ɶtj	7�9E|��%A7����^i��T�(Y�3�Ǝ�R�}ev�fj���܄;#�#	�n�S�MC�j6蔕�юP�����@B{�P�D�փC��p6\���H�IgZ����]1Q{��\�K=Հ欔��]o��=�q�
�е_Y�"��-�\�X�'�M�J]�"i��/�{.u�S7V�����~��~OZJ�u�[���IDJ�\eu�7;+�<��扨
��4bT�~ҸcD�3��w���V�QR������x�s�gV؝^�>�b�;~�����k��`���{�B
���&q�-l�u,��A2kp���=,�����Ŕ�EA�)ڷl|��K0�/��kk>�)���L&=׿�!�=
���i8sҀ ó}m+EM��
�zOv ���}M�C���Q�7��E�-Ƀ��d,?<�M!�
��$Q7�q�G+�e
�V	#���,I+J�q�FL�e�J�Tn|�Ǖ��Ő>�ޡ�٣J�͔Ӈ��d��b2k,w�n�.A�@�7�?V:�H��Xf��%�.����ύ;ྰ��%Jr��T�n�j:�_������r#X�킱~�W��{$bN�:��q�F&�Lv�류?����S�+��ˌW�8٤���fa�"���?�9��&ɉCT�*��SO��a\��;�33Ү����;1��<;vk�<�� 3����*HXW�C_B;ھ��$���L�E�q�VZ	�H��am����3�E9�r�������hڽ�6�Ԛ����a�+qp�鞢��ߓ�K��S(��mp��i�,���͖�A薘�VH!�ay �}8�G�c�JOՎ�^Em�gV;����ɸ�Տo�Ұ'����J�ݤ���V�$h;�eh��·3��߲jQ�kɣ�Y"(S�e�c����}J��|Eް-l���NBR�+jh
��K���})�BȨ�O,�PN��W�+2���
��oG�'�B�i�d���<e�W�|\�]��:w�vb�1��6�W&doh�	_����e�Հ����F��'1΄Fv�{�ł����\d8T��RR.����нU�����Cɹ��Mi��,�]�����/��&���$=�0��vm[	��>r.-�S�/a�⢲�B\���
���=H�"&@]?�r�e��B�F� #}���\:v���E��-�
���[9P�ڙ,�Z�����q㺥^�=#=�� &���	���SW��ɞ�ka����>'s�C�t^�&F݄�8+k�W��ހ>j�!��s.d���FQ�ZM@�ͿM����Ċ�\�����@�}q�ƨ�����]�M v�-��+�O�ܹ'ԡ˨;9H���z?.��kZ�O�4|�;U��'��,�9XyR�%��N: ��\d�4g<�ץ��.���mAÎ]���<I��Fl�n�P�R�k{�6���﨎�e�s�w7��쿂���Ɓ�����K`~�-�(�ѿ��J����Fs�����zy����B%4 #���Bz�����PC��?#��Va���B�ZR���T��An���a8����ڔ�*�U�B x5i�
H*��Q���A<4N. ������Hr"WJyi��Ǯ~�;��ں��CVD�t#�|���XgV�'}��P]�H��?pCA���l��a�+T�m�S�^f VPK�Eu����"
A�����#�����J�Q#���b�/����xH멪p���d���[D#��_%NP^�+�S��S�I��V�X��Ѥ�ؒ!��m;v�6���u��^����уG���[,"ڟ-�Y���qI�^���C�#�pĭ��ܸ�5Y���r�T0����q�w��%�[Ƹ�ոꟿ�D��J<i�+e��0��@��xH�J���WqlDV�G_���v�lɢw�S�$|�D�f�Ylz�k����_��d�'^��F����9,\�+	�lĥVU�#�RLa�� �o4�'K{9�
~��R��s��`�SX��s/G��z%�@�����p <Z^���1J����>e(C�$�|��:6�.{ZU � ,EA����k��Ez_��[1�:�u���6M��h?��;����uH:z�����쿌a��+�o�Y�&�vz	�n@d�J�� ;@Xio��ςAb�9zԋ��y	�f���E���.�Y������~���Un�sn_��!I{<|C|�`�.��R���@�ӎ_$߈�˙)'��{%{ ����3"��U�屖����y���3��[y|G�R#Ñ�U�"Q�q'�]i&;�
/ۙ>�#2��G��I��T�<�H]��S/8��4A~��lb���%	3�ʐ�<Ú��-P{�E|��eِ�V,���	��N(��ۍ�}Z������t�N�*�V{�K(�������i�ڒ~�KY�%�h�7k5�N������>��Or��h3w��U�(���N�J�H,+b�����������֙��J�,�p�ȍJ�Sr��0�\|p!�mTŤhF�_r�q5)��@H��{(:�[q�ܫ2��/�jeUI�o�6g��/V�qL�_�7Dq9���j%�C���+�"K�<WL�5G�-bY��~i�/��XROc���K�ݳФ�'����\T��%�fba�X��}����|!I��Ʋ�w���`%���Ճ���$g�3����ʀ�~'���B��ı��cP��;W-|G��S~��Q��J���Κ�w�������q�}r��f�Yǌ�L�>?���.�*��X���Q�f�X!K��DxV*���I��9�^aT%;��F�83�,����Z��l���gC����咫ORKD������R�}�ˣeR@z_��'^�њg3����9���b,W�ˢ��t7Tr�8�g4��l��������ZAe����(t	�d;y���I�z�����/��A��n�?�7�(��tB�h��΄L5�!:�೤����(�(Gɘ�4��1�Km�Ą,U1��5��6�%�(�W�M�����7c����icsv����ɺ�������������P��ׂ�W�瓤�l]:3e���F�M��Ͻ��zd-!1�`�4�b�j���� ����nk-_M?��6d����Ʃ����g&{k���@j`���C��H�6�����OH��g�%�X��1M�,��������ה�:>]��۞9;\���[��".��X�2�D_�6P]�m�"e}�/eP�.q1�7҅z����ꋳrO����鷛��*DƵ`eq�7���<�$3�$�]�����XҴXyDh�Ϭ�03��=�o��E�!^]�s;�B���ŧ�����M�>p��)�^�\15M��qU�G�>����M�#Z }�Q�beG'�7
��Y�%�?�$����ދ|�14I�GUR�J'�:�,~��y��̸�L�����4���Dh$�;�w�S����������!�F�����R>K|�C��ܡ^_���vs�ED��%����m��h��"�.ی�6`+�-�W�*_�ר�� x�譧	ȕz��ٻ�(Brr#�̵ZH{z��܇��8��ȕ[17eB2�3�}��T�<��3�س��΋#��|���q��Μ ew�iD�*�/K�R��A��h.-`C9:%����W7��i;U*��Ym;}�޺�9+C�hD���ɽ�� �{'�̦P*�V�V�/CN�X��f���T�X�?^�(9P��u%R��/��A�7�P����%x�~��>
������O�x������v郼�>�[q�$ع�%�Q��8 ��ZdEI��E�0�1|�N_�:�k�}$ܖ��&u� x^�?N����r.ģL]"G��fj���^cC�M�p�+-�tH��-Y�٫L'0x9	�َ��>>��4���'k����ݱogJI����)K6�-�*5J���W>��Voa�_���#�����w�T�$	�Ó��lG�����_"e�dqf���Z���9��n�X�Gl�n)�_� ��F�ƼE�'8Z;9V�~ �����s�n ��=4��R������B 	Ǔ�!�F?�euNk$��J��H.��p �
�E��-�����k�z��[�M�4�c���5�F�S|��-�H�*@z$�p߶����8b+&+�&�����9�{K����M=�XV���\Lvb�4H�XFzyvn�f�c�E4�Q.�X]�����V�F,s;={��X{IF|[�.��
m�`@k7_9ُ��&a)�W�{2�� �D̀��� @yUMfw�ڌl�F�)��U̮�y�\d���~��Upq�~�8'��&��j/�U���o/���HG�]]�CDϓ(�-<v�] ؽ/ES�4�'�]����Q	�jbʽ�<����x��R��ѽ��N���	1�zNU��Z��Z5����2�!8��w�-{mܨx�2������+�������h3��5�5'��Ƀ�B-��|2A�5���|�5B �K]~J- +O*.�M����tQ�l�9�O4�JK5x��;w\	�$���5�5����+��~��T	��CZ�('w�qG�!2(Z�7��I/F6t2�aU��'#_�|�qƃ˶�Y4C겅�K��LX�`�z:������%/�XX�J�즣K��C�Qͻ���\A/�%�=af�O�X���}C(��WAIR�������=%�(�O$��Ut���t��;�=ײ���Ԑ�>�qc}Se�:-�r��'G�+�Q��R�7F#�d3b����O��3wv��}��fJ#�y�o�ˏ�J梫���*�g��e~�����f�2K�Ynx�����l���a��T��8���C�g�	؍}7�����d}����CRX�z��B�Y�?���X�<Rms�_s�^E�5g,9�蛻t2�7x�$,�����}t��uM�gAs�lq8���l}���A��9�t����DG��M��E��/�rAAE��lJ�Y����]nO@� �� a�xy�@�n��|�(^;��n��Y��ӑmv�,BW�º6p�(���M,9ݺ�J���͗c`����1K�G��ǚΧ�Yv��g�Pj�q���瀹m���3����|��q[���@��'�!~�a`������j�|G�͌b����nxM�^�6�b>���&D���%�{8���g䃨�G��U@6%�v��>HB�g=X�%�@1��Y��M6��I&b���]xg��f� �S�B��ލ";��z�������[k]#Q"��D/2K�.ޅ�7�g+������L�O�Df�~
���.D�-he�<v7�Oi<N���qu���
]@��gLD5������Y�r���<�����|,:Vx�_Ab�$��q��S��<y��6��K=��'���\F��nB����p+X,=��}�ףŝ��9��r,�� ��8���'�R�G!3�R�0�ЊLMޗ9n�Ҙ��`�p Wb�RT$L���dt��gQ<����ͺ�9�-@���w��%20ٴ�y:vY:l���_�Q���>�x�yb��4g�/�yA�	�s�5KGX�ʖ5�S�2T�@|�/�#�1L7�EH`'s�S잝�y�I�/Kd��&-3��n{�`G}�Q���4�Q�Ѻ�kܛa9r-����v�x���X�6O�R\+�uC��?)�:��ٛ�ky�� 5���,�O�Y�s���ᇆ��f�VT�X��h�lA2�gC�n�������v9&V�ݳv�\2�9e�T��ν=n�� S�#7���L����Xiw�u�}M^@8Z ���̃���8���-ʥ����=��ZWr����"��~B�d���-Z��g�A|fIzo�����"����w4�r7����|�b���oPEtaL	���� ʰ�IE�:
�U�|��!~��������(־�7|7�I�F����0�?ѽ#nN$j��#��0��裇��P�0��<����#m��fzBu��W4�t���8>P�0q�@U�wJ�@�_!��Ǌ�k�k�D���MY�j{��Ӯ�O&�ׄ�XD�f;��:�����;�P���&���	���G8�)�g!h�/ırS r�3�2k�.v?'�U���>Z|���d��1l�jO7�%c�<�I��IS����>V�#!>(P�(�o11��])9�m]��6��A$��5"e�?��*�P���f>M*�1��E9��1�T�R��e���*�¨7�;�6��?ƍK�p��򡈥W��N�\��P��L���m��#?3P�D��N��M��z��P�����L������P�n��⴦ec'�,�C�^�n�1�j�:S����Я�IfՋ��z�C��KyP �5�$F��сxtE�a�r���٣�s' �gA%��f�c��;4�Z���;�}y��Ԓ��a��\�(U�w��(O�gZM����I�lϯC#~/��h�՘ݪ��2�d^k�UQ�8{P���=B�������Y��F�RM%��m���o�0w��Ĉ�?��S�Ŗ҄L�[Ze\������Q�A �v8?�(�h�i8	�N[#�9���h�)�Il���5�(�vW�:h_}��O����v�Y�]�(ף#��5�vA�کh�D�R;��{��@��h��'��#�dl\se�_O�/=,�`����aY>��1v隕�ڥmI�M�o>��2_Kv�y��=E��.R�\��:�q��3��Ďu�v��+[�˗�9dW�п�� ��qA����H��s勰���7��	�9FЎ�4�kG�bF[��x��*���4�#����b�x@o��n��Aw*�W�[�[*� ��||�<j2��T��N����wO�]|A���0���Q�juL��0R�)D�%Ē�-a�'�Z?k�Q�B����#ý��J�+}�,o���Ɔ�B�W���;�H8��:����+�\��R�}՗<�K���F���8.�]����_A_)�A��ߟ;s���\���߮+�4�g�5���+Y`����Ù��ʤߡ�C:����^t�8w!�W�H1�L&p�e����z:S�摈��~��6],Z�F�ł�>��,������b6
�vx�6t]��WFw��+c�X$�yw$-��̧A�ɩ��{�O��kf����m����N���=����#�2���u�]�b/�ۤxYmY�2��,?,��>�G��P�(8v�Z�h_��w�Z1�̇�T���u*�6G�tAL�ch�;�ܚ!����TO���<��7{�Ś�>�.���j!���f) ��K7rV���_�?�A�8��O~��@����_1����ZS���5���KM��B��#B���T��-a���D���LbV�C����.�����,��n��~'+07t�b6r��t��t���4|�f/�[����['���@jn���J�lT���aa�N��9-y���G<w��͉���TH[��bI�c���dx.����R�(��nG��p���O��cJa���0�2t��	=�~# p�{Ǖ=N�L<_a2��ʹ&��:�=�/�;k�35и���/Lʁ��/�����(�{A�$�g�E���s�;C�i��ƨ���Ų>�}$.�g���Q�
xV��M�~�,�߇(I񜰙6>!��`o�B�/V�R��>�D~1NcdqАLĤ�D"����y���;��P�@��G��~G��5�������0�j%h}�8A�2��~�X��֛j)w�}�vg�;� �
$2=�З���D~)�#ό�߇�/8�>�>��ѝ"��JeY���	=��EUy1�Z����������G�L�Y�S��$o+`�����3|I@4��Q�	��D���9*��E�@�'%ᇄ�3��N�F}�yL�D�-TعN�?�@ۭ�eF���n�}1�7���S�{�*���*ғ���i���(���O`h�r�h���~�B���]Kv��z=>�I�W��W`Z9��lx>�t�HJނC���oٙn������e��N|_^��2���  ��(�(!�e"���fN��k3�p�`��0鰻�T�I���n� E���DƄ�Hc�u��ն����o\�r��:(����M�����#�u��:npYG��MF xOd�O�ОJ��g�M �$г8�J\� s}���O���T֐�4�q�.Y)F�����\��Sզ��G�R<��������)�5�n�R}����z�W�|��qv��p�U�k�d��c��,������鈳"U�M*����N6�]I�u�5���Q4_쒻j�KwH��yΣ����(x���Q��u�`8�~j}���|U��kU<�	)��$�J��˼4�#	(HaH�! ��y�R2�+%�i�'|V�B�5au%�G�	���R��֧��c�w��0LLk���lxf3�����90�t3ON�xS����'ka�I�)z�+��|	��EtC����x�a����
륽i�7��:Tųw8xE���
s��0���h�4R��0�Ҋ��7�C�J�j��>,���M3ZD
�$˯Eq����_�q��gz����, ��k]*�A1<��-8���n����>އ˽�IJݓ���5���J��Ek&5�O η�����U�9vӂ�sX��%G��a�	�U�!X�x����^r����諅:>O�C���r��
��-~��[��΢�:v�џ@g�L�up� ��X*k�M�؇���S��^���T�a�/"�G�J�m9�&e�}����O��xaM�æ�V:3�\K���,;kԜ<��?�uc�6�� m%"s��H�G�=�G;zf��.��s�L��:jV�عHxj m�&�m�9������������6�7��s��ѹC�I�pj����D�	<����nS�(��'c�
%Q�f=��GG�A�V��P�0ɛ'��_��h�D�{�4��m,�FV�h������Oǣ���������t���a�V�l;���h������䰙�UQ�����(�0���p���^}�cA��0v���g�� YBWC?����
��#��}O'YBBnvO�\
N��W��h��
�[%oA,��ڴ���dgA]�6�W ��\.*@�U��p5�1�	Q�џzd)�	Y�4��$�������9p��1Q�v�&��Ƃ������ ��f���;���q�W� ׹�����`�k�x]9�O�ָ�i֩&� �ǈ�=�������	,%=r��S�j��=���=���E��e^�\E@�M2r����׏���P#�?��e���d�IvqĄ��ySrP�2�f�[Z�����qݖ�^��=9�r&����Hᙍ�5�C�k�m��t�s9�tض�& 	�S8em�Wr�M����!�&sh�%�y����:��M�22��瀀Pɥ��z�'q"�ګ!q�	��MZ���m�O�� &'e���c�ڃQ�?�O����n�46n(Uߑ>'�D<,K>�y.+��tj���k4�G��ѝ�h~4��:�CT����װF�$��
�R˽a�p�o�n�k�c-s�6��B8�������L����۹>.`�r�-`�����W��)���T�ռ�� z�m�و� B�/#����z��������/��ٖB�p����CT;9��5Ü����[���1���`��< r\Ki��*�7�?�TA6H�.ZuL�P��EWD�i�8���c;j8��CJ��DuIo�6��3���'�"TP�����C{{8��G@�kT��r�'�^�{JPo�u��k�\i�A_i
���-����%���Xv���؅x�MI�*}��f�@��[�2Ű�%H&��ef��'��I��m�R ���0ђ���'T �
6#��Pu���^^տ�}ѽ�^{X'�9��"�)`���;��9�^z�C�~pM��a�p���]Y��#��I�0E�$�F�����ͅ_ ]�2i����>8�JvfD��	G�d��:TӅ�RiJ�W+��V�f�_�lI��a&�w�Xr$�����ml4*䍤�q_O��d>���f�D�OP9<j0��Fl~Z3O���>ݒ�v�)�('E�G9Xn~m�1y�.� �uMS����-�ޫ鍰�zq��;u �Bq����NI�Юe��N$���tB�.��� �#E;�-���\y�zˎ[+�p�g����R�"7p�����3aH���z��-��⌛��+sT��	�p��Ǩ��~�>Xcꅡ	]b [M�E6$y\�f��E1�.ew'�����U"��ies(����g{v}:|(��.Q%z,�@�7_�����P�)!��{_ Rð��S����U����'��3fխ��z��y�XD���Ë�_U���'�e&5�}/i����ls�G>���%��u��<c��]���/rCV4��}���p	G���
/<}�I�'�r����Cy��w�}	�IN�e�G��Z������'O��_{z�K�%���@��ޑ����\�h V�5i<.���k���=n�"na����b�?�G�JpP�+\�������U�j�a+���k�fG�1J�u��ĉ�\��N��ӡ�"w��Y�	��:l�!��鰷/(4��q��2e*i�$�I��6�-�.�3�+��_�D�qsMq��X�Cכ��%��KvaL%��������k���/kشX&�y��KҰ�('�TR�\Nq�%U��f�H�X�۫}Ш�;��I孲C�@���^%H�h�OE���p�-���'�Ҁ
m0�s�i퐒��Ԫc�F{RF�-vm�T���Z/QT���D�r�Π�/��<
L���Ş2�A}�'�f�Khǆz�x������l3*����ȴ�s�f[d;K�L�x�p�s�����aN�3�3��8�� �5�����*�L�^k��QNk�u�R�MB����K�Ld��R�Wb_`us^��WgY�,�h���B���[,�����'t����{gn�l>�ӹg&��ǳA��jht�{�5Q^4���98β�/�5�A�j���%�FQ�n@�|t��`\�>��ي��"��U�(KGɒ#3à�
m{��,O*��o��6QE�(�fM��ۺ>s|��:�cmɥ�2n�����Ǉ���<��2�P7�"�:M��Q.����3߲	� 5��1������d�!�)�`�;:���WjI[ܺ����n��=M��g6�.��E"�����D�Hó�8�����.�����yh�ԭ5a�.��w��>E��x���|hɂZ���>�Jh&d+TP���F�Mm�Y=��*�^�X
qJ�ý���n\�����o�F�Q���"
��F�}�(,Mq��2]�N��SI�P�6���&��#�_�Aqk�2��s�C�]��uKN Lm�߇������#W/ck�X���q]K� ,�w��L��\F^�%MMaf�S�XzE)}�QJ�3�Z<.}�$�ܳTW���(�����!kY"����s���tV�,&>
��8#�W�Nk�6S�!�s&k��,��R��M}Y�	�=�T&��E�8)�q�$������M�Y%1�#|T��Y'̘j�3���l�? b�c��G��4t�%U�c�'�V�,ɇhyJ�?��d�2+��T�z40�ύ��&n��e^�U�����Av�Fd�k�H.�R����.k���-Ǝ�b�s��� ��z)��쉭���w�G`v�=-��������Bs��{8e��7��'zq����"B!P#��\��Mzc����0��Ə�]�8	Bݿ[���T�O�#5����Yx����ɔ���Ms� p�!i�.*��}�A4�.������@ǆWBhi���v�.;��к�\C��D��tX���&Nm�'u��PU�����tC9[=�d�Y2�T�Q�x�g^^�fPC�nu��;�'wA��Ѫ��㋸Uhマ�I]g��,��~tx@a��h ��je����[<�j��%F`�#�O��ADI����P	\ќY���&e�/���yutu�x^�An�
�>�{�D�6Σw<["ҟ8�Q�"�i'�^��C�_}p��4U���Y�5�j]k0�g�������+I��Dư���p��<��J4X��#3�Խ��8��p�NJ��%Wi��V�6�_�<m�n)d��w���$te�^^~lrP ���2_��d��b��Å��9���#�l��XMm�J������g)�'C�9��A~�Gl�k������KP���k�n��:�8�Q���� 4����F\���e (C$� �29�.s�C ���E9]���*i�VzWXe[)��m<\�.'ܿ`3'��s����H1�z��d��`��Y��+�^�Qc4�n*��f��B9P��Xa[D���b�lԃ�yf�E�.����OšvĚ�M��sf�'���{4�|�޳.�*[xٸ@�.�_�U����)��{�+ ж��+�3�q U����,��q8U�����>Oy ��JP É�2U���I7M'�F�&3�x/Ӡm�*⪒�G
E���ғ�v�<�{�]�Lf/0Y[49ܾ���`����	n�ʈ��<�s��%H*�=s9�]�ݖN�i�H�	��N �ۅ:�Z�_���zV�l1.�"�{x���8Ǿ}���[u�3)�{h~��5��:�����D�Gt��`tC�]�� 4�ᖌ�J�E�+ZX�����ӎ����3��W�$}\�~�J�ȯ��D�\t��eF�`9��W�T�i���n!��h(2[8q��2�:_�brI�7�6_U��ՙ�i��_�;	q1$\�b�C��#19K�{5L�S��%?���#a�Y/�$XJ���wNHK��}М�(���\L�X%TCfZ3�X��}�*�����I�����+��E�%p����)��)�+?���JS��Ų�����ĩ#�cHmk�<�-t+���v��Q��BL���������z^����>���}j�f���Ǆ���6��6̫*ֲ�P��I�cf�K��xN�헃s"�1
GaL�0���q8+��4���C�诎��	m���9劫iRCCe���Ũ��J��^R8��_�A�^�I�g����I�����;,Od˚�[t/%�� (g,�@l��L��?���A]G��t�3�K�-��������/��A����7<���ؒl�k:�`���|ɀ�V��?���	�(�axɐ��XV�)�m��,M���-�u6ϗ0(�oM�H����h�xV@ck�S��F���������ϸ:P�x<�(��d`�3]A9�>�7��W2ϵΨ�r�!)w�`�0��Zm"j�ux�������ncd�M7�"6\�Q��:���
?�ɹ{c��8/������6�*h��eHyC�g�f�P�1E�ǃ������K}����]��1}�~�~�SGJ"&XY�P1�ꛁ���]���"]7�/]I.iI�7ʜ��U�h3O֘��y��.'D�&�ei[P7�?�<��g� �d��ZҬ�D`�O�kB�DLK�E�*�7�U�\�T�V�Nw�N'bu���\N<��vΞ��ȃ
Yڰ��������0]�i���pv��=�����?�|Z(��_`�9��4��,R/ʒ3�l�ś���TV�d��]~<�Kp� ���R�!?��d��Y2�����E�t��:�/2����0�B�y���:7��75�Q09�>�������gƘ�y�(l�>��Kr)��!,�S��YTC��Ei�[�d��7M��`/�}�JCS�!��Ĺԥ�2d��-��!nF�a`-ǅ�0���r�QM���2л�l3>-0�Ax+�ۦ`��V�=U,��Y����E���DFkD/~>5�\j�e�6�YSΜ�$m���7�1�p=�d��W�%���Qn>�Y���%�&!?R��I`2>R߻?���%�nj?�S��Ѐ�租��FUFi[�h2p@��nG�̎И�����y��,0-�Ȓ�ZB��.�"�3XMg�&sZ�C�g��f�r�o����N��"F�^��.4K��Ƃ�|�S�N��o;[Zt����;( Ղ�I�,
�ִ|6!{!	���l���U�i:�7��I�읎s�SAO����#Y�,$`s��}VD�;���~R�0�M�vn�#j�1���`uB�:4����T>��0��U%h��+��!
�>����k����cM%��V��Zx��q��o��XM������E��_>;��u�k�{+���Dܒ��)J�Zh�#!���rvA��]�p�0�v*ZU�s�>��3#����5Q�P�8��ɋ�7ߌ��>+�#,�IPMo�ie����9[%��G�P��ݭ�V�Ϻ�e�:T����{d���PS*�����l�ܒ��]K�e1.�*aQS7⣃6��m?�����`�L�W�4������L�Pm�[?*�D�ʚ�mN�Ѕ�y{'���s[L�b����;������"VI^hwl�ϊ�j3�h��V�<��\.��X�y��t� -0��<��x^�UE�����Sb�	� ˶6%.��N���6Z���;��e�nhQ�K�v�c���y�b�(�`�Z�����l:���I"��A�#���C���%� 4�8��ʁ���B{2��3�Y�~F�I%�UE�5�o�C��9i�
��S� f��[E��\Ӻ�X���\t W&P?���h��	t�5[#!���=��C�lВ>5�v"��h��7���%����Y�C����.?5����|��7JH�����|�8'�3���[s0;Kzǈ=�����3a�ܠ����1u���#t�����\�������vw���HE��|e�.rH��:\4.�����0v+Y\[��߈�u����E�K��q�^c�Ϫ�H�aH������N�����й������b1�;��_.*w~�?��9i)bp�No���nL��w!�����*�,���[<����c��y���2%w:��|����w�lך}Q�@��[V})�~ ��x5<��
�?��QR{F��B#�/�+h8�,P���ncu�M.�a&�_8�-�L��+���)��}��<�X5���FW�8Y�]�6��J-e)
����2ls����o�ʪ���_������ `�_����[��aΤJ�`Cd���
�����#ٟ�Z�1[��p'UչP VzJ�"�瞑;t~���]wpF��H�IZj��������-C\
E}Z�!L��6-�F"K+neX���w�ڠ*�Aa+Ó�T�?��Ve\���^m	���M�h�0��?2���ź���ۯ�&m�O"2U�d?Wv�>�$G��|�s^#���_ȁ0Ὣ���T�t�u�j�G}81L)�P��p+��Z!������TzN���z��"����M�ٕ��!M��f������r�I�J�W��GX�E�����,�C�*V9�A:��֊��*�6�.Mb��`Վ�7L�6�6-�]���A���OObsC0�1���o,姾�P����i�0�<mb�C@�At��*�j�����å�F���?�rI�@L�[��J��l��*8a��5N���-��%��w
]��ru��ƀ�[��4��Bc�7kdS���2X���V(:q�G�l�p�/bڅ�c5����|�ݾ�t�n�=�t7~�a.p�&��N�7N�a}�p�d?d����=������2�g���ۘ �T�,Q/��u�Js�{�:$��fE�pN��G��?i������T�Ĳ	$M$Yɀ�������~�րߒ��qP6	�VË��Bj����O�̉��~�rlco+󐷿��l�@�y>�^�&WeP�����R����}�� ���6��S�j܀Ƀ228�.!-�\H�j��^w���v��|j� �l2�k��E`D�*/��N��S����)�ʄ\��H3��pUY&����p�E1��������
��+�LG�M�Yv۞��B+�R[�Vx;3g��403��O��Ow������P@(���n�3�������$΋Dg{�p�N��@]e�
��Y��1���{Pu{Ѽ'�J�^�ߔ� ޖǒ���hMS�4���{�%��KA����AGD|�BD0�)19\�xI�"���U�g���H��Y���Be��N'�������$g�D��s��ǐ�P��F˄N3�I3�nw`i+�]�:�IW翛YI� �����)�S<�u�"�uꈨE���� :�ș�R^/������uGMH:9SJG��ZF��,OO����5�Ig�� ;���\�W�}C�VO̊WTYAA�ߒ/�9×)�Pf��8\�|�L��;͝���<A�+q)h�np�����z*�����r���ߛ`����1�.R�G�����ܯ��̣U+�����ݹ��F����5�֢<�^7j�jR�QK����ed���S�߮/5H�`%8Z��j�L��
A�|��:6u�4B��ַ�߼ȹ	���H��N���R��S�V9�i2��V��5���nywo���z�r�c)���@�ks~ léJYY��|0��O�3x~��0kL��܇g�֩|�iE�w���_xg~���C
֡~i���������0\E�
>�[�%$�O����_�5݃7����%��ذt,$��M��/|%$_�q6h?�jC������]�,.����ɾ,^��*�s��#�������h�>�����fJh��Ӭ��)0�}�|k1�
���#�sq�%ƺ����mW�X+�G%�䜠��t����Gࣺc#l�r��3�_:��.��o�rrh��ҡ�~��m����   �   ލp�F˸�$�R=�1�#l����O�ToڬrN�'|W�DC�O���]�e�����:Vؽ�Da�w5,Qlڿ�M�F�ilZ���T/f�l����!��TI\&�L	���I!����һi7&�����o�x��f��T8���,O���bM�HR��V��x�Il���>yUJ^2_�Y�C�b|ެTf!m�04Jܴ�M���F}�*�K�	_�ts�\`�D97K�p��T��B�	5?��0�)Ҿ����6`�C�I�m�̵9��]�c�B�L���C䉹|�z���#CR����_8D��C����$h��ѻZ�\�)�Y E�C�I0<ĆDY�*]0�|9�)ˀm�2B�	�V� 4C�l��,ŌD3��!��B�IY �z�ꊘT�\h!���1ݰB�ɯ>�h$3�Ꚋ7��H��ZLB�I���I(�JX�t����`���C�ɖI��D`�YU��=��@ax���>	$EJ�AF�s��ʻN���QD����O4��V�d�27M>}b�ǚ�ug�O�� �J�-D�.ez�,/2�\�@��d��O��L�\�4ᐛ,5�șv薹���AC�>Q�1�S�#<Q4��-}���"��990m�g�<QP�I 2  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   5    މ04�̐��%�R(O5f��p��'l����I�l���   ��@ӌC�A+,ɘ�I'\	~�`%Ϲ>   �   ލp�F˸�$�B��>�1�#l����
�޴Y�:��O��d�����	�����"fŰu�pph��^�wS,�ش>G�6$}�8����
x��ј�R&?&����[���x`&�j�"<�C~�����Y,~(��v��e��W���%���36ڱ�-)?aQ�E��7Xp}BJ�8���D�5{>���N�!��X�Ӻi]�V�Ϟ������ē��.�-!�ph���Ȯ.��x�ȓ�V@".V�>��`���G@�ȓ]d|z�	�i.j�i$e��N9�ȓQ��
��p�GCO�kk�����ZG�<��"��(VX��N½,�V=�eH�<! ��/q��̂0�� n��iI@�<�P��i��`���?��%b���P�<��*�=E�2�:C�"�D@�0b�M�<���c�P�Cc٧o58L�1%Np�<I�"ϧ3��m��->n�a!��o�<���f���'$«h#�+WfD��h�'��Ň �¸��O�=y\������I"Qf�n�󦹤O��7����rX$��N�1^n��6bD�_��➀��I0��B �3b�F�d���
q�9�'t�Ex�}�'�R�j���2������6�|���'�L�k@ ��<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&�   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ����Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �'F>�БY�D¥p�N������?��O�`M ��4u&�̧O4���k���W�ID�4��B��0<�bH�Q���[1!-}҆K!7�[�"'@l a#e��0<���ʟ��	�����l��}Ҁ8@�؁���XѮ1�'T�����F�xu�����"��'H4�����(0tnРl=��B��L�m`���%�O˓3v�h�����y9��Z��]͆�7oMeM8�'�- N��A�{��I�2"Ȕ"C��X�b��{E�ɩ�4�b�����uH�%V`��K"�
j.����	��@&?��|27��� 氹�G5S��Sӈa�I񟔇�I&I��0��Q�V@*M�gc[� ���?�4�Ӭ L;�EFO�"�J��ڙ(����\�`⟜�S̟���q~b �1f�^`Ke�4Ac�c�&�(�yR��5I&���D�R<5��
��
��y�H��V.�bĨ�'> ��Υ�y���%|G^X�5,M� k ��S;�y2k�d૥߾����	���DIA���X���.X��@�T�}t�b�:]����O.�D�OP�O�'T����j*!tةĄ _=�/Oi<�q̌2s^��S��]F<ձ��Ԥ/Z:\���s_��R2��s�ƕ�5��	���w$ៈ�Iܟ\��Iyʟ1O�8�d�3hjq;�LH�&�*��.D���f�Ƙ0�b����%H�d|K$�'�Eڦ���OyBLz?�ɟ.�8�Ό�}���O�b�^Ě��'��'��<�B���)� h����n-��ðiO:��f�'JX�J��dт8#d�p�S�
�b�M��M�ax򠋄�?I�yrLV�7�|U`�!�9�� ��.�y�V9*8=0�#	,3� �H�����?�2�'PL1 b������h�N�MX���ҫl�����AC���j

G:Ÿ��[6R�u�������	0a��$ڣϒ/*0,lBE�¾l.�B�ITQVm)�D�w��ѐ&�~NC��-+�����(��[��s�+˿0K�C�I	\̀�'�.Y�XMH#$M�?��?��퓨)c�A� �Z�P���O�!!��ċqO��S�� ��z~�i�"�V�9b�A�]��L{����yBI�*.D�� #S��+�^�y"�� �k�ፇ6:���y��M	���D�%/��0�R��y2�Eyֲ��Ќ�25�p�%����L��(��)cL�*b�*E���"H`�3V�TsDK���\�)�3&.�p�_��PU�HݮB�Ɂ2�����e�*Y�@����O��C��sy�T棔(H���q�ːl.FC�IZީ1�f�,�[��ȯ(0C䉺I�
Ĩ��H? ̑�%J$!���O2lE~��M��~BaW�J��8B��Ũo8�TH����?)L>A�����I�SH ����g�4Ȏ�2��B�	� s�9�S��+29�������.�B�	5AF�XR&�4*�ب��P�R�B��eN�uR/�P���N�G(@��������� �5�ج��Ŏ�m��t��J"ړv���D�d 7$^ ���(ƨFf�	`��2�y��'�a~���|Hh!B��6$;����y��A|l9�e�c�N4�1i��yҮ���#B��.φ)cѡX��y"�R�hF�y �ޙ����w��+��O\�G�d��̾��`&��[2�M 7���?�7g�����'�����p$��
��3�S(=G�	��#D���ԡE��9�ER�\�]�`$D�p��I��R����WK	�}{S�6D�h����+>�8�C҃H(5��A��7D�d3 ��5)JD����m����@�<��)ʧ �Nq���]�^�qD�7UJ��'������'���|�����8e��h97\��4��BA��ybcN1n�Y��D&����܈�yr�O8
"�P Ɩ�A�E ��*�y�$Kd�8(rA�@�U޽+cNε�y2��h!u±�(
�Iq���W���Xá�����U���J�j�AR �?<2P���g�O*�OR�d �3}�+�����h7HךnО0�#���y�n�
�����n�hi��Ŋ�yB�]7i���)�m[�2�c��y"���bH�H�mL1{�����?���'>���R�I6(Ӏ�:�`W*e�8=i��DR0�?U��-˪�lD��QYP�ן\�	{���pD�	l����0*�:2���q`�(D�H��.��xh1�I̝e�v�&�3D��s�״X��9��H_8HKf2D�t��c�[���3�o�+�.�'�+�j��>�P@ȓL$L��G�B��h���O~�2��i>��	ݟ��'cH]��N]4Ռ���D
@ifU9	�'���l�5rg�=k��5��;�'C� �c��
7Q��ٰg�0�2��	�'B@1b+��C6��C�J��&!X�J
�'6H��J�.��)rr�N��T,�)O�Dz��mV�)��oӴFX��b�^)Q%� 2,�d�����$��>y1�*��X��N�MzS�!D�� L�
Uh�9w|1f�ƯU�8�e"O�Q
�#�sd���F��
Pk�"Opա� �t,�D���L�n��k�"O��3!L�:H�nt�@b�U6�S�|��,�U�t�="r��b�ւT͂|�$�˚S��9��l�ڟ���O�C#�G2:�T��%�,'Y��Qq"O� *��@ЀKD)KV��yB�P�=�����⅍ 6<�îK)�y��V�B�"e*UFԬ|teP�(C���?W�'�Q3�H	*rD���)+� i0��$�+?��u��T���0���+��9	�
�����K���r-��,�Y���u�Dq��6D������&U���/ �I�4D��I��-�"y�H\%T
 �Y��0D��@r�J�-�IYA�;q�9P�j0��U��>���D��N�Z0-A�Ќh)�O�)��i>��IڟX�'n��G�O��Iu� 41|���'���뗂�9gAJ�
pGX�!� �	�'�J5�d`�;g��!�G$I=^�jH��'Vؙ�����pBK�]�8
�'�@xbA�Ɯ{JT4�gd�WJ� �-O�Fz��)����y�m���<K5��	���	N��y��ԟ�&��>�����t�R���)�&,1Pb3D����:r�s����Q>��m-D�4A��2HvajC��%|(:e�(D��XGH�4\f�ɢ��:r<8aG$D���1�+��e�0�W/r�t�q!#�d�r�'��(C�'�25jca�dՔ�j1CۓY�Fea�����?a��L��҂��GF��`κ4�6�#D��H�η�X 1��ا� <�4D�P���{�d����/X��]`s 3D��1n�3ey�h2�!ƾAۼ!Yt?�O��	�:P����ǀ l cF�Fȣ=��O�k�O�ݐFL�nr����ؾ!(Y�'�"�'5j\z��AR򎁺�`Ȣe�'��ݱc̜�R|�w�:�`��j.$��B���P�AbЎҴV�tm�ȓ,'��۷i��p����$�˭EZb�D�� �'C���T�œZ�n��m�?���I7?��#<�'�?)���dч:��Z���&�Ԉ"��ܫ.!���d��Ư�_�v(�X�(!�
M¨�CLH<+3JA.Aq�!��	1E��@kE!3�x���,^.@R!򄔨g����`��<�3���l_��=�HOQ>9����2{��q�D���ȡJ'	�<�1n̆�?!���S�'SG~��$��:\�'�� ?�
���)������ʚxa��d%B2N�Ʉȓ ���`f��{��MQqoJ2\q�a��9/�qQ�*jN(����� ��ȓ4���+#h^6yR��Ka+�;���'����$B1��$�0l(e�H�e��D��<"�|��'���s��9��;ޠm��ǚ�]��@$"O~$��?c���b��ۮj�D��e"O���TcL��:�0d�Ue�����"Ot�� �N�����EG>�x�9��'��D+L��!p%/8R��z��z�ў�h1�,�iqn�`I�L������MX�<���?I�/��8��b���i��]	%���ȓ|'�Mk2΄���`��Q<Eh�ц�Ԙ���'j���x���%�L��ȓ#z<��Lט&.|؃�E�J���F'-�'<m��Ӆ;.y:�8�b�9o���	�N�"<ͧ�?A����ѓ�m3H�,x��Gnǉf!��<l���s���rWG�q�Xx���� �z�f�5 2Ր���,�(a�"O@c��`p�)&��#A�+`"O����퀰s�P\�"�)M��Q�[������ӻtU\9�	�r�V}�0S� ʓXG4lP��?�H>�}Z���mH)�7�C���%B2E�c�<��K��@:@A7f�(4�	B7k�E�<	��<F]� �,¨���Rj�Y�<���|��h1�fJ"XB�8�'��V�<9�R,[&�1�t�@qz��P�ɦ��O�����O���V�<~{F�tH�	P�jY3�'�'���>��;���ӡ��7\�'�u�<�I�>$��C�ω1l<y��)
t�<i@YK؈��= `ei%�q�<��(�9W��a���U�ґ�5�JH��x;�:eِ�1.��]ra�C!� MD{�n�&���nc�Ԇ�d%#%�)!�F(���O��D4�O\�
����;�*� S.�&tx�"O޵Jf�3|
�z'R&��E9"Ovy)�gą�.E���1d]�R"O���p�@�D3^��b ����5�	��h�zȄ�Ft����攐7�����'������4�V�D�O������i�+�\�N��l��a�ȓ"��j	R(�V.͑r��ȓY��1�(�";��u��6@�n��]zT9���d2��񦄵=����1�
��g��?ޢ�����'�6X�'� #=E��'[�p����Z�s�@(3u"��������O�Oq�,LS�꙽w�lZ��(4g���7"O^���h=X��a�)�"&/��S"OR����B�l<hd���\
U"O�9 ��P=�!y��ܵP��D�r"O�0�� �[����)�O�P�|�6�	����D�>�a��:d����ϒ�&:���^����@��O� 
��YN�"��Qa��M�H�	�"O�X�B�E�[-�rb  �ޥ@"O�d�e��\����͌t�&�!"O8ĪG�ĲoC���a2�@,���'�����a� H�3r^e�bᑦA�ў\F�8�u,:�H��Lp���F�,^~�(���?I�v�)˖��?H���	G<?�ȓAX�I��E 1̽xШ�N�r�ȓ_��rGݳ_�m�A�ػLp�B�I�P0��W�S׼�R*G(EjƢ?9�퓥R�<�5mєpf�`�j�l�~�D�%,���L��p~.F*�R=Ҥ����퉖����y�&��i߲���H�s�����y�BY�����\�m^P�ˠ �yr��/W���aFیi�ZIa�eP��y���>0��Ö:8;���.����$�p��(��y�AI�2��XKg�� �ΜHR�d�������IL�)��0R~`a�~�)s��ݼ)�B�ɂJ�2�Ks�֋�hU�@���C�I�l�yc%�L;=�2�+�B�$Pd�C�ɽCd04I�f@!T8�4�\�kbC�I"P�>9q8�U*�,�(�Z�O6�E~�k���~Z��d�*�5!UaO.O@�����?���L�(�a
�|�,I�vi��ǐ{�!�ĚS`��*J�t�t��IT*a!�DN�k���fㅃi��GH�[�!�N"�­p���$V�xS2Ǉ������O>����I�|�yq���'al��e�I>p��#~B����kjƙ�`��}'�"R΋�?���0?�6�-^KL����$�va�U��x�<yM�1qF����!c�h@#%a�p�<� &}��̓1b���te^-+��c"O����DybP��7�R/R ��ڳ���h�=H�C��S���B�J���'�
����4�$�d�O��P�8i�C���g���P�;(�����ƪ�:$�G�$7>�	e�7q ���Q��q���%U�����ƶy:�`��3��\ぢ�R*�q�f�1\�J���:�$<Y���*̦���-�5u�@��'T�#=E��JS.������6#V
�?���1P���O�Oq�lC���	1N4��TO�$
�a�R"O�u��*t�"%�a'I2q�n�f"ORl�C�M�2t��(PGZ9/؊M�"O�����S��<���3hd�hc"O��2�P )��bV�;�	�1�|2�)�
y���:��J7��+W�|��g��x�ҵ��m�ϟ4��OԀ+�X>|��l�a߄j�z��"O�zզ�>=� �K���!��Ċ�"OP��kԼec��4Du��iE"O�����͉�T���蒉�H�x�'�`�D\�,\f��SCćm�T����K>
�ў<��4�.��L)�ҍ_	d�@	G��>�i���?y�l�r�K n��u�T�����@��N����s�4��m�4�Iٮ$�ȓ+����X'`�a35m҄-m���~i���pgN�8�#��AQ��F��<ڧ��'%2��ڤ��z���0�#<ͧ�?y���d@�|��٠;D�i�W?6�!�䑺Rx�9�&�B�1�,+R�!�D�9qF(�\
2)[
�^S����'�x���L�DSX�rIцO���`	�'0��`S,Ǖ'T5�FGΔD��I�(O�aGz���M�9w��Z5���(��MC>f��6}��>���i}��>�u��$O�F�!Ǜ�H���0�B�?���?1��d�����(+���O�O۪��T�P�_�(E�iг/�J]i��d��h�����l���3��|*S� Bx�Y��dǙY8�-�6Ƒ|�'b����?���F��dʹI˜)0̾\�����D5�O���WN,����C�r\Y��'���A�@>_&Z���V�-�&D�'��ِ�'l��9O��6D@�0 �׵\|z�ȗ�O�,)n�$�����Eڕlq6��$��"~T�ʒ��y�+��i���	���<93.Q
P�4�%ɐ0Rz�:��i������OV�\�jlp��΁8��M����'X�)�)-?	�A:+�X��¢i�|*q�Jk�<��,D9�"lr�զ+<,�Q�c�'p�"�c�0)��<1G�;q�dCB#F9B�d�P���OKb�'��'Jp��-�-3%BU�umń#ߨR4"O��(R�<-��	59�ʧ"O�iC_gx5�#*íN	��ڷ"O8��a�
�����Q��"O���,Ű"$E�.� RH�P"�'7�#=E���"CE$䃲�U�38�X��T� �����W�2�'ɧ(��T���_+!����_��P3�"O�����mD�}e�������"O��g�I"'c�`�6+������"O���˘w1T��5iw
�$��"O�ͱ�(�Q�:�� 4Zd�U�P����DܿK�f����/S:d�ȠelA�A��X$���I����ɣe�C�(-P&��O���C�	�.����'�� .�#��B�ɻu����!,Wإ* J�>m��B�I�l��%z0�F,G'�՛���)O���Vy�v��D@�`��A�'H���'�h��4����� v�f��4�N������$-��#������e�)Zh\hW�(D��01h	L ������*6X�p�+D�� b� �D��J�����E���v"O�����,�����`F0�HK퉳��T���Q�V�t/�0{��}��Z��O|���OD��<��	�Fw�-�b��yk�e�\�B�ɨ
w�-�!DHP����V'ZX�dB�I#_T��'GS"7�	�3&��J�(B��1p�0�D��P�B-�fh�x9B䉂:6�x�7Eߌf1fe:�o҇L���dTx�����c��ڣL���3�hԡ4Ib���OP�1s�O��$3�哄J�J�X�f�B�`�C�I&W:H
0EL/`F,u�� �>?�C�I B!Xݚk�/#1L� � t�C䉨!i�CP��2�A$��N�RB��!e��x�B�J	3Gb���ƙ�,ʓUڑ�8�tD2}���r��3$&�:��Z�3���?Y��0<b�g��@��_�;Y�@b3ms�<�Q B�]jv��¤1�J�R��Hp�<y�f%o��Y��̗X��e\x�ȓ]����E�]�XR���لy�����	;��ހ(9�$!`N�#YE��ޙe��	���	~�)��R�@�ys�\���a�O;LO���禅&I"���Wg!+n�`v<��즡$���	V6���KW��<.-���B闇 ��I��~�ɗ���|�j��%#W�}�#p#X��E0�kY����FT���h��~�O����!�4mwJ �p�]-@l޹�W�g�do?���9Oh�1Q��h�vB�$,������J�JA�#P�%�Or�O;b��P��"�蠠Fs��3�R�ݦO�|�g��BҶ ��C������^�p�E�ɓZ9��'���'l@�zM�0�ٴx���v(?1d|�c$ ��'�А	J��k��锂[��Ucp�*���hL��X��-?P�O�s���??Y$�B�<��\�U�ǍqR�����Y^(��+O�}!@������l�ȥ��IB7jp�h
�<�H���9�~�KV���?�	�Ayb�	�]�(��d�ZiPy�0��mh�$�İ?��̸��꓌�>��;�#�[�<9��Jc��˔�n3�(��3B�IlD�����e18yq�b�nR2C�	�W��L�s'�]&Ҍ�P��7`C�	�>><��L/)����&ÓFaXC�	�y
(<�#擶8<��@�@�:C�I/��DI�T$����F.&
C�I"i2��O�w��d�τ��B�	F�,�@b��8_p$��ܳD��B�IZ�R�C�C�Q�PbP�h��B�I7,��r"��'����C��.q,B䉜L���QD�{�D�JP�՟0^"B�I�
82��U�W!Б�ňR�B�ɿQ1���-Dif����7�#<���\"}�*��]�̌��HǀBy�U2���:����F�2�TMs��L���0ɲ��*apX�����1=~�DY"I��0]�� ����� �C�/�\��1��0%Șt'͞�m�VY��-��3CL�{�ĉ:��0��l��S��6�@�+�5X޸�ʃlϳ*uj���,�����h�5 b|b�6(�����=7��)�r��"<�T� @��� �R)�`n�/s�����
P )萮��1*&H�p��1T��s�_�p$yb��!cdm��@�8�(Q1b	�u�̃CA�(gtly"K>��+�%-F a���g��P$�@H�<Aw`��N8��@�8.�>h�E��~�<iBL(�>��s ��`W∢Rd�w�<�㬀a�ƈ8���0Qz����r�<�T�׎.��2��ȁ^�,$b��p�<9�a�',�)��_��f-JVg�v�<�'��3PE��)qO��X��uz'OJv�<��	��d��R�X-%Ǻ����HH�<�b�Ǽ��%�ë�n�"��\�<��F�N��v%�uq�}���l�<)m��R|����"KX� :��j�<yb�P|�1c"��$H�jM��N�Q�<�@fS�mg��p���7i��-�M�<� ���C���xU�P�b@ {g�HU"O^���^->Uq�;guP�"O8Y�E"L�LhPoO_g�,k�"O8R�%��/r�R���~�4��"Ol`�J�5?�(C�됛 F�R�"Oh��L]�p�ք��1�i"O(��0I�jU%�U�ՑE�hH�"Oz��O��n8�ae�Xw�� 8t"O�1�j>)�d�h$�::�\�#v"O(�6OGN��1�)�4(Ph�"O&�Z�Ӡ3��1{ ���2T��"O ��` �	Ј:D�<(����"O�Rխ�9�p0�'�r��8w"O�XQդ��P�x��g�\=u� �"O�$b"�՗Z9\�� #׮��y*A"O6�٣c÷qK��Xu��+_uv)��"O�SQ��9��Հt�2"OX��L$BM��lhO|�c�"Oȕ�`��-��	 ���d`�1#a"O2��%�N#?��[�l��R��(2t"O ���o�9ql �{@��{� ���"Od���)���@�k���i�<|�4"O^�0$y�y j��~�`�"!�yr��`lŊ��A�����	��y���"\_��{a%�V�ٓ/��yB'��`n���a��R<i)��R��y�!|�b(�v��+u��2�@��ybbN�`:Ը�LW�g��Aķ�y�ˬ-h���=a��a��?�y�&ۜ-β�e`��O�: �׃��ybo�i�~ �4aؑK��)1�/��y�BJ�9⺼����B���%��8�y�1*��c�6�����-�y� �uU��m:֨����7�y���(�l t�4����)�#�yb ���,�J�.�0a�'b@?�y")��~��]�?���V����y�+��R�b���A�=A�Ԋ����yr��w����&�K�t.�+�y�oH�,��R钀v�"%����y��to~��%��gθ(CmN��y��N�5��9P����i�Eϝ�y��_)��-yŋ��J��Ò��y�A�4L�#�ܝ�� ��y�F|�u� ��t�T0R,ۊ�y'� ���)n�%r�9q톦�y2 �:6�up�/lc HBa&�$�y2)�.Vv@�F��-~�Z����y�B�(~�xCT��xy����#8�yB�=�"m�w�*_՜ȋa� �y2�Y�gO�\Y�j�Y�J�@H���ya�>{ؽ���'�A)0��y��7�j�q�kO�J?�`t�
��y�B���@ D��:20ś mM��y��!����f��+:`�I�gG�y�&��,�bE�w��05t�;�]��yR(U*�D�eO:u�1��#�y�k�3(������'J9:���y�E!ɪ�`U{���CO��y�!���̚��	t�|@��M��y"-ϻ"����b��X�>�顈���y�OW�^���P�o�:GR�Hi4F��yB���>�ʤ��,�4B�h��"��yB���� xF%6�B	�Ʀ���y
� ���v�Ę�B$�ԥ)�f�@�"OVi8 ��6pR�K�>2���i"O�I���F�,�l8�c�:|�p@R"O�8� i�.x��i�X�b�
�"O���2W���W�M�(@X�P"O6	z�
9\��ZP��$K:�}
�"O�m"��Ȼe���"�)d{�Ԃ�"OjWnڞ �#0�ҵudvHs�"O��A��֘;
ȡO�zD0Q��"O����!W�\;�MS!D2���"Op�l0"���1��O M�~ �"O� ��2H9���89�ԐSf"O��)b�W��0X�Bk�7,�
�s�"O|P3����������O�R���"Oru��*�zP�<�
�&tEJ5�"OPd1�N�w�J�ǋD���u"OP0�D6E��!Rċ!i�f"O<��'�ر{�Ђڰ
�mK5"O\L�B�J�sp��VK��t�hm"O�� ��!{z��SJ[�v1�	b3"O.��SJٰ䥸�nĂ(:�"O��ࣦ(H�V<x��V�xU"Oj 0��λkچ�ɦl�6;� 4�"O氉 �Al����4kN�S_�a"O�M�V�Ҟs��T��W8YAK "O$L�o҂x�6��〙I�1ڄ"O��ѕHh��0���ķh�N5��"O�U��a�"D����ˉ$_��P�"O�`�	ܴ=�ʳ�L#\��]�3"OT��F�+�)��l�*�"O��6+Kw���0�٬�x���"O>��q�.�p�+5��?�~ݛv"O`q�`W<<�l���>`�ZX:�"O`a(��=y����D#&����"O8|�ׯ� I���ڠ�V�?���8�"O�T�P_��"���0k���v"O����[L���1f��a�"O����+��M��895�y6Ʃ`�"O�J4h��n��AP�c�`'�Q"O�q
��֯Rv�|�g���"O���� ۳v�,,{�Y�R�8�"O�Ö�����8T$*����"O�\�d��L��l1�d�>Vh�]k7"O��@K�<k��a$D�-EVD��"Oؠ; �?��,Ţ��+D�j "O���F��X}4�H��<v%��c0"OLl�ueS9F���RkA�D0�;�"O��aF���LU�L���<^��p"O��0��W�?$4���+Ѣ=�BP��"O�D�s/9$Z���%��q�ݛ0"O2H[�b? �j�;�&�Lmh#�"O��"g�Lˆ #�CO.\N�;F"O��)�d�*J�tAT�ZgF���"OJ�I��C�6�Pxه��}8
��g"OTZP��)h&��o̱)�4ằ"OuX��/Ww��(� ��>�P�Ib"Ox����,.pP`�� Ա"O�-�G��+��"��[�ԕhW"O�\�����~�8=J�J�(0�Tѣ"O��K%��z�zD���N(���"O�L�p�)!0VA�Dh��-4"Ox=�Q�N����RG?ZK�Ч"O�qhVI\�R*J�buE��$Ap�ڡ"O(A�`������S��`�`"O� �Y{&aO�F��(��ԩF���A'"O`��TD�1qfxY{'��Z�1�%"O�T�e9J�vi�g5<��=��"O��"A���S`d�bd`�XWB�#%"O`Q�N�I+���hF�1��峓"O�Xx�+��q�@<��GZ�J�,�"O����-�J�65��� "|x4(�"O�< M	;9�̙��Q j:0�2"O��p ��\�����)/��@�"OFij��� %|!���X"�Db"O� ��J�^)JP�e��+�h@%"O>�4�SP�ᚷ���I�p%S�"O�q�WDQ9K�p�DeQ29 ���R"O �jDB�-ɳ���7����f"O��+�2�0	��V$	��0��"Ox|ZҤ�R��"�a�#�l�۰"O~�Ј��@Hk���7�D���"Oȵ��܇o� q��/�_���I�"O&��D���!�|AC�8��u�"O��p�ѫ.~��2�N�%{v�;�"O:�3 �)!𨫲��0z]�"Ot5SHF'jޠA�D�l�ж"O0 g�m�n�0T"�8r��ur"O�Q����V�Y�$k�:a�tL�"O�iS�ڈ&� hr2�H�V�B��p"Of$�LP�"�v}dL�
{���"O�&n��e��(�G�Y�	µ"O�D����;|Nq��&��Sq"OҘВB��/��u��F�<|y�"O`��s���/·>��7"O4D���5J�x�0�`��_���v"O�c��� ��S m�}�@Q��"O�����QHhJ�#�e�.�� c"Ob�CeA�!�2��F��F�: ��"O&�)�"�r\0�[�d���Щ�"O�p�3��?<d,��D
!F��x�"O��N�,��lp��R%s!�\p�"Of�:Q ˙;-Z�7�_%�cb"O:܂S�ɷ]�w ^�$D�X!"O�,�C	��>�� �IL��P��"OD���L�Q&��0F� S$"O��ӄF(&�uȦ�����z`"O��q�'fU�#����� �"O~��g�\���ӂ7��;�"O4��¹��)r�! }h��G"O�I���G�r���h^��"O��)H��5c7/�S&�A��"OV���A!*\��6�MzyP��p"O�E�s�Ϊ3͜�*��ݕsr�y��"O������0$���R�=({.�P"O�`�q�֝u�Y�2G��Dz�(�"O�����u��"aM�w��}��"O|���m+1���)uZ��ei"O<D��aϋ�a���G�Xq�G"O���k�N22ǈ��+�"Ot��3ʐ2&�䐣���"`����t"O6�xѭ�0K�.IS�/E�)�hp"����zt��͛N5YvM�^i�'�����[l��E�B�N)�'��g�*ZV^���\&|�X`8�'�ܝ�ơ/t
=�c�߮!����'��`�3�e@L��"n�i�X�'B���t��=W���#aoG�
G��	�'��M!�"ПLN��0�>L`����'�����	o_�{�.ԏE���p	��� �T�4搥!��Q��='z!�P"OR������kH����>3|f�pR"O�]���S�.�>���"Άdl w"OBx+���U��dK�2PT#"O`)B���UM<u��ȓ�1J��ɕ"O `�/��y`����|��"OL�������bv
�m�dt �"O�M�A���"�pJ�&	���"O��SEFN'�Ը��c�a�:�P�"O(�2e/՝
�,�r�kP��b$"O�4�S"Ӂgd�ٙ���unt�"O�u���E=Y��o1p�-�"OjPX�h�-\��]��i�@O -�'"O~���*E�W�di��/X�6D�a1&"O��h5�ؐ?�zՎ��\�r�� "Oq0���"p<� �������Id"O��+0,��i.��Z"E ���@R0"O,����!7�\<��AB�u���""O��(�KÙ[�fQ�R.\33���"O~�z4�?S���c�+�$lj8�U"OV1�à��x\!%�#1��A�"O6��_&s#B�u��6�"OZUJ�`J��tAk�F@�Mp]��'sj,��b�,Xb�yjg,ߖt^�Y��'��X�����Z���
�LB�~;r� �'���a�lҨSq^��q$ÈHiLPa�'�)Z�hP����4���.!@��'�����њhQP�2����'�t�)D�Hj�%�s��7*c.l)�'.TtS!̢ɺ J%
\q�'A��s��A%B�ATj�.��a:�'̩C��t���┫�� ]�,�	�'`��ǂæ5�����W�.P4�I�'��Lծ�;�9!I�)[(@�'���!���FgB�|�j�'f��+/̥VjX3�#�9�P���'�<��C�_�x���gĴB�L�'�8�@T/:�D���.�K�Py�'4Π# BѠ��Q�C��-0=��'&��1����oI�%�Ȑv]��'za�	�ZfB�����|��'���B�"DL�9ϗ�M.$;�'w���Ứy��С挒q��r�'�ZMyƃ�O���a`XY��T�
�'
�	�q�Q6�bq@�Z�[:���'A�e���<����3���pX��'���F�D����2(�*=-h��'����" R'N���B�7�l��'���CM�8���+A*�%
�'5��AC �/\uh�#Wo����'G���N�>jװ�4��k���S�'�\� �ZC��-�h����'�b]ص��z��k��ϓc�f��'��)!�dG25�=R���4\Z�'����RH�4l'($A��S�"��:�'�`�A�'ϻ}(��4!��LBI1	�'i�*�W.;�:%#�G
.H�r��'��a���	!d�Pr Ʉ�ډ��'��u��&�)a���ʆC�kf���'l���G	[�=���ڑk�2�n(��'N:�y�	"���B%s'&�k�'��	�2م	�P��p�^��X
�'&pyO� �"]�!��H�����'T~<�Ύ�/{"-t�U{��(���� tlu�L3q{b�#Q�@b�2"O���Ưv}4YB�k��
M�)�"O�� ��	4�>�EhM�y@�m[�'XV4XtE�2c�;�EC�_�fIy�'�� �鍲K+\�@�]�
<��'*I#�T���V(2M�2)�
�'Z�b �?�8f�V�Kj\j
�'�:mH&�M�xy���߼RP�u��'B���W��j1lLm�E�'QșQ皈R�vY 1d��.��ap�'~&i��,��ԑSuF��-��J�'���!]);��Q�']

�	�'}Ԑ�����@�`�aԋP�a����'ȡ��N��%�GmZ'`����'yؼk@H
�1�`-Br��8�{	�'E�ٸ���"�M[%��.ZJ��	�'�"`�Q�[	j+�� ���"AH�!�	�'� �HB�)<y�@�W�7A�Dlj
�'�jq�kY9$�(���̗v�$�' l�rO�&-|����A�;h��s�'�Aȷ��7utB�!!�ܞ,�$�@�'���C��^�~�H�bJ�$SF���'���i��_Z��� ��*/�v]+�'~����A6� h{ B�p��)��'ڪ��]6�"�X�ϋ3@��'��[P�T�s�	sǊ]�4t{�'2H1s��A��qҫ�*Sg��	�'Iܩ��_N�xy�'@HE���
�'ۜ�;d�y�\49 B�0}��
�'�9� f[i��M0e_;dxP,3	�'2����	F�8��B,U��|	�'42 ��TÚ�SE�Ɣ
d� �'w�P'%Ƀs��|�g��9�eB�'�
��
�I3@<�I-��a��'��Œ�JQ��`C�1[�L�[�'�xa�5��t�D���^?%G��y
�'��b5K\�5������#l�$��'{��9��'�z�+ �Ȅ:5�e9�'�����h	I!~9p#$�03�%��'��\�����}۲ˇC�_���'�܍��h�{場�WLėPǶq��'#:l��u*oޫ2�XE�	�'T����o׌$��'R�*���X	�'ǆ�Y�KȳXdlU(�`ɺ%�����'���0&b<h��ㄜ�"�ݛ�'x������?d�R��e�H�@���']��bǁ��E���Zb�����	�'��2���z�0�T�P�W�Ż	�'HT�A���*WH�t��R�I�~���' ̬���K1LĞIITf��}M4���'s<�rk��a��Y�ǥ�@�4A�'�@P�N_+F��F�7A����'|XA�\%9�|�Q�ͳu{z���'5<H"�	C�!I2� oSԬ8�'�H��擆-8ƴ{�΀�l��%��'������م���nD�`�~�:�'�u��'�E��mRR���l�'Ih,�Rj��S�)��D9}G��'k�īSl�(b:�)���:�8)��'��4��Ԁ#8�1�b��N��1�'��K�84 �E`�$ۮN����"Ol�q�čGv0��ʆ� � Qc$"Of�!H���	p�䅟Y�
�!0"Or}�7!�Hg�c���2��}A�"O� b�[P�
8x���ʡ!�+X�^� &"O�%�!���xl�S+˶D3��5"O��$�3f�䪰��Q$:�p�"On-b�L�"�*P����q6H\P�"O���e!��az@�Ŏ/"�H�F"O��Q�E�8���2��ز9��"O���F� /%C����ސO��zf"O2�J�.@��J�1�Q�l�B�"O4� ǋ3Y׺����Q#t���"O���Qʎ�(��� '��~~�8D"O��:3 X�%˸��P₄u4���"O�pR�Ɠ(p�����>6i���"O(��`��&a�J�St�Ҙ#�Nxx$"O��b�G�	Y��Y#I
4�V�Q"OFi��/$m�#Q�&�B�z�"O8�80i5G������Z���"OJ���'Y�5vRp�2��;w�x��"O�e�w��s4ʩh���7j`�y�"Odh���O�XheC%��f�Rq"O���N�V��ʂ"C�J8�8�"O��0J¦H���T) ��(;c"Od����[?&��Dt�-,�����"O��YSG�3�@ڕ��!8Q^�r�"OR\�"j�!Ǻ	F�Y�p�pm�d"Ol�CF��>�ĉ�a��4^nB2"OV�@��A=Uq�iu'K)x��d"O^�h�2��hs�fL4_A���"O���4�V�Sp�T�EE�pm��"O޵�W�H�>���ۀA�]���"O�`XfG�=�
�Co_�Y��(1�"O~��U��6_  �,��~V�"O��s!��'��<Yc�M�Q �"O؈(M�=��Pea�<+�!��"ObH@u��$V�xѩ��&uDp��"OT�B��	N�|��N�O~�	�"O��外�S�֙6�SPK�Ѓ"O4�x��;y�&�B�d��5���"Or
��"^�H,��E�.~��`�"O~�5��6d�Ѐ��[�ʥk"O�d�Qa��S��yP��'���Q�"O(��Ė!!!Rͻ�A�s�:�r@"O�p�@J�l�*Y��/�
����"O�q�����A��&&��e��"O��7M�,�p���E�p�D0��"O,�%&
�4�Xd� �U�.�&�j1"O�E�Ŭ��S��� G_E�~�YR"O��Q.�%�n�8"�Q�o�Ƽ��"O� �eڇr�~���� =��C�"O����ޫ'����"O:v:&�Q�"O���UH��WB��tD�)H$�4�"O��H�W�@��K�/D�=p5"O�����L 2aI
��<�|m��"O��y@��s��!`�(e���3�"O>(2H�)��L��B4O�Ҭh�"OҌ���B�PI9!,=Hoef"O�0W䛀H�F�Pp@�ZZ���3"O�m;���+[�B�s�kU�T����"O"�� ��ԘZ�*��L�ٗ"OtɁ�mM�rM(%* ol,Ȉ�"O �������@Fׯ	���;%"Ox(�0���"�4];@���;��������o�l���G�!�4x���"��'�LmS�դ�05BA+I��ح�
�'�j����W�Z���BG����'��x)�"��;'P�1���?'�h��� �jŹlΰ��!�I;@W��v"O�m�d̙!<NAp��:Fv)��"ONp��.�!7���9E!ج�0�e"Opp����r���4��s"��P�"O����i��\!���TH�+r�]k�"O��	B�*ph!G�}�u�"O⩛���w��8��]	�ĸ"O��[�BX��Ph�$�m�0��3"Ot�V�C�(P]�Bc�c���1r"O�����[���Q"��dxڈ"d"O�$sыIg��`��=
d��B�"O\Q$��2D� i ��.pZ�R�"O^U�"K�u��P�� BX�`"OZ��wR�6�Ƀ'#B&AZf"O^�ك�b�b@�#!
�'+0��"Oʌ�b��8�$��> ���"O�]�@�#/(P0�:8�0Q�R"O������*��|���X�9:�"O���/�� �V�1C"O4�)��n�[�`EmS��xQ"O�:� ��j�<<���#�嚅"O%Ň�89EM\�r���@�"Oq�bZ./[�HA��R�XA��"O��yH'W�|2F�^,�Yڶ"O$A��/3��4�7㑦j��""O�Ջ�N,l��G��u0i�U"O��҂�6NX�gAC-M$<�!"O�u+#Q8$��p�Q*ZN���"O��)��ň�!�GW �iS"O&�jvf�'EXx��L�s$T5��"O�X�!��е����;x)�A3�"O@���'hE�t:��7J#�IH�"Ot���N�IQD��$��m
�$�1"O*t�5�	7|z�Ű�����$"O|���D͍B�b0�ւZ,<�M�q"O&ũ�؇m�|�$@�Ht��"O����cx#P!H��� t%{q"O�P�է�)V1�C"0����"O
�!�O:A5N�L��A ��d�<�ERZo��e��)@(<�`�b�<����2ѦA�gȁ;N/�d�E�F^�<����-Y0�����EH�öM`�<Iw�Yw� �
1��Z����d�[�<ّ�Z�j���&0�b7i~�<ID6
����DEɤ
��q㦝z�<yE;/�T�i�$��}Ԩ�I�E�]�<q%kL&Jcց�Y�L����[D�<�"
�4"X�Yb�Oӄ����c�u�<��=tļZe��>p�I�[X�<A̫Yx�5���/k�M��*V�<�O�0"��]�&��eHAi7!�T�<���� 4�ݠE̡N��5��F�<�ShE�n_�
%�6
|�{d�k�<qюD��D����\�F�:�'�d�<1 ����9�X4�bС���k�'Q?
�)I(=�`ЪL�
aPz���=D����Ȳ�|9�4
�6+�9�$�;D�PK��<�"|s¤ƴ$�x�@d�?D�@r�gP�qUr4$�`������;D�	�f��`�)�(J���15F;D�h h�W>p�+S+O���y4�:D���)��
m�&�ÀYU�|��h;D�̘�oC>��ӕ�^���h��&D��y�.L�w��S,-��1Ҭ&D�� @�CGΒ>���T�G-i��"O$͂���z5���H9�"O�9��U1GS<|��`�7i��q�"O� ���Ha��K֏��}	�4k%"O����:3�H����"����p"O��"R>C���x#�!Dʎ���"O� A4iɱ��=�u#�f���H�"OLt���M"dy�A��hP!�h%!�"Ob`�w�@&�$ �5��5Z8����"O��c�/�.�bH;�/�!S�`bP"O�q*��,q�`Ccn�LCPI�"OQ�U'�,#��(�!��G��v"OT��TdŲM���r0��B��[�"O$)�3���q��,y�@��pC��u"O��`�#|b��/��N�Xp"OT�j&/G)5��a$NT�$h�j�"OD�� nȥYT���r�Y�k!�t�"ONe�+�#)<�1� .<�8��"O֨���Jш�����T怢4"Ov���$މ?���[�$O�,m��"O���t�fj�4�a�J8�hd"�"O�K�^�o
�ͫ��HUu���"O:�b$�ƥXC	ԅ s|�+�"O�	���Ul�)��G�MpL0�"O���B�2�b%���Ū]T�ّ"O��Ê�h��zeʑ�qW�Ū'"O��+'�F�t?�p��k��I�Z�;f"O�`����f�(�k�'ОZ7����"O~$H�-ÒFN��fD2Y;t��"O�*bgZ�#eb�S���s�:��"O0equ	Ku��(��P�,�� �"O"�����(�Eт	[��"O� '/\���90tA[9$yʔ�V"O�3��%[�� C@�g`���"OE���C-h�183*;_�1��"O�Lj�n�:��x�5�e?�U�""O��Ȳ�K�yL�
I��5ȸy�"O�)x'Fɛ`R\�h���V5����"O�X�1�N�\���B��G>�	�B"O� �r!ؤ���nt�"O��Q��F��y��

VP�!�"O��YbO]�|,��;�G�]8��Zp"O��pB/rC*c@�j�||��"O�YeIY0C��lx����$<�c�"O��0��KU��U��)1�\+"OmY�^᠔��хh��1�"O�.-�>��ӯ�OP:u"����Py"�ց-�j����
E�b�Q��KZ�<I�-s}�}�D�]��p���V�<�6CQ�;l�У��+~6�0�jYi�<i�g]�K{F�X���[��-Z�<� L= �lQcs#��:���ѵlXQ�<�0(#b8�X��aX $ìzr�_T�<�A,�K���Ҡ]�) �Y6j�P�<��F��Px�y!M�Y`��N�M�<Y�͆M��$��U���+��1D���s�F��ˢ�Ӭj�ȘR�a5D��� ުw� 񂄍Тi���kw�6D�:�g�vhLŘe���fc� ��9D���Ɔ��~�C�'s�Uː���yr�%�:T�T �&S,B�@�W�yr���V]ա3�,_� )�Ŏ�y�U1�6��f�*{����G�7�y�*�dxi��9ykv���M �y
� �}�r�32L~)�+��+9֩s�"O�X�eaC�*S������-J.t�!W"O8iXt]�R�2�R�)�����ac"O�0��DP����"o_L���"O�Q�F�/J�f)S'�4Lvh�if"O�y���D��|���T#qj�أ"Oh� &��jU�:A�� Ag�x��"O���E��}�# �2G�*�B�"O�+V�$ ����3��d�`"O���I|"p�5M$1�*d(T"OV���� )��1��)�*��"O�I ����.�2 +S�V��Yx4"O.|S!�E+b���1ʋq�t�*5"O6�k�ُ,�F@�R/D�&����"O|ԙSlO�oB9aڅ8�ZP)�"O�JTIU�@�����`F�p-�y�3"O����ھ�\���aC�(/0��&"Olժ�ӾQ���2��],��H�"Opd��@�l�%)� ��!:��"O�j��@g�`�ѧ���QPz�#�"O�E7��Ba�	!�Ղ����hL!�ğ&?צ�w�Tz��	d�S�`�!�Ro�^���A�=d�p9SaO?.I!�$֑"���A�Y2)ZU���Q$?!�D@=l�d��R.. ���cD�!X�!�մ�H����W�f�r�ā=S�!�Da4YٵBW�C�2���d
<�!�Ĕ��0�-��0����}!�ߦ ��� gɑ!��XD��2!�!��+-�����=$o�D�t&�:�!�$�t�j���&K>cM�!���@��!�:pk���SK��H��#��<!X!��RA�$��S�PM�T����-y%!�D�C/
�@	�-!�H��/!�d��B�pZ"JՕ:�k��(j!�Ĉw �����\�|@��P?$!�;}Rp	��>8-��SEN�T�!�ď<^��1�ȟR*v�y�C��%[!�d� b;��B��8.1b��O�!��1H8)�b ��rWk�59!�ڴv/\]qE�F�!ZR�qEH[�I1!򤂟g�A��L> A�Hz2g��3<!��>�Z�����<=0�ك��}4!�$-2l��Fk�$,��	��'!�[$�\�p#״<�xB�Е)!��g���آhƞ7�4ٱ�D
!�$�4Xޠ�Z�M�j޸��"ə'�!��C�3�Tx���+���v`�	,u!�$VXQp ��ER�I~�R� �]!�'Dz�9�C͕ NK�.�>o�!��	X�y�T���$l�7-�6.�!�dK�V�^ࡢ�O t�~��W��1c���Q2%����G*� 	�y�ƍ�K�\h!��Q��`)��y2ɐ�a[4aR6J��F�vQ�����y�$]�vu��1Oq��j�5�y�E��9���c΀�Ha��⓭̲�y��~�4-�K;O��T��y�X�dfDyh��+�R�+$��y�)X�T���H� �+�
�yRaTv���n�a����oܱ�yRV4�2�Z7	�V��%*�yB.ѝC*�;��ǊK�hA D@I8�y�Ő�..��
)q������\��y
� ��3�ˁ',�|��T�6��3R"O:�20���)��H�#��/�
�"O�;��>.0,Д
�D`r�QP"O$	)��,0r��
l��(G"O��Rq�Yte�e��!Zv��Zs"Ov����F>Ґ� ��Y���1"OB�Y��M�?�2�;B(G;|�ȥˑ"Ot���n�Y�T[���L���5"O�١�� �*�U&"+�vh!#"O���fQ!�%Ҏ:��ܺ�"O �z���;X\^U
c�T�d����"O��zq�!��U���M!p�*y#�"O^�[�� vv ��l�b "O"��VKC�_�Dp�2�K�Y�}:�"O���G!CF*``&lN�&6�� "O<��mBi���딵 ���v"O44)C�w��9s�0���C"ON�AP-A0{^�8�S��xMA�"O(1a %��l�Y`-���D$b"O�p�%o:��Qe̝�n�%qd"O��� �6y&\Y�1��#��4"ORA+�!9�୍�Kj���"O��R�&O0מ`�u��!Q�F�@�"O�q�b��dx�PBʨ)��Ht"O��k�	E�8�<�B���9wԆY�"Ob\R��Pl� 5%��^)�"O����":,xH����5f���"Oz��f�Z�~���&��j�b2"O�P�"��t���@��U�I���"O�	�ĆWdI[Ч�	`1tX�"O:5���J64���E-|�
�"Oj`Ñ�ٛO�~m��E8���	�"O2��Ȕ)��i;�jJ�{��2�"O���"CB	"�U���_M�¸ s"O2 
���TM��p�_<)�H�&"O��A��wla����>�@dc�"O��¤,J9{�Ta /N�mn�e"O�E;V��R�,-ђ��eHL�ڣ"O��b���AK���N˨6.�a"O �z���i�t�W-�}��l�	�'0��j 
'"I�0��k�D�V1 	�'PR1O<I.�۷�������'��؋ÃC�y���C����$��'by[��� ��y"���8�2�'H~}�r�>z�����'V!x��'fl��}/����J�G��p�'�Z��dF�c����!K�;�L��'�ƹ���ڟ?}H�"�9Lp��Clli22E�#�Y�����*(�9�ȓ<@H���;#<����@=k~�U�ȓ<z`ј4@"���4�Q5Bb��ȓ4�������7~�&�ᆢM*?��هȓ	�Z)���$H�Ѫ�z�4��q:�-��aH�h"��b���-Ņ�K��1��N�F�{����p��qɦ��Ug�?`�]v.р��Ԇ�Lr��q%O��IZ��G&ZO�цȓO�F+�/E��¢%D� ���ȓ~Z
(%`�:ak(!��#[SX⑆�5�`qp�++ʹ��j�	�:��~v<�"���j�t��!C�X���ȓL�鲖-�-d� �va������'�.��6S�5
Mi�^�`����ȓ1b�EJ�'JX����P�|��S�? �I�q��0XX�QE5lL���"OX+��ւ0�Q�BʱpiL�""O��e�O�8�|��N�{��A�"O�	�p%�
�b@��o��`-.� �"O4aZ��A0L���mF-_ ={"O�H���5��"��%��uh�"O��Q![�b�ܰ�UJY)b|�9�W"O���&����p0�IY(5mX�"O�=��+��TX萦�Vtcj��"O:1�f�-��Y(�'a��z�"O�,�aN/r�H!��ՙb�B �"O�lpvjE� `��pq́�|<:l��"Op���ِ[7��i��4e��q"O8���L�7Ϙ���mJ(<�^�ҥ"Of�y� �4��,hcmW�<���"O�����U�^$b��ј /nt�1"O ����T@�PY�F֛m�<��"O4��)��>U3��C����iD"O�%{훏=J�����d�s"O��@��(OB!�G&ȚH�B�"O�Y۴�A���t'Q�~�Ȓ�"OB�i�nR5v�"da�*/��諒"OZD�%X���@��d�p���"O�ȸrm��9?� ����3"|l��G"O�ȉ�ňu��Ԭ�1�"Oj0�A��0oS�A��A|�4*�"O�����)�
#FL�.�.�S"O�d���?�jq��Ŋ�M��tK�"O��	#N�o��a&5yb�R�"O<��/�jlag>)x�Y�"O��gm�t�0&\�J�F��"O��J4��X�"4�$��t��!#�"O,̻Q	;TRL$G>`ؼ��D"O�m�U�ԓ��5
�Ě�?r.�!"O���6��lԮ�+�$?��"OB}���Q�mm.|q6F�C��9A"O|��d��{٘�C��R�R�Z%B�"O�d۴A^�K�q"G� �r|�"Om��6���"������8�"O�%�G�9"�^��W-��N���B�"O�р��O��0�T�T��"O~l#����$�j� �P gςD��"OT�0�(E�r%z�Ȱ,�/Q��{�"O>����PT�ʤ��"F|��"O8d"�bJ�h�*�V$R#�$
"O���0�. �4�#d%�38����r"O�<��A;���:"̙`��Y"OBȑ0`�7/����d���)�"OB�C#N�^���֧S�4Ő�"Oh���
�ۊ(0��w���"O~�Q"$4~TY�Q�]�� :�"O�l����?L�ģfM�f�~��"O�Y�L�=5'h|0�,ճ4VH�T"Oj,)��_�@�h!�U��7>���"O���@}:�P��R4��9�"O�}Q�\3-��}C���S�E�$"Ol�H�VFLp��Κ+
�#"OZ1j�%��qXX�0ЏN�l� �"O�x ��I�"ۆOL܈�5"O( ��	ӷ!���� �O*��Q��"O&�pW�H�w�C��k��RC"O�$�V	^��,�q'X7Β�9�"OT��`����Ԓ����x�6E"O�p��i�hÀl�$��$/@P$s"O� (K�äy	�%��W�`:l�I�"O2�SԮɉ*�X�X@`�.9�<�"O�T�B�B^���1勨[*�IpT"O,ȥ�@�JZYB�uh 1R"O�EiTH�3c4��aaB#M�%�`"O��;��/C��,��j�08J�`1U"O�tJ�흠|�j��Ɇ=�Qʰ"O�YCgȤl�|	P�MRB��@�"O<�@U�����O�T��U"ONTD(��f�`pB��P�I��*b"OA��*�O
1�+I	�D"�"Oz��p�Ӧx�R8���T*\���"O��O��1����Ôx:��"O����-Oz�`�fb�!9v4c�"OȄ;&/�h�F��"쁍{ �y�"O�+�ȉY�\`rT�3\X���"O��'��?	�!1aBP�0��<:&"O������a���BG�[��I�"O6)s׀/<@��b��|�~@��"O~�4o�<��"@�o����"O�L��W�q&�\..��%��"O
�+��ո/g$K,��V���"O�у��
�P�ؐ3���NuH%"O~��0#�0�(l@��Z@p�,��"OrL�N�Ao 0��g͊D��R"O`�	F�&(� t�D;��@b�"O|EIR�O!/�(Q�p�Ȩ�y�F"O�U�&%O� ՌE�'C!�=1�"OH�2U�]�u�2�	�Ş��D��"O����X�4�l���$�& �"O�	�2i@�Vqf����6�@ih�"O`L�v@�8����*\@�S�"O�!f�I�"tKߩ\�� 4"Onl�ˎ�^��j�'Bd1�"O�=��K]`ae�1(-��"O�D����+)����cĦi�P�rD"O.!	���`��Qb0 ن����"O@�1��&!XeB�� ��Aq�"OV49�;��Q� Ba�}�f"OP-)�L��N�F�E��AD����"Oޅ	��D�o�T̹�f�@����"O���A�4c��hj���?n�X�"O�)c��:A�x[��M�W$l�"O�e�X��L��#2*m`�"Oh�Bq��1iKʰ`R�#qU��"T"OX��L�j�ʔ�t�\�PT��S5"O����+U?�vd�T���c��J�"O�4��?W��2�mݮy7��j "O�)A$�&),.hra�G&�(M��"OFTZ��(NSx�a�����JQ"Oڥ��j
z�|���E�U����Q"O�P�(~�[�V�m�:I�"O��%���
` �A�kd�1��"OfajĤB�~��Q������[g"O�p�b��b��X'h�c�.��f"O�16�W(3q���a�n%\9b�"O:\A�.ɹkPޑ��A &,r"}bd"O�Th0&�V�h� �'1`z��"O�� �� ��pBs��W��U�6"O�-����=F��n��fʸ�$"O�$�歋/R��ؓC�~��B"O�`g�&��y!��/8n���"O>��R��+���X#�VY|��"O2���"�7��)�6��65l%1�"O� ��"���1��a`#�5Mvd��"O��и����p�A.%����"Ob�a�d�R�պeL�*�5�0"O�`�Qlˠ&��ps�X�����"OrTk$���=����f��[�D2��۟��&Ҭ_s����r,�Űw�W�nQ��S�!��?�]�P2H>����I�6@��iS�U$#���XE�=���Q��(h.d �!잙V�8�QFS��II�7@�{S/Q��*\c���e�'M*iI���?I�����i�����紴{��	R\�����O��Op�d9������m�yI�!SgFiu�d�C;�O��m�ԟ�n� Z�hd$D=�y�jM6xۼ �V�i��tbc��ĸ<y,����Ob7-
"s�h�OO="���&�(\�丰a:E�ph��OD�'��<�aDׂ3�`D�"K {�"(H��Ϧ�������IT7Llq���3�H�kl��x���:�\`�E/ :ݛ6/��?a�����'�?7�@8{�H�E 1V�Tٱ�â@����O���(�S��(T�J��~B�\Y�$X)Z�<Y�id�6m)�SϺ+��:oM
1j ��84����L��I�s2��ڴ�?����?IO>��o���`�)��k�,����Qc�����۠�5#�O�1PUke=p+MD=x<�@v}��O�o����2��xb�7'Q����"�ype�`�Ԁg6��>/D���OXx���	���'�����ڗ�~!'щ]��y�5n*$� 0ףԠ|8�`�Y/#��� oӄ7-�Ǧ]�<��?ݕ'�,-sr�F),k�iæ�u⎍c��U�����'m"�'ɧ�4�'zE�.O@��)��n׌�*��dc� ���'�� �ir\��;��C�~���I����t�ju���p�����.\��i��(0��P�z��E�S�>�⑁�N��@��h�S���գ,�>�����%bۄB^��~�A%�S�O|�An�W��y���N35���(�'�x6_צ�'�J�K�f����.�)� w�h�3z���We�33���?��o5ԙ���ʊ6Z�I��x�O����D��w^�Ԛ� ͟�JT����H�N�d`Z�.Գ*yj��U��ŀ �J���Ϋhj@���HO�����'A��u�B�$�~�AA&<�����/	4�Dए5n"�4�|"=��MI�(���/p�<,���s8��Xش.���i;��A�[�����敺z���'���ĩ>q(O���<����e� `�4+������T��z�iT�Q�"�x��'��	>Tv9�!&Xk�61�@$P=�7�F�PW0��Q�U>?x�)��̄�H-.��%��r���¤�}Ӏ�P!�'�op�2�$=���2WWM�tE��'�
j�V��T������Oy�'��	�M��4�f)�7�X�Wh�����{Ӝ�,���6M��"��+���7���׊�N��&�ȅ퉂w�� p   �   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �    �  �  *  y  �"  �(  P*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms��a?Aab��jD�O�,P���$�0y�x�����A��j�w��}�n�W�R��&R~��YBd�*���$� y�~`#_|X, ��o��L�#hZ�i$��`N:�`�O��t��XF{b� �v5��-��.s��c"ճ�~�Ƹ�R��!dH���J���7�ybf�9b��a��Ƿ��P�F&�?!D�V��|�¬�,�`sgb�i?�"�%̓@_����duP2��%�y��K%i�i�J�PLQ�ALR�>T�D��f?i�f��."�O=b@�V�DS ?G������_�h�n��0?I��Iڂ�8�L=*���ؑ�]�s�z�*5�X�L!LԢ@K��=)\9��_��0=�F�]�"�vT�YI��I!G�&\5ўԡD�U���T��*]�QHh������]�p�hQYB�G"{UlՊ7�#D��ٴ
L�K䱱"�D �2-94J�O@��@Bδ �)ۂc�T�ض�O���`ӣƠP��/0�jD��L-D�ȹĬ��s��+�G�����-��k�ڈ;��O���b�/O���'^�~(�<A'IL<{.�Y$�j��ط@Hvx��ٵD@&T�D�2��A�!,V9H��Fe�r�G���D�f��$� �`V"�q���S�˓I4�yb����l�V�Ha� �"�TA��`M���#c)��5{��!�L�����ȁ�g���ȓ�rP�5�ڛEC��!dO�	&���	%}(�X6 @b��a��Y�;���)��40V�e
�Rw|��&�C������4�|���62�V�h�����8@q�'`���I.�5��é|�D�ۺ��'�J�(���j���ɕ	��s:}@�S^�}Aw�ܟ2ܠ���� 9�
7n4N?���		P�8	����P�v@��l��VCY�-��Q��[n E{ @@6�QTbóX�4� �Ɇ�~2�J,")��"@a�"� IZ!L�-�y�	]5'�ҝ@��(�Ҽ��"���?q�(�$^����*Ż(l(��Ue?�r�K�}`k1��Pd(��f#��y��{�ir4�
hjR\���=���5
�v?Q���f��O��@Q�$��@��r&�d�f�#���1�}"���$q�Ț� �����G)~��%*������H�_HΌq���(z�bi�C�'��4" ��k��)�(����EI��$��͈Ȳ�Œ8'%
%K2#4U���0k2�� ���������O�]f!� �a|���W�;M،i[��IW�#�^% �҆ɐ��J��v���~���IXFr�8�Q�)?
@��l�E\!�dٛ'i�*�KCRi:���ͶZa�x��S��~��f(6�)��ii@.%�I�{8�ԏL�$�����2)B��"!i�d�����Ed��°��Y��1�0�+T
�YFB�=,�~����)�n����3�Б���I3j��rd�6ў,��*T$n�hЈ�!]� �6����ȓ$�Z��� bBE�&��d���$D��7=:N�X��M3��J�i�	��̞^4�2P��6�´���S�'QƀRp��;R���P'F)H�.!��'��4���R01�g� xt|�8�*G��x�#����o�Y��gQ1O�٪D��:R\��f�/V��4�""O�b�@�TY6�G/\�]� ��"O:P��F��'j1���20���"OR��!�CY:��-ƆO}�<`V"O�����+]�Yr�͝�]�5;`"O��C��,���R!�*v4�@"O���e����4���|V�\ۤ"O�P�#/I.��zU�y@�M�G"O��iҎef`�b��z�41ia"OL�P��
eڰ�B��>h�Hȡ"O<����&�&,�Co��`�����"O�aQ�ٮAf���ݞA�a��"Opy����L#��1BM�4%�U#"O�,�l�>p���$/^IwbA�c"O��؅��&Q�H�aM�>?�dr"O,aYgi'A-��BR�:=���Qg"O�����gH���S"ۼ#�H�5"O��@�#S��I�D�23��_�<�MG�:�m ��/x`�hq��W�<��hڜ&�|�3����"@p�"V�<!�o�?l��aV`��a�j�ծ�Q�<�uG�\W ��𩛔mY�iNTQ�<��l k�8u���֐<��%y�e�c�<A��DIU���'�s
ԡ#$JX�<���<�
�H�I�X��a��o�<��\�-7�!���>Uɀy��C�<�ŊҞ10h��> ��Z�j]�<'�H��z}�Ì%�� t�M�<Qe�9��@`r��5<xt؆"CH�<�QW9<ī�-�n)�Īs��\�<)r�Q��,K�� +���
3E�V�<1s�=f\�zu�7�Ig��m�<�uF/��|�4k�+22n�t�b�<�pbV�D���I�Dg��|;A�a�<�W��3��s�	�t��}ZG��h�<q��ƌ65.x���k��5r��K�<)s�
	�j���zP`C�<��h !�4Kfj,i5��ˡ�@_�<��;yFy�dϩ�l����S�<YÈPV%Y�@ͼg~9��OS�<�5BZ/Bf��{��Գq#�!���CQ�<I�i��9�X= �)B�z@0��Y�<p/D�'"ȍ'�%��cU�<�4��#m8d���K�jn:<{�I�<ɧ�
T	|}Х(īL��0�A�D�<Y�j9�p��q!��ܹ8R��h�<�q�W
��:��$^�ʙ�EF�a�<��e�,gV�l�����\XȔ��B�<1��ڦ"�䛱�ײ��=�Z��ȓ<��(�Ǧ��*<��.)a��E�ȓ-
�CF ѳ5a�c�Ο?q�����S�? ��@BC��B�a��c��h�"X�"O�a����4�@K�B���}��"O8�ā^!Of>p�3�C t 9Hp"O��G*B�zD�4!��$BY��"Op��A #+:�� ���$._�D�"O�9����8�Q�M�DE��j�'��*H�9�4�fEE�_�6P��'U��8D!WQ�\HQ�^nU+�'���1`��	h,㰭�Y��Ls	�'����͂�mϲd@@$C�V��r�'8��ʃ�ޒ;e���$�EO�>��'Q�H&d��b{�0�T�p˄�	�'s�PC�-!Nv�h���}�Y	�'��};'�@؅ic慭t�� ��'���s#�G���k�c,i��0��'�Nx�" O69J|��iׯn�^�K�'�l�z4�R�2L��` BH�pN0�'!:̩s ߷r
��3@�"|ծ|p�'Gmh��6�^�B#�x*�x�'�+o�61h (%�.!�U�V�/D�` f��L��0��8T�Y  N:D���� ԛH9��{� ݔ�����&D���M�mJP8�癢k���R��%D�t�%!Y�,@�i�v�X�9ž�Zc#D��V��Q0����o��P2�<k�d D�� S�@G�����Ֆ.^yȆM.D��A+�9Æ8��F$�>��`�&D���5̏�u[̑�Fj&2[4A$D�D'���+J��p��#g�2�1!-8D��+A�יఽ�T��_�m`�1D�|�t�;;8.<KAM��ۅ1D��p�B��JΊ���",)�<�e4D�|�*V�Ghn	�R� V�t|��(D�h�T�\��8R$����K�f5D�x*HѰp�u�@�b���W` D�j#���>p�C�D�|8���"D��� �I�q�M��Gn"<q��!D�4b�)ރ�f!���P2���j@m/D�4�P�Y�Q"P�2�O�!?,,��7D�t�J�!>T^+V��5T`�i�6D�<É�/�nhhuD�#B"��F�2D���I>���S3IC�	��4J��5D�<+��1i&�ɡ&l �L���E3D�tᦨ	{�``2
ϯ`?|�!"�1D��xR�^�����O���"s�?D���!!��m$�I�ɉn��B6�!D�`('�M�N��p#d����M�W�,T�pr�*�@����2hֺuؕ"OVaʰ��t�`��p
��=`"O(��LP$aVV�q��<]��"O�aJU�[�?�=��L֋xYv�bR"O����*,�,@��V�
_J��"O�x��k�X���"�l�n�Hq"O����+��"��vȶ�Pq"O���O�%��ՑD74�|9�"O0���x/)��O�2���J"O��c�m�ϢAc �H7'�2� "Or�y�̘�{NѨe&םUBB�k�"O|�
��%0�2� %	&@ȑ�"O���𩇡 G.<�&���t�"Oq@�I�l�\ �B��r���#"O�<�7�ɞm/ؘ�oƱP�%x"OH)H���@�Ne9.��sz����"OĔ� �ק�r�{�NS�Fx��&"O� �X��N�C�j��5��vq>��P"O��a]�- ��kN
*prmi5"O��f�/�X�	���2F�u:�"O�Ih��B<&�
��6`<ƒ�k�"O �r�Ā(�5��-T�G&��W"Oz0���ә/"l�L 3�Ģ"O�8v�s�NԺ��:����"O�A�&^�81h��t�ڏ��$�A"O�A��dY������GͰTy.�֎{���/B_X��J��!h�؀i�̋ ;���@�=D���I��xz$��:p����<D�HL��X����ؘ��=D�4�hC/VD�(��׾�\����1D���c�*����
	�N�[�,1D�p�T�N���l�e���Z�,,�e`2D��@�J�q��(`!+�z�<�&�1D��P��w��XD�.��0��*D�H�
��q -H%��I��;��)D���g� �?ab�i@E�S��}I�,(D�L��	�_��9�6#
��:D��)��˱H�Hd���D�RJ�S�'7D�S��=6Y���E>aT��'F!D�x"��ѐ�j�zjN�M�X��� D�3��A�z�$��%@�8���+0�1D����ջ:ڢ�B��wv�]�� 2D���	g	Ƒ�wj�1�#%%D���b`F�gyn$�fǋ�q�~	��I8D���T?���4(=�����8D�1�%U�{o���*�C�f�X"D�<�%2BW��"M ���K"D���eN�']*mBC�ðSx&��!�"D�<��X=Lu�d�򩀼-�"x �@!D�T��Hߺ�HT蜔W{4dB3+$D�����={�Y�"�P����!D� �r�¤��K&g�q4�a;SO#D�0�2�^����ĭX����ej%D�t�c�F�<*4�&�@��׉!�$��(>l�2�T�<[bI�.�!�ć(hЄj�-�t �S�!���[��y U���`��M�@!!��!#Lv�P�ǒ���D�c!�Č�J|8��_7����:{�!�䈸�h��򎊴 ?8\�[>�!�]+�:1"Q�I|%��*�+\1!��M�U��JE}	h;Eܭn!�Đ��x���~�B��E�Q!�$�_u>9��A'�H �&��!�DL�,Hi��f
�~ɨ��U��!�d]�����N	~ D ��%v!���������3^�L�Bp�	d!��-�}�ģƪR	��Y�J*D!��ҺsY�H:�'�
S�@��e�,V�!򤎿b��� B)C-�QY�D^%N�!�d��GG�p6�ͷ>�!�5^6wy!�M�-P�G�0k���4D�c!�D:/t�Ȱ�)�]�@U�c��S�!�	'�T���Ȱf��DI����#�!���}�$�2�"�t�`̹��1	l!�Ǜ.������ծC*�j$�\j!�#�$���n�q�*�qFe!�!�ēq�"���'��v�L,_�!�ǣy�$A��DK�X���fd�6�!�D��5h�q9�LY9i�m���Z�mN!򤐖q(�����c��	
"S2!�� ��YC%N�o�Ha$�_��-Z�"O
m�ǩr����cA,lF$�V"Ou� ��T�
��ͼB+�Q��"O8S�a�HoFMA'FF�$�<��"Ol<!��[4H� �g�'|g�|�G"O��qA�hS8g r@E��"O�`��F`��81����:;�M�e"O�y2kӜ%y�,�����u�S�y�L��0!v��-�,�xt�K(�y2�F$E��qeO%#�m��,S�yr'�)dH1���I�$�h�� �y�ĝ�*9�y���mn�Kw�Z �y�n�
s~Cbd�"j|X:N��y~"����
^t�=j���"�y�"\�������[�h��˻�yb�L�k<ܤ)��N!U�H�f��0�y"DՍ>�D���Z�i��4��N��y��*ֲ�r�j�b���� ���yR��0�p���m\7G�t��)	��y����44����ד��X��mP5�y"�R�
�ڡhӄ	z�24s���y�oY8NJ�aǠQ�_N��j�7�yB�˭7~)�Ώ
w(�����y�K�ml�@��L�Jxu���y2DT�%v�!����i+.�y2��>��Â��z�����H��ye	/l�t�D(F%$)��ē��y�,�aH5(4eJ"xp!Cgπ/�y�)�Vvx�n���8�q�[e�<YaD]!5�СG��eQ[��z�<)ƍ_$1x�]%�PL����Hs�<��`�*��Bg@?Y�S��g�<A���cĸa���)z�J�de�<Y�*��26D��N-5�P1F�Yf�<I����Vd�Q,C7����&l�<��͊X�@�q�P�;�,sÉFk�<����C�t�2䞅~�)K⢛�<��/@�R��|����LdB�*�*�f�<�!嗍i�L�Q����Y Ѣ�dZz�<Iqi%v�*T �K�8�r��Nt�<�s�QY�����/"2Mra��w�<��%�0S4�jf�0Ht�Bc��]�<�TŃ�[;TTA�Z�7_�i��i�r�<AB��5q��i��g\-K.n ���j�<�U����y���ڏ\��2#�M�<� m4���cM�Y/TAb��J�<)���/	z���F�'t�>����G�<9$�Ƃ�ph�#Q=��Έh�<oR�}1��镎�D/�I�Bmo�<���b�b�B[ .t샧f�k�<�&Nƴh`���"p�$��m�N�<A$�	�:��R�	C�]��� ��S�<9���2&ּ��k�>f ����a�t�<�@JVj-���!��j��(�U,LU�<���?���!�Ο3u ��w�CQ�<QF�Y0��`�O�tl�"��M�<����?Ճ��N���s���J�<�c��$�j�Y��;)�� 3�@�<B���q�y�VMA�6���"W�x�<��ME�'�j�뀮�0h.Hԛ��v�<Yr��r�D!�#�,J����g�<Q���)��4��l��Q��{���w�<u4
��ib�ʇ�72Z Qb��r�<Q�'P Y~`�&H>'r ���,v�<� 
(	�GɈe����M/T�ӥ"O<���CF7,��
�6\��A�"O��a�NS8V�j�s�H��/� �"O|j��"�%�?D'x�yc�A��y"m�L�X��4Rv2�dY5�y����� �`�)Lš�-��y�䍘��艕E��Q�tY$+��y��է=זѲR�L8:�p`�ā��y"'�.)&����9�`A��`X��yr	�<0�J�QC74�Hg���yb��ZLɸ�8)j�#�M��yr��C�8��c����9&#�$�y�@� ���m&�6��I]&�y�B
CE�I���M����k��ɟ�yr�X��	��*P���V��yB�I<B#�)��D�>U�n8V� ��yJ0� �86&ݶ~1��h����y���=äI(���oJą!Վ���y�#N�#��/Ċ`:���f@
�y�)�9U9�s�T�QHErD��y�o�>�4Ht����P��D�y���8M�5cnB et �H��y����
x(cAK����F��<�y�JK�,�B�˵�+���S+�y�IC�:m�[��ҫ �j�9�,� �y�D f�%�C��x��$�3(�
�yR+��	�	���O�h1�廇�T�y2B�T�\-��	ozT1�J�9�yB���Sj҄
eH�{�l=������y���5y.�A�u�΅c��%X���y���"
���1��Tm�FEc�$�'�y�	�>�x(P�OY�c�f��@"���y�߶[plْ� ��u9����yR)&?8�䙑��X��1�r ��y ��`��iK��M���1	��yb?�P�8p@�v6 	��)���y�`C$P�)Т/4�ZH���y"���'�<�襎Pc������y�ݙ��Q,U��A�#���\��F>l�Q�]�o�� �n׻�FĆ�#ڞ�˴%�Uk*�k��l�(��R�=���׆>p����H�%���ȓ$���+7�}�A+p ɐ�����%���>k�T(���^.�*q���jM	��ٚ 5��A�+-{����+����@�fYD��	�%'n渆ȓ1��ņ�(��h�I������)z����P@�#fD�<���ȓ7$���>z���0�Ɲ A� �ȓN@����M�'�6�C����$�te�ȓ�D+�L˓��\�D�V�4��ȓ0�hx#0��,QN\�'J��&�N���ҺRF�
^F��9mH<��5�H=(qcA�,���&Y��l��|����#�W��т��O/U��ل�E*Չ��N "��XB��èC@ P��o�6�aP肍Z���1�	I" ��-��}`���QiA�d^R ����t��i=0�
GaI>yLl��E�ʘ	(d��R�Iۧ#�.�U������ȓ�~�۷�^0z�m�Q�F±�ȓ^z���"I�q���c0d��Y��ȓ��@A��Ch;aJ�5�؇�l�|�@�(���W�G���m��S�? �T�W�G�2m�p�K\�vp�R"O��Ô��*?4�<r%��
�x8�"O��SRk��
.A�Af
�M��i"O�,��_M�vL[d�M�PQZX[#"O~�򢏂	X�(8��ċ=o4Yj�"O��P����B����3Ȍh�"O�<�Ǥ�	�F �գ=�N��"OTM�ğ�>\�1y��Z	�,�"Ob,�ҁKZd� ��@�2>}h ��"O���f���<��
۝OxUp�"OD�fm�v�F�����e�� �"O�}� %�6,a��3[RV-9e"O�(�F���{��(� �J�ɲ�"O ��`�  ��   �	  �  �  �  B&  /  �9  �D  �O  |Z  de  \p  /|  Ƈ  ܒ  ��  ��  M�  ֲ  ��  1�  ��  +�  n�  ��  ��  ?�  ��  ��  �  ]  �  � � i   ' �- �3 : T@ �F �L "S �Y �` �f Jp �x # g� � �� � 5� L� �  x�y�C˸��%�RO5d��pJ�'l��I�By��@0�'�F��A��|�^{���OM4ؐ�Їv�lh��Y�&7�C1Jɜ��AP�Hj�%+5#]/AT֝�ҍ�"�x�S(#�t�	0�� �Pp�h�� ���rI�	cUhm���>>O�|�6k�p��`Xw��dU�O������q �P4b�d��A��$lkL`����t
��Ia���9A)�9��=n�<;� �I۟P�I���ɘ(ɼ4��M7P(� �c<w���	���I�x�'���t��ϟ$�`J�4j� ���~���eFşx�	J��ß�ɵO2�y" �l/>�(fLѓXi�q�Wf��y��+N0�*�XҮ t���?I�[�qV��q�՟>0�����uH5�Q�]:ʙ�襟8�@dܚ#�()`�ҵ�,�B��O��D�O<���O����O���1�S!O2�A��>b��'h�/6������������'E6�@ڦ�޴!��	�1�Q�V��9q��w���b�ԭE{��O��=ke'ԥbhE��P�o9Aϓ�OT����f�9���������G�'wў"~z#m(@d9+�nQ��"��u�è��-�O`@����]w��"6c��M����[y��p�Ҽ1����2��W��8c���)�n���3	���B`�I�OѴ�����:�	�>���@�QS�.+g��Rte�'Jt��9�D�Ob�?�'+zI�7��4���:A�Kx��!�'�By�ЭB�XE��,��u��+�',��k��0��I�m1ܩ��'rʔ��b1{W�^������B4]<�}ȳ�Q�l���7����hO�U{���.;�  X��"
��	�$A���m�	؟`���)�y���PtFi�/�1*">C��g*@�I���}Uȡ:��I0	�(C�I�d� �*��Y� ��M�r�ȭ�JB�Ir>��!w�Կ:0@����J�V�?)1�S�c��jshޘuZ<L�S�Z���Ix������	c~��{�r=��eY�� �$��y��˅"ب-�`y2�,��mI��yB�:_���kR/I�n$(�r�GG��yb V�"C<$R��G��h���y��E�=�hY��
�����d+��
P��(���1��3B���1vz$��S�lp��ǟX��K�)��60��қXQfY[c�˳+�VB�=`߼ �%�S�>�M
�q��B�	�?��[E#��'z�p�u�ɿ{�C�	qR*��4l
b�`H2È�@�rC�'7���(5 ҙ?~���DҠQD�O^H�>Q��U�<��O��9E�9KQ����/�.C邕���'��'��6��1�7��� O���T-T7*V"��Qi<J㚝��A*O��1�cd>�;L�,X�@#od�5�rLߔE����*O}#��'�r�'W`��D{ȸ�V(N<;$
4?�I�X�?E�4A@�O�pE0��/ ��XB� W���?A��'�6 �� }���M�,/�Mj����d�;:���$)�s�0�'@�P2��R�vk�!�����=��!�	��t{��/�|�"|2qI�#>�f��h϶US��Ӗm�D~"cX�l��=E��E[
�`��	A�[��8��Z������@���'��O�1��Q�E��1/R$%��
�' h0��|��'0az,�V/�A�t	�*{�dyr��O�@G��h �*w���&'J�p�H��?Y�(�3��'T�4�'.╟�"A��f�(��2d���҈cM9D�dcu�P��x34��2�X���$D�LS@��M�^�:ԫ0�h��=D�p�Ňhܘ���T-z�|X��'D�� bl���֡T�
�`Dꗈ�<�1�)�'r^���J�-�$�.�%��0��j�<����?����S��ݡ�<C��1G8@&|�.)i7O���`�׊R00��IW�ܸq	͊J|!�䗊4؄���F��MR�c�6��P���'l�'=BX��g�62Й�C�\� w���q��K��
�'+��˕��!��;a�I�G�VM�I>���i��S�\��O�j�Xa�+3����DV"o���	H�	��'6�!Gx
� N��o�!5��4S��
�V�����'��Џ��	�X�䅐�I�k�&�S��Ǎ4paxR���?��y���	���5���ʬ�����y��g*. r�I��",2&a����?A��'�D���6Pir�H@�8^i\�*��d��nA���(W���Ǫ�5�< �*ӥ$���Iɟ��ɽU�t R"�"��gk�r��B�qT��5�W 8B�}����/��B��9%�s�ݠ2S�ѻ��T�K��C�I�wĵ�%BB�B)di�@� V\ޣ?� 퓍h�)�� ع�b��!+ߖ3X��NS����D�Iz~򏒟,e��'�L���������y����5�T�B�v,�"�y���R>��A�!RZ�!�f��;�y��Tkj�!��<�8؅�=�y�,�-_��S1C�42�%��P���s��(�7��i��p($(�-Z��(PZ��h4N�����Im�)�S��.M�G����".Si�kI3D��Q�F�P$�a��њe`x��F4D���%#Ю��И��.
�~q���0D�� ��
�1l�thwb�=@Ht��F�.D��� ��w�@�x@Oį d�Q�L.��P�'MU��'
�A���w�C��]�������?ɍ�L��JfQ�)��x��bV0p�`�*��!D�8:#i�!j��)0��Ӻq �a%D��b��-.�b�卆z 5 &.D���)M�j�Rq0��.������-�O$��Ig7��+�7��s��_PƢ=��)r�OT�X�F��B�t�� �O޺��'4B�'�F���(\�R��š�a�z�'�y��U),*p�KSq����'Q�P%coz���銫DNr)��'��|!f�R�i�L�S-��-��
��dGb�O�j,�p��:tDɁ����P{�u���Ex�Ot�'��-"d���%��R�6L�%D�B䉔�+*׆L0������!8v���'y荺a�c��y�e� ��u�'�T�r�`�Sd��u,�u�Y �'�x�)�N�W�δrga�p�$+O�0Dz��T&,IL����� }�F����5"c�99�
��I��%��>u�â��X8�{sk�X{��3b�*D�li�I��Ut�����3*Ȅ�h)D�,S��/qÄ	���[9����<D���'�$��r�O�}���&D��T�;���S�KH����&>���r�'�:���' �@A�צ���:���&'{jqb���䓧?a��L�\3�ޮd�z���ET�=�d�{q0D������0^�'��Br���/D���	�Q�`)�QcLr�4��,D�PqAψ!8�I���8���P�e(�Ox��I�ls$%�R)��N������0q<��=���c�O���c'��=H�Z�bK�|T^-���'b��'�jx+��C4\��[����
�	�'QP�;�A�5��x�%*�
�b�	�'�$��E��t�t`fC� N�N0��'
�A���r�@y�֡-M.����d�~�Oo08FC\�0��Q�v��"K�����:(Fx�O`B�'����C��	;��v)n��e�!_�C�	�P<�R�X�DǤ���*�;,rC��&��0g�ˁ}j�s% ={nC�	�t��X#E�#M�9���$:��B�I�h`���ľW�TYG�Z�mG�ʓl���|�Q�f"�<yN�#a�DP;�LUyʇ6�B�'Dɧ�OK4��G��`ʨd٢­d�40��� @��D%S6%9�)RE�2S �P�"O|E�3��&��`�����C��	"On�V�I�/Y��ң��b�|z�"O�� q|�92�kN#K��`࠙|�1��΍�W�E����e%`mx�K��~Q�I`�	�����ON�R l/��i$�^1v� ��V"O��nV�H	�r�ۃ�$��"O����� `6�iӳGU!xᆌ"5"OL�30ʑ>��|qQ��&b��,ٶ�'Բ��Γ&C�Q1��c�DxR��&�ўLIK6�'!�ݨr�ؖN���Da�5^q$	C���?i�j�lx1����V ���a/׭%�D��1����ͩ�jȃ7&�'m�m���0Eq(�V	�Tc�fR� l:�ȓb�d9�'O�/$zx+���j:�D� ڧ�$Icf�6n�0�+G��,�F}��-K��"<�'�?����D�"*&<�7� ���!�ƞ7!��J2b��w����Nh0�G�I!�>0Ȉ�҇� eR�,b�`B�u*!�dH*�"��Iţa���DJ�6�!�d3`�$ٓ��t��ъb��{�剽�HOQ>�'�<!�X��dg�C��U�BA�<��M"�?����Sܧ9|Ѡ�\�0��M0�eƪP���ȓTp����r|�X�2�C>U��X��@�n1Au&V9���J�9��t�ȓH�p]��G��j��� �L	5P��$���.aY��lV��
����$�D0��$�71<�$G"~P���F�k�^���H�.�|��'N��Oծ1��5V�,�F')
I�ȓ+;�4�*���r؁�l������).>��G��@�f�:��(���XL�G	De�8�P-�;<=�Q��Ɋ�?iƉ��kX.��Vhڔy���a�Xt�'.d�َ��N2��!�uJ)ق𰫉�-/����O��d�/7b2��%g�]&�0���<c!�䇗=Cd�:D� %�`Q��u\!�d�!���
�&
B����0@L6hR!�˹;��ŀ��Ph�,T��?">џ������2G>ܨk���,�����<< ,R�O���O���-?�A���=-)���0P�b�D_�<Y��s�`��%�[g��!E�Z�<9�I=�tX�G�k գV��W�<c$S5�
�� E��eF���Y�RB䉪(�nE�󣊺�PX�#� �U���|��LZ�A,������ ��K�Sy�c	��'^ɧ�OY�Pk��!x~����ʗW��-�	�'~��ir�Ӭ�\E)`�PDd�b�'p�X)1�֠�ݣBO|N̽�'>zUC���cY��1�Z�%�b���'�H�cE쒛U5�m�6%V�2�܁�M>����">��t0<q�EK�zĀD����45���1���OB�?�''�����j��j��H�C�(K	�'s�	�S[�,;F�V&@1l ��'��8�sf�8
~$��iG�A�4�	�'����A�"Ore�׀c�6��� Y�U�fPc*X�CdU`��E2�hO����Ӫ<زS �hvD*'��'vcxD��韐���6�䲗G�5A��I�#Z+vB�	>�=���2i�t��냜n�B�ɶ`W�`	A�H*z�ah��*2.B�I�Z����I���@�b�
!ܢ?A�5m`��$��'UV͊s/��Y����"2���S��,�Ib~B��N��k��]�\�R͠DCִ�yB+�6%�dy�&	
�,���+X2�y
� ��	�.΀y��o�Ը�xf"O8T�Ц�1g�*�x�0]T�
@"Ot	�n\�ȉ��)dZ>���Q�����哮\�%��<Pe�g�]#}�0ʓd��R��?AH>�}*�I��*9�0�n�b�����
�]�<�5C�v.�j`�ę%��mc���X�<���(z�=ku�?8��m�%M�U�<�L�bP�\���6+)�؋%M^M�<��
;F�E��
�W3 �h���d��1��O�� ��OȌ�G�G����)�������'�'���>��GO
e�������t�4�RWkKQ�<�!C<`����%�ȑ5�۱�V�<ё��j%z9�6��X8��U�<�%"E�'�%I�)� �~���C�Q���R�b�ȼI�/��1"�&�D���D{l�͈�܄bFоhϸѡ���t��1se�O���9�O�I+�F���@׮D��"O\x�rF���0%�sgM�H<p�"OH\ȰA��p!���s䌲y'�yc�"O��ٔ�� iiT$ #�.�<(�g��%�h�|�	1�Z�3�<�8�Ʃk�x�$�'�Rh���4�H��O@�)�Ո�B9$l���?�~\�ȓ4�z���V��B�[e�Q_����kP�}����$LAJ�;�aJ��d��o>��p���K������Zذ��G��5�Gn�*�<٪w��|Ӵa�'T�#=E�Tb͍_��Y@���i���J������ƈ���$�OƒOq�<��sƁJ"�� �O%{�<b�"O�U����J��AK�,�t�p"Od 1����L�2��c�Ɲ'�>�*�"O�X@ƛg=
���n�(���"ORs�ٵY����Eڿ$tX�(�|��%�ES�i�9�4��'�!*4;!g�W��(��e�П���O$hp2� �7�<��+�;V9B�"O$!�E�ՁZ���S�TIX�Ӱ"O����bO%���1j��:ij �"OԸ�G٥JaHвh�F^�M�f�'y*�$n�ܰEί5��@3�$Dvў$r�O$�Z$^�	4�ʀ/ƐZ�"Mm������?y
�M�$�M	u�dP��T�[�&Ԇ�9~B�B7��_��Q2�ȇy�Ȇ�I��AQ �37��L�w��Vt��ȓ1Ŋ����Ak/��p�O�-��HF2�-�'![l	Cw��g ��T;����I�H�"<ͧ�?�����AM Dz�&�#[�����m��X!�d�3p.~Ic��_?C�̭��k�`�!�$K*I
P��$×6¸���a�,�!�d�	�Z�@�B�+,�*ڒ��9%�!�� s�Ԙ��+ �X�����<�創�HOQ>%���S:K��s7�/M=H��<��#��?!����S�'z�ހ���)\I!mͺNu�]��Eb����h�G��P��&_�^�͆�DD�)�b�ԉi�Fe
L��[3vy�ȓ=���H��ڃe�0b�D̙��d�<�!'R��t���B�:�d��g�g�:��O�#D�O�$B䉥���2m�"�&���'Q�'���>Q�
ӹa��S�0Z��-�`�i�<��L�>=�p`���R�B���e�<���=gj�1��M$n�D!K�B�^�<!��1�~� �G�t�D3KR�����f������ (�nzBȒ#~�E{�kF�҈�Rqq��Y�b/x�H��IH�y���OX��5�O��b@�͘�3�ڗ
5�h��"OFD��ɓ	"<�A[ �`�)�"O� @�8fIP��h�rr�H�0EY�"O���p��m��H���`����	��h��B�M�n�c�ʚ�6����' &IJ��4���$�O��3�V`�nLq�&2���f��=�ȓ��1£Q2M}8Tae��*(��ȓ=�L	��iÚN.�$�Q���Ԇ�0���E_�pIH�
��V5���uz �2L�f�K7O-�$�'5�"=E�Th�M��lX�iB�l���Zb
����v��d�Of�Oq���S�A�Ct��	��O�o<N	s�"O�q��@�(�Jj�4�J�"O�p�"ءiu���ɘ.V8Ȉ�"O�2k�2Y�� +،~�HXf"Ot�SF��	�f!2c��N�
ĩF�|�,*������M�c�;�f�鰅U�T�L��@�	�����O<x#��&aY�ɢ�E	�)r�8��"O�p�%N�w�2�TNNcS�a)&"O*�Av���E���c�Y�O7�h1`"O��#��0G
2qp'I�C?���c�'Yh��Յ-tbhҵ��(c��	
 ��(�ўЉ��4�:8����X�Xk��W�t�����?�t`�X�ă?"�ڭC��]+YB�ȓA����MR�~�
<�'j�*g��؇ȓ_�8�S��ݫ�r9�'�	�{WJчȓƖ]׌��"�,Dσ�
dr�E��#�'c�60�H�0����@�S�°���q�#<ͧ�?9�����^<U��TBSj��T���� lN�u�!�� 	���vmD�g_ؠ��+�22�!���Uo�P�ǫ�U.P "� ��a�!���2*�`��ǌ1���`gI�!W�!��͌]BxӇ@
4�VX!���剠�HO>}�WՑx�� ���)r��]��nY֟�O��'{� I�O��'���RU��&h�^�@Fꖫw%�����|R�'E��4o\fу',	@��	3���O�!1ub���KWx@=S&�z8��Hg���(a�C�Q#��Ozt pB�d��š@�Ȧ����� ��'&1�R��uK�H�4�j��[�U���pR�����=+�ӆd�:6��ab!&��	�(���OLyr��	M.�b��T&n�hUr3#����D�7Z����O��?�	���� �/����2c�"���Aޟ0
O�Hp��,��Ku�X��S�O)�HeG�, �5�&#􌩜'&*Ѩc�l�Z@�"Ă�}N�?-���׷p�Lia�	"W#\�(6�s�`S '�O���#?%?��'p�hI�*ʿ��a��[�4J�@	�'Hz��$�*6�\�y��ܸ���1��$�m�O���R$LK+jr�(�f�!��V.D�:��O4�i�O��/�Dۍ2�bL*��[	ˈ�y�IO��B�(vb^БF��	?�f];�
��ܜB��*S`<h���2Z�8��wE��]_�B���đ���N1���T�&=~B��&[��C�M�>�y`��T�G����B�����H�`��62�؅O�d]F-�U��O,���O�d6��ӹUWh��"I��K���YR;Y�~B�	�`��Li⌙�9�`� *��.h^B��	-�H�	j4=��X�2B�I�
�����* )]$)B�ɫ,^�B�	>��c���\Z��G%/;˓`ӑ��BC�6}�@�;/K��p�f�9pX�g#�'�䓓?��0<i`ߍe��� �q���A���S�<i��	Ǫ�6�f�hDO�<	C�BAQ&$+�O >aЍZ�-b�<�,�U� a���`��|
0d
ax���/O@�X��F�IT(pmާ!�f�8 ���o��������n٫,:�����u���������� �f�("CL�L��!CG�}:0,�ȓtҸE��� 	�8D�UX�l�,4��S�? �eHchwѼM�dbS<_r�U"O�Iٓ�CJ�Z�i�&^�C���蟆,�J1�t\���.e{l����=�O��)�O
�$ �56ȑ�sg��x�V�X�A��6�zB�	*\�]z�BAg��(5���TB��
�^���d����Т ��qm,B�I��\�!!UQɞ!���%v\C䉥B��Y2�!�J��	y���vj��dCZ�������oT,�^�*�B�1i�cA�O��:���O���,��5LL:�r��}���F �sLvB�I�"���RBM��#��NDC�Ɂ4Vm��5��ج?~:���o��|{����R�ƥ���<W�t��ȓN��T��C�0[+@y��%�5
`���'<�"?	Ӧ�g���,�������H�b$��ꓧg>�'���'.axB�T`zl�����^��pӲ��4�y����0ǎ��KƳWD�"�ۍ�yR �����P�KN|����n��y�j<Rf�a���K����E���$ry���i��1�G��J��3�@W����O&��<���kz��3����l����)V����O��xKB��>�©S����;8�@q�!�����&�d����|B�NЗz,!�4�W�4��ɠ�~��W;���|�t�l��R+ �(h�E"P90�0��󢝣���DD�d��KR�F�O��$2�n.��I3	ˍ8�`Q����]��RB?ٌ�9OR5�5�6n2X{�їg7b��e2[��-��"�PD�O���On�I$�Q�^Δ�j�.�a;��F��O4,�v�S"u�>=�]���"p �V��8�	�:�.�'��'xHآO����4J��� �Nז�
�KN�];�a�'6,]�I�x
���٨^ �aRG�2U�V����W�3��5��,̔U�O�s�X:�+>?	@��p�N�t��>��ٻ��AV�/O�HW���3�ӲB`�E�%&�?
'���ܘMP"�Dۇ�~RF�(���?�	:6����2���zD��+��@h"����'lba��	h�����*��=<)2#�1_��B�Ɏc���ᢍL���}Ba+
?@�B�$^Eڍ���Z�"��%�2/�r��B�	�s�`���ՅT��Y2D,%fB�I�~;����i����27eBB�	C���̝�yN�;Ӥ �cB䉸qU����N*@v(k i_	PC��,A�R-:d���J��ɖb9�C�I��й�MZ;.B����nC��L��(�� �v�>�P�$ԥp-C�I�e�
@+f+\/�t�тc�[��B��?'��]�LΖoJ�M��ĲR7�B�I�O&��+5&�% �9��8lX�B䉍��lJ�)]/W^� Â���!��#?����?���?!�[p e�� �c���<W��)�i�b�'Z��'>�')r�'f��'�0��֣&���aƥO(jغ��e���d�O����Od���Oh���O,���O����̟|�6��3!&m��X���¦���ǟ8�I۟X�	ܟ��ğ�������#��l0n�AS�
>�d�K��ז�M����?y���?��?���?!���?	��ZI�X���ϦJO8���0����'�"�'��'�r�'���'~2��8���ps�^8(~�	3PB��G��6-�OD�$�O@���O����O��d�O��dY�B����ʲf~i��_"9!BAn���H�	�����Iӟ�������	�0���ٱO�#Ӿ�H�	��?�~|��4�?1��?Y��?i���?y��?	�E;��nbԍ��K{N���ÿi��'v2�'lr�'���'���'��ഩ�B�zL�Db�	Jzp�
u�j� ���OF���O8���O���O��$�OT�Aw'ٴy�<�Ec�_C@��`l����	˟��I͟|��ڟ������	�i@fH�B��4�Jb#հ;xt��ٴ�?���?1���?!���?����?��qZ��t��]xμ�����3��i\�I��'?Ib�̘�CA����P�f��D�6
o}�T�\��D�'�?�'LZ���e],M�J`,A����s+R֟h���<��O2��L�8#�'���ÝA���K$�w���-�28O�e��.X�ў���<lǿs���I�������'e�'��c?��	|�? ��UjФ)� �r8/�L��"��<)���?�'$�.>0dQ�B�N�U29:�ڹu!(ʓ�?�e	�h��1���ҟ�cR1O�l*�n���V�B�
5c�Q0Q���'b"��:&�  ��d�g�:K���c��O���'��I�p�?�'ڸ��v�^�����2�D���?i���?���_5�M��Ov�Ӆ��^w(�\0���0"�TJL�"�A�����ON���O����,oe�5`�m>�0R�<�rY�x�'���	��6^͊D+]�dp�A���Q�.��ʓ�?����yB��h����i��8�<x��E�"a�oܠn����?�p�O8�I>�(OD�[v��3�V1��ҕM�l�4|O���'���y��ʒ����=G�"�'��Oʓ�?A��y��{c*���S�����%�:�)��4��$��i�֘S��O�"�����ݙ.�ּE��=J`b,
�:���D-����dK2|O����'p�H�`��O��$�O���'��S�`�<�㒓=�|x�K+B���G���<��O��d�O���P�L46�5?��5����G D�K<�I�J�0����g
/�?��)�Ī<I��E�:��� 	�(�L-㶄�4�Oh�'��'�r�?�y�([�f�V�C�N�cRp��u�<1,Op��O��]���>���d�9d>1�Z	R�X��?J>D��Fay"�O�4�	y��'Ny�O�)�vHKTK�;�t(���'�B�'���'��O��	��?a �Eg��T�^�{1R�����T��ݟ���b������O�KSl�������`�yn
��QJ�O2����7I�7m ?���Ƚdf��Sc�D��Z�bͺ�,K��b�9�?�-O��O���O0���O4�'9z�c�jF�*蓀$����O����O��$&���O���f�g������]�2>(��G�O��D8�D'��)UN87���(��HP�x�vyh�\7l�(�U��OE+v	և�?�V�.���<�'�?�%���:�ڶ^-K r!��*̀�?1���?�����dE}}�' r�'n �@3�R$J��1k�6|;$�j��Ģ<���?�M>!�^2}�����i�	v��� X)�򄖧S& 1Q7���e��i>)j��'��5�.��)�+l	B�)���U����ʟ���ɟ�	w�O����2i^=���{M\x3s�#��"�>I���?����'��d^�n��� kB��H�M��	�'(�'�j�H#�if�i��I�V�?�Y��ڨ(�X�)&H%/�{CMS%�'�Iş��Iџ��I�����>:.ĈҖF2������"��'F듗?���?�J~Γ4M�@#WH�`�p�e�w,�/O ��OړO1�2|�蝅p�R�a#�\8}�y;���3:�7MTHy���LƜ������$Ŵk��(�s
�HkRx3VJ��-�D��O����O4���O�ʓ<��	�4�X ��ah���=נQV�럀��G������O���t��k���T�d��N{��d�/��6�;?iP��@��i4�㼃e
�2�=�j�>]�@���ߟ��ڟ$�	��`�Iٟ�E�T�ɯrp,\�C���87�;�$[�?��?��Q������l�	O̓j�>L�A��X_|$��(IF��$�$�Iџ��	J
H�n�T~������D˖j��cؑ� ):D"�1��Iu?�H>�)O8���O&���O��KW�z�ʤ!��=��ݚ�F�O��D�<)�Y�8�'B�?m��
Ƈb͘)�W��a��<	/O���Od�O�c�v��gܲr�(��m]��9FkG�-� oZ���蟖ha�'��'IjL`�b95>\)"%g�_z��A��'d��'b�'�OB�ɐ�?�b�� �%�'Wb؝�v��~�Z���O����OF⟀�'�b�[� � ��k���(b��'G�(���i`�	�ED:P�r؟@�'/s�pr��`��JE
��t�����wyB�'�2�'�"�'��?��3�%I�DU �	�	�%S}��'���'.��y��'-�DJ�g�k�G��H��(IRj��!r�'{�'��O�BS�i.�$�H`�z���Oc�}�'�I�dz�Ƽ�"�������D�O���3�L���V�L�`�ue]*���d�O����OX�g���Wy2�'�<9���,�0=�7�B;C���1���<����?�K>ٗ	)j��q�V��H�  [bm��Z*k�x��K��(	�i>u�`�'[�ΓZ���E�<bۼ��7/dFjX�	韤��˟l�Is�O��dY{���w��2h*m����@f2,�>y)O��8���<�Qo�9Yk���΍�i�7i�֟��	ɟ@�əCx%m�g~aF�Q�]�'Wn���W�,d�~� e9Gph�I>	(Or�D�O����OF���O��p�*D46Ȫиa�5��͍cyb��>A���?i����<a��B�V��ܘ�h��4����d�O���.���!�|q���F�D%��� Q5��T�i�h��'� ����a?�I>y+Ol �D�@�1�����"�?"6�+p��O<���OD��Ox�ī<y]���IW�? lj6g�s�J�pPV04�,rD�'U���<������*�$ԳT�ݪ�1�e��>ix��x�i��Ɂ?̤�V�O�,�%?=λm�⍹�	�[򖌱gB�����؟��	̟���ɟ���j�O�xt�n��H�ɢ�-p�� ����?A�������	ʟ��<�T*@0^��j��B����a�K�|�I��T�i-7���R7M/?��¬��R�I�(�Ǜ�l�f�""G��?�D	!���<I��?A���?i�o��M�8p 	b�NZ�M�3�?	�����|}"�'u��'!�1?���G�ξW��glB�.����d�O��(��~z���0����T��|�FYȷ-K�UJ��7�H��z���O
�I>q�M�h�2|����	j�8�
��?����?����?yM~�)O����2N�(�u��-�($�fA�%M]���Ol�D�O��|�'M�N� �DȘ� ӂf���.ɘF�2�'��a��i���(&���i��HA,0�SK��m� ��'�8P�T���I�����՟��I쟌�υY��@�+#CM�JA0� @��w���ٟ\�����&?Y�I�Γ^�fH1S+\x�ʐ�ɓ8����ğT%�&?y�����y�����E��RR�����4!D~���^ʼ�)��O��O���|�����}��F�>{YpU�#m_�Bz7�'��':\���O|�d�O��V�|`^��7m+Li"[@nV�kE��x�'����%��kIץ)0���Q�EjZ˓]���Xp�Ѷ(M~"P	�O`�' 0��n�',�8��eX:C�����?���?���h��	�` ���̟pn�%�I�1� �dq}2�'M�'5�O:牒����!��Ap�mR�A�g6�D�O���O$�� p�Z�Ӻ���^��� L�?> ��A�8$>����Y�cT�O4��?���?1���?A�I^r�@Ab�y�.��J�`�(e*O~��'�r�'%��T�'x� ��e��d�g�4�����Q�������&�b>�����W���'��!� �j �[�v��s�]~yB�o����ɺw��'��I<;�x��g�J�+0�Pr�NG�n���	˟���H�	��ܕ'�@��?���܎	��ai��O��)�s$�7�?����'��������<�¨:5���F���tE �B���秊�'O��$\azJ~��w,j�
X�<�и�����Q���?����?����?A���*��$���f��;�bּ���1�'T��'e:�����O�b�8�d��� �q2�[�LV�T�q�=��O����O�,	�E|�N�s�^YQ�(�m��E��!�/+#d��v�H�j����X����4�����O�����f���Mϱq�Ȼp��9�R���O��t|�	jy�'��Ӕ)ߎ-�
���%��.vJʓ����O���8��~���#��ЁO���E����> X2�A̦;*O,����~�|"IH(~�LH P�DZP�I)��	M��'F"�'Y��4T�L`��|aj!�Ѧԛ5<n�(@�@:8��������Ɵ��?�)Ob�dQ�0�Yȳ�>�N�cc��8lH�d�O���	g���A��˓��� pص�5�T���O_TD�c$�'~� ��䟨���x�	Y�4k �	��OF#y�V\�Gc�g��I������&?�����ΓF6�)"�A��D�!�Ϲk�z��I���%��%?��f��A��\��DKR3{H�����hk<D�	9N�$a���'5��&�d�'���'���Rc�s"��C���)�$�'�'��Z� ��O^�$�O��D�Ck�l�t�μyXTa���qHr⟈�';B�'��'{rԸ�*�>}��D
�KF�[�K�X�l��+H'&�L�lI~�O�����y���bR���e�>D�p�k ˉ��?A��?)���?��Iq�\�$�F:1�(I�K�\��D��O��'[R�'���$}���i]\��P0�(8 �U�Ba�OV���O>���	6�??� ��~��	~�Q�jY">]m�HÚ#�� ���'��<����?	��?���?4�A�=�~$���Z�
�ͩ�O�?��Ve}Q����~�'+��1��''��S@��1wEJ�#*O�D�OؓO1���*�e�8)�lQ�4�� ����Ri B��6m�oyoΆJ� ������Ė��&e9�eP�yj��36/��H�R�d�Or���O�d�O˓��IΟ Z'E�>/?�HR�B�FG8J�W��h�	I����$�OF��`���4Txx��a�eB0θz��؉Tu7�"?)��h=<�I?�S���GB�X�ĠU�L�]�`Q`�@�	ş���ɟ�I͟XD�dB/}eh��.�<C\47`L�?���?&W�P�������r���l�� H�lQ�D V[;�&���I�����{��n�M~Zwˎ<�CH�af���(7���3���6�fVk�	Yy��'�B�'⫏�s�"Nu	`jN��@U���'h�U��r�O��$�OZ�<Z�-��)�F�`aM��fҮ�z�yy"Q�@�	Q�S�	�qf�4:ω�@6� S� yg�Y�֜� �T����f"�LP�	�9�m�⌌'������^4�%�I⟈��ٟ`�Iv�MyB��O� �k�LMW��:����Ym,�g�'��'�����<1�4�I��ċyh,B��̙������?1K\��MS�O`��b��zK|2�
�O?�	����Z���OKɟ��'_��'
��'B��'��ӣ5�z�z���F�,�vE\"O����'�2�'�R���'�23O��G�ÿ*$����ԓ7�\�s��'�b�|���D
*��6�O|�TG���Y��aQ<"j�պ��'wt���P��#2�|�Z���I`��6�@��K�e�����I̟���|y�G�>����?a��YR���E�(`$��`�B���}���P���I̟X$�\ʳH��vK�����V=�{r�wyۼ[��	׾iZ�i>Y��O��ɼHd�t��b��&�O�M��D�O���O���0ڧ�y�͖r!0���钐- �p3���?Y�P�d��۟(�Ij���y�nO$t�����nC�X������?A��?���z2��P�4����?
�RxI���u�hw��c�
&�n%/A�o��p$��'�'eB�'��'������,6L�p�M�*Д��P�HA�OR�D�O ��"�i�Ob�I� &ws�9�(T�w�6�Q��<A���?�H>�|B��؈Qɐ5̳iZA0��]6�l`��Lx~r胶(b&��	2pC�'c剐r�ܲd*cQn�h CHڥ��蟠�	ǟ��IX�'QF��yr.��<�ЄӇ�#�I+����?����'r�	џ��I�<iR��:,�� ���:Ppu�rF�=BZo�M~�%Ke���E��;��A���j��-�7LW�+O��iE�'���'�r�'�r�'�>����"� �__�a�w��(��I�`��Op���O�D"��="�t����P�P�QQ�+@�:�O���O>�ŵB^@7�5?�;"ʬP�L�	��u�P� 5� V�\��?ɰ+<�ļ<���?Y���?���i"�k��D���k���?A�����M}�\���	j�t���>���S�1d�4��\��<��������܄�0��6=?�MQ�hϡ2�LA�X�* %I�)����?�� �'z��'��`�I�!�fqKrl�+P�l��U�Z��\�I���Iϟ�&?��'�D��}m�c�%� �@���S��y��'[��'�O�˓�?I��mP*�q#���y#�A�2����?���kθD�޴����!蟬A�ʟ�Ћ3�[	!�B\��#�|h:ucC�'��ϟX����l���� ��H�Ԍʇ �B������G�o��IП��I֟l&?��	ޟHΓM����C`Y���m�� /�,0�I쟄&�0&?����ܦ���!�r��.�u�ѩ��Q�p�	9\��y؝Z �|%��i݁�'�?���M}�t�T��4S 8cJ״�?����?!��?���OS���'eb�'��m�c+ �b%�p�>�PFJ�r��':6mK�g`�d�O���G}�4��I�B(,)�T�Aq���@���F�'�rK����c������:��{�*�ə$�r5x�ÂnN�H��6)����O��$�O���:�'�y���,(��V"~2�駪4�?	�Z���	��0��Q���yr�\�wU���!k��_ؘ��&Ƈ6�?y���?���|x�D��4����,�[&���;T��/R<x*����df���f��������O��d�O����O��� _�>�J6	�;@~-k�oZ�4,B˓~<�	�������&?�,l�R�	%'T8dZĢ�H1>)�1�'A�'�ɧ�O�j����.-�d��t�؛>V��3�:�ź�O~�h��W"�?�uc6���<�uS>�
�3�Q�i�Z$�q�-�?Y���?)��?������w}��'h�h��"H�q#�4'za�0�'L��$�<���$�;( #�ꑗ5�LH"եڇ7�՘��i��	�j)�ț��O�ȁ&?�ϻ@H���+�#x�����.z�4����\������	��	T�O�(yB�)h\��&�)� � ��?���YC��XyR�'�1O����C�.��h��o��@ו|��'KR�'�t	H�i�	@=���5[J��.Y�[I �2�Q+�$>��<ͧ�?����?��*9x�:E�HJi���G)�?a����\}��'��'2�ә%�3cA��E;P 颎ĹQ2ʓ���O���O2H,2E�ȩ9��Y �)Q2	Q
	0 C�"8Y�y*���������lA��}{B�O�c�Oм{J 1	���HP����OD�$�Or���O<��2ʓ)����~�@��iá�dݩp���?���?����'�I�������K��
��u���S�d�Ɵ��I�_wZ�mZD~B��� h�a�9Ɣ[���2P��ڄ�^/���D�<Q���?)���?����?q͟ Y2f ��j���r�@�;=��e�ʷ>I���?����<)���yR	6W�	�aJO-u���c���?a������'xΕiڴ�~2�zj��v'�'kڨ�bC��?��`(hv��IW�Ity�O��k56�%X�,,���c1'�X�"�'��'8�ɇ��D�O|���O�$aeC��M��b�
���6�	Jy"�'n�|"�Ӭxn������YW�* cмR�	�SAd�Z���¦!���J�v?��'8L�W�]0|���2j,��h��?���?q��h�b�)� �`�$��H��=���OP�4X��'͜��?���?y�<Ox$��ʅ'<��p;�U���@��'m��'h�iK2��&���A�ᄺ;�4���q�m�*�V���E�>od��|�U���I��P�I؟��	��ː�+�p�Yq�\�K�V�ayң�>1��?a����?iP/�n���A�&|���ߗ��D�O��+��I�$ElN�Pt%�Fx���`IA �����@:�	� h�y��'�t@&�|�'��P:u�?KD�#�JW+Yg2h�S�'���'�"�'��Y�l��O�$�Cir���T�G�P\��j����OX�Ȗ'hB�'���'�V|�U�R�!���U�[�z^N�#@�i��	�o+�=�C����jۮF�a���O�eh*ɔ������֟��I��<�I���D�o�b?�0�G�-ĭ� ���?��?��S�$�I�\��E�`޵��+��^���E�A��" '���IƟ0�	�[<l�a~���w��u��GZ,W#l8�ߛ��$�k֟�r%�|R[���쟔�	�� )�fH���ռ�
%d�ߟ��	vyB�>��?�������J�A1�Wq� �Ʀ
`u�_y��'��|J?��Bŝ( �&uY�f�<?Qx�0�IT�DВ�U�p���z2��O��J>a��*�Ĭ;'-��uaT��sM�?a���?����?aM~R-O���I�0��s�k� j=�Q�H�-����OD���O:�$�'�b��nn�)�CIѹ> ���F�F�IF�|lZd~�f/:���S ~���5�h�J��S�O�^@�
���(��<q��?����?���?A͟x�HG��8�8)��CDϒ93K�>q���?!��䧝?��y�a�(,�PS�̞�!�j���?��������6�Oȑ�5��t���� ,Mb�'P��ӑ�m�6� �����O*����Px��b�&9ǈ����<���O����O��,��DyR�'���a�F��);�bF�: ����<���?yI>�*�|��;T�!49��{�[���P���x(t�];i����p�l��IEB������k%�@�O�M���$�O��D�O���$�'�y�ڹop��`T���1��]+�E���?��U���	ٟh��d���y"d�0m
M�4(bb �ȫ�?	���?���=�F�ش��Ċ�0 ��)���uا G�,#��N!.���87�����$�O:��O��d�OZ���9Hp��+���`���Ȝ'�6�!�I��d�����%?牽G�^5)��V��-s�C
3
�4��'6��'�ɧ�Od��	��Ѿi��+v�V�e���3gC.:��OTu�fN[��?�-�$�<I��Ŏe| ̱�Ŝt�:`�ch#�?1��?���?)������i}2O|�FfR#�=��I$q4Pyq'�'BR��<����$@���:���!���Qa*1U����i��	���,��O�M$?	λk�V��Æ9C�D���)\$����ܟ��I͟���ϟ��Im�OB��q)O�RZpe­~�|r(O\��H^}��'8��'F1O�ɡ��
�B��ŋ\>Y�4�`��|��'s�IoLou~�@:�D�+B%t�.48�E�o҅9�,՟@B��|�\���	ٟ��	���3D#Q�K0ܝ�0N�bV�]a��G���Imy�A�>�)O���*��͝�`@�!�q%TAϺ�@��cyRR����ӟx$��O����CY�j`��Aa�3Q �c�K�&�F �fD~��OZ\��I0)�'Y�i�HaJ�ꑀE�(b�B&�'b�'!r�'��O�	:�?��h��B����0ꂬ����c��㟸�I�P��|������ODEA�+w2����2C�
��m�<�T!��M+�O$
sg�.���!��	���<�C��4@Cֽ�"P۟�'�r�'M�'���'��S��hC�Ƒp����	�	<��}�'6��'�����'�;O��;W�܉`5����	��q��'U�|���d��4���O�4���m	��:��!����1�'ɼ ن�[�8BA�|�Q��S�d*��6rm���3o��hb���ߟ������syR�>A���?���x��E�����R`x�$Z�1�����T�D�I��&�DJ#i3Z�ұ�2Ie~�1��DByBKG4j�(� �Ø%�O�,��	%��$N܊�1��!K��a��%�c���'��'��S�<Q� T����f�����t�&g���$�Ob���O��0���<��+�1u,bX"�ˉ  ���������ş(�I��r o_~�-(�����+�-�
 K�tcqō)��p��LRe�	iyB�'g��'���'��'q�L��V����h��Ʌ����OX���O�������b}�
õH�VСe.��;����?Y����Ş�4��G%�|Xl-) ȁ
�|�����M�_�P��G��8��$?��<�*
cID]����&� ]��9�?!��?��?�����	m}�'�4a�Un��z�+4��$� ����'�b�$�<���?a�'��X��R:Ix�X&�D1Z�U����M#�O�h�U�J9�����d4�x�3͗�,T:6�,�����'��'�B�' r�'�>� ��U��%Lg�yчw�n��_���	?���Oh�D�O�c��cN�&^��D�T�X�W[�hz�j"���OH���OVx�	bӐ�
�d�3�o����9A�K^�*x�+�&��S���������4����O�� �̈��n�N-z0yC��)ef���O��M�Iӟ��I̟��O-�Y��N� �
���!4��!�.Ob��?����S���8�8Y�7��%bd�ag�;V�L��A>y-��3�O��	B��?�gb,�d�� 8��rB��m��q�mC�8�����O��d�O���)��< �'�8� �Aκ8aL91�����?���?��^�t���uN���C  |�	�c&F�n]|��'s�Aa԰i\�	:
�(��Ocb��O� \1�����c�E�/f�U	�����O����O
�$�OZ�,�#,\�[^���G.Y�E�ܜ�&&��$�O��D�O��?)�I�<I���)!����=6�!T�����{��r��L�anZn?�eo)Mо}!%�G\�0�e	 ԟ�Ҥ�[SWbLq��RyB�'��Ȁ|A�eA�+N�EP�E�͞}!B�'�b�'�I���d�O0���O��t����6lˆ\���5� �	wyb�'���|b�Z�qE�����9U�<� ���5U��	3�T��B̚��L~���h�<%���ɴE[*5!a#"�l���؟���۟��Il�O��D �SN�8�/�([C��G'׎ie��>	���?!����'i�dZX}J<Z�DM��*��K���'���'�� �4�i���z�J�!�O뎚�|m�Y�bOՕq<�;B��'�'��ğ����4�Iٟ�	�$�(�l��Pǆ�k�(ߞU�8�'듼?A��?�J~J����i3i^)L�$�89D-�/O���O�O1�b���eX�U�&T�J��؆ŏ2.�V��H��?3���s�Zy��9C���E��*i�A�BF�2�'}b�'M��'�����D�OiI����P���@���:}6T@0��O��:�IXy��'�2?O�*��;B~�� �7	����6@����,`4��
3��d��g��ì��tYRu���A�!��O(�D�O���O"���O�#|J7��r�L8�������a��\�	Ɵ���O��'�?	�y���f;t�3"m׷(��8I�� ���?I/O�
ujb�d�la�y;����VK�4��*R.Cbx��_
5����N#����d�OF�d�O���ӊd?|�o�vҰ���i���d�O@ʓ\�I柌�Iٟ�O,���?��4���Q�WHdA*O6ʓ�?A���S�)��H�@���{(�0�3ea"y�D��n`U��O��)��?��I ���j�c���EnMy�@�!��$�O���OL�d5���<1G�'��cS�D�"ľ(qW�:H�������O"㟔�'�� /�, �׹c˒��Pf�";�b�'n���Źiq��9%�Ƌ<��
�0ţDi�Ā9��e�%��d�<	��?���?Y��?�ɟ�I�����sĦ��AػZ�$R���>���?����䧌?����yRHL('��}�t��w��H�/��?q������ڤN뛦�O�i2(ݵaj8����D�����'�҅6ƃퟴK�|V�|�	���ؿU1����ް�B�%L۟����p��ayҪ�>����?1��qX�$��1Gf�d�g+Q1+�� ���W�h��S�-V  id(=3���3	C�� �A+O�l����BʀT��,�)�&�?��!m��#�π�7�|!ri��R�R�z��OF���O��$�OТ}b�'�X(�#P'yF�1'�L��k�������I۟ �?�'"`<�G1:�I�w��	�LE���?����?��D�)�M�O����B�I�3vn����@�Hph� S'�x��K>I/O��$�Ox���Ol���O���U��,$�mɁ�o�a�B�<�TW����ڟ �Iu��4S~%$���>%�	F�I�k�`Q�+Oz�$�O��O1��� b�7l$�M�<�d���2n��`)㗟��a!�0e����M��qyb�Wr�A�#�gm�W��'���'��'B�����O�`Bd�ȥV��$��(Ġz]
I�w��O��-��Ry�'�?O�dҀ�^B��Δ�SMȭ�3	�
%���<!�N�"����@�S��[��@�g�B1:���U�~��������I�4�	�\�I��F��ݍ$���w �q�b��tb��?q���?i^�|��ӟ@��k̓[T�b�*_[:��0�x��&����ߟ��I�Gp�o\~��m�$�'I�<z"�K5��x�k1@ӟ�C��|]��S�l���pc�Q�8F���`�%������I}y�>��?�����i�0%j�ه��s���as.ؘU��Ieyr�'^�O�'�e
5J2�U��O�j�-����J�нCrGP5h��ʓ�׮�O�E�K>G��,�VhpcC�Cx)Hd$���?a��?����?�K~+Oz��ɠ] >}WZ)f:)�|�$�<Y����'��ן��s�ِ���Qp!�����"Ee�ş,�I(~@*�lo~�d�nkP�~
��:H�bA�PDg����&
����'X"�'���'���'��3� r�3�%�82_tqbvk�'��ً��>���?	���'�?���y��,��%�B�b���Y�]4�?������'7��X�4�~↗�_�x׫V�] $�p�l�?���~�b��i��~yb�'&�eZ-q�0L{��Ɩ>��(u�\"s.r�'"b�'�"����O��D�O����$��z��Eo��r���¤(�	Uy�'��|��,x�j�)]4o1Pd1A��|��ɧt��)Ф�G�wM*��|����O�T��'��i{�̆T-Tx��G���Tq���?I��?)��h���ɚUT��Y1&ܑx�̂2
3V���CS}W�$��F��yB���X��ᛆF/��Y���?����?���sX��ڴ���J#w�ؤY����k�OQ>�L3�dQ<J���|�T���I����	֟��	͟ Pc�=o�Ҧ�B�4�8r�*�ny�>Q��?�����?�F�F� MB k����ũ��_����O��2��I]M��X�ÔU�F�&��dMrQV�%[T\˓{�&5qq��OxQ9M>i)OL�j Ê�	2�X��͙��x�Ä�Ox���O��d�OZ�$�<qX���	H�n� �j1�`&��D��ɟ��?Y(O�5?Q��p�b�K�)��cq�OZ�Xl�Y~r�E8?qB���:T�O�#s������ƩF膤��*F3"P��'w��'�B�'���S}"�p`A�/s,���m�/
����O��S}"T����v�xBJ}Aᇿd(ԕ���q%�$�����$�	;O�ln�a~� ��RP$�hvaP���ͳ�&%�&�r�n�̟L�Q�|�^�b>�I�s�LL� ��]�=+!/X
h�0��OD��O��9��%��E�Q���a),� �TBy�[��I�0���Oâ@d�֟z���̑�'֬�6l�>Jm���Ϋ�����B���?�`�OHȡ�o�V(&Az�c��5���O>�$�O��D�O.��P�-\r.E��HP�R:)\ă䮙��?q���?9����?�+O��ĝ����	<��2c�� /�2���O�({C!a���Ӻc􉞔�bc�1ʃ���a��vΜ�h��9��F���ȕ'/r�'���'�b�'��ӏ8:=�s�B"N;hpu)��jD�'r�'$����'7�7Oh��B�ȫ=$�	�o:�J��D�'D�|B�����2כ&�O�ewG�A}xq�F8J�^=��'u�Y�A֟���|�V�D��ܟ��r+�F���N�#�6�S�k�͟L�I��x��my�e�>����?��
�X1A炠 оTA���Eh�K>����O�$$�� ���S�B��ۆ"R�g��ʓ �}��h��M+���T��?1�'���& λ%u�!�p	$fB@U����?���?���h��I%�t�{!-�	��B��P[���O�(�'���'wr�|R�'i�M�ih��C��5=n�[D� :T��'���'1�K�i��iݡZ���?͙��;a�� � ӣiz�xB�Ϡc0�'�I̟��Iӟ�������I�� d��@ΊQI� @<~K�x�'I^��?���?aH~���C�N)���͠\/P �stz��/Or�$�OʓO1��tbRǆT%(�X�䍌Pil�qS��52 (���<��F�o���������"`X����%�� C�vF��$�Of�D�O����O<ʓ��Iԟt�UI�~��!��ڙ7�P�j  Iҟ��	P�П��'��'@��B�����
+@�a��I�|�ði���$$eS$�Oir�'?%�;?4�R)��T�А��� ��H���d��؟��	���^�O���i��/����2�0@\�����?���
��������ܟD�<��+ @�@@�����5�Lq�6��T�ʟ���֟����B���'Zd)��@s-.�Pj�/>�1f�J$C�0����'G�i>��I͟����6@�i��� DG}(��Do$��Iݟx�'t���?����?�ɟ�� �'L��w�:#���S���'c��'ɧ�$;�pJ%�͒d;)�j�+OJ@bMQ6"�,f����S l@�̊C�I���`�T@R�RV�����^8D�	ß��	֟��	H�ByҦ�Oy�%M�Wl�t �#��U)�'���'&��d�<	��H�j�І$_Ȥ0H�'��jW����?�!��M��O�!i 'v��D�S�7����@�:y~P��ӸM�F�d�<����?���?����?qΟ�[�#t���[�H��I�<}�j�>���?�����<����y2�[ƒl� ��;����s!L�?�������'7}h,q�4�~Ҡ�IȘ��_��t��o�?I��	d}8��O����4�����?F��L�U�D�1�HY�5&ʣ-$h�D�O����Oʓ�����	�DI�.܊9��(�GСIRU����l���d�O���1�d�<|�,�7p ��ru+$'�˓ܨ�F��7D0�(���� Q=OhU)��=&ޤ�,D��0�'b�'�b�'�>e͓o`�����|i�G �*E����$�O����O��hΓc]��:�j�ԅ�(M
���s(U������	� �z�o�n~�J	2u��O��y�� �dD9�� ��9O�1#K>�,O��D�O>��OJ���OJ� �]G�"F��iY �Վqab�T���O���O>�$7�)�OrtHHISx
�%�ύL6�d:6��<)��?�J>�|�$��z2тQ��
Q*�zŕ;l",kٴ���@�|���'1�'?�	�S�6l��F��(M�2��!v�`�	�������	ܟ̗'��ꓹy�%�1J��_�l"�.��?����'�����I�<93���־�JDC(������$o��n�L~r*�>�@E�0�r�
�n�oN�� B�C�o��aٲ�'�r�'���'B"�'>����k�⑐G��- �4��U
�O����O�d�'���'���OI{ � �>2�v��ց�#��'���'��'�u������Io��
R� �v�n���H�"Z��en�/!q pR��G	}�>�U8X򾭲҆ {�T�p�j�K!�Q#�l�%5Yإ+�Q2Rİ��3W�E��M�kΚ��JU.��҆
\/Y}��&-
�eZ�d�%��%{��%2�H��\z��Y$}�����(�3=2�h����;sOn��-�5w� ��Х�����7e��K�*�v�T�i�ȪP��1ggęSe�T1IW�����N�[^6�p�ʒ$o��r��Ǧa�6��&�=�9�Y+}?"�z�E�wf0Rȗ.{:�����B1	�15Ԝ�z^<�q3r
I�x�(��`�xM�2)��
�XT"	�g�9K*���#ꉓA��T��Dհ>����� @�f���N����㇝�S�L�,%(��DO�g��X�Ԗz_�0`�	I5A�����Fɏ2 `)9��	|��$����x�LH��ix� 6L?U��8@A&�.��ge�*@��;F��R:�D��j��B"�a���i�0��eL���J�`��Y{Ǐ�F��@@I�,y7��U&"L�1 ��9�ď1BA���D9|�&h����O����O@	�'@���pAT$��e�G� �69H��'��'���'Y�'��(U��Y@4͕�|����� @���1�Jޟ��I�M[��?���?)7Z���'���V��NYH����5t�e��'��$��'_�'&�S)e�*����ibҐ'﶐06CO��֠I�I
�M���?a��?	�\���'i"<Oʬqui\����&AY�<vt��K�0��o��D�O����O,E�%�l`"�5��@��OR���O^<�'��͟0$��r��B�mt΁8�n�	qg�D�s)�Qy��Q�>$�b�y��'���'��S)o�D=� ���%p$��1'ԻG�T�DC}rQ���IR�	蟨�	nkD��(H72ז����p� � �DP���؄�v�p����0�	w�S��MG��"�	���H���ȟ4�')�|r�'(b��:["��('�萋�.ϐW9@��U�r��}��'��'�r��m�~�j*��jT��3|Jf�Idc߬1����?�N>����?�	\Ř'�b�kQɔ�nM������(|�;��?���@�Beϓ�?)fY?�	ԟ��I�nչ���"
��!Ǌ��'����ʟ H�N�\���t
�����YF, |�1j��*�?IFa�<��I��f�'���'��ſ>A��[:8�t��uJD�oO|��	��?����?�$�o�'��!,���L������קs��XP�N�ϟ���Ms��?���?QtS�\�'E"q��a_��������M��'��@r��d�|2n�<	�#��i�׆%�Ҝ��m۔B6��Ըi]��'rR�'V����O��I9$l 9�*J�(����`nM�N��⟜�A؟$���j���Iӟ��\e,��,%d�a;F�:8�L������	��S�4�|bK�T��y�� ��60r4�+(�' r(ɔ�y��'"B�'y��?�I!������K1�d��FT�	ן���M�IWyR��a��u�ݡ{��)Z6��#f���'5 �A�O��'�B,O��SCp6��5�	$�x����[ws��$�O���/�Iҟ�'&t�y`
S��%�u/ʪFV4�[�e�\��Ob�d�O����<(����1v�T�QA��!��!QD��&(��d=������'7n�YL� S�"J�4��"Ōg��İc��O��O�1��<�-�����O��݉?{t)P�"X�YzF b'��9WJ�OD��<)R��t�'�����)֢<������Д0�`Ѫ5�'a��1D_���I������d�Iy�̜y�fŢTޙi�t�8�
>3"�'���U�#<�'f�1��F	���ђȍ�_"��͗����O
�D�O0���O,�S���xD�K]�kZҬB��F�	o剓
*P"<ͧR���͓�?�����(?d|�s�E4�Θ�'��YI�6�'r��'��E)�?e͓1L�x�g�O�&kX O�t��̟�$���I�i ��?��w�*pZ��;lܔ��MI45~u����?�����|ډ�bӌ~JdIk��4>@A���#�'���@���y��'��'J��l(����9�F��)Df��[B��ϟ��Iw�Oy�-
f7�%�V�E��Ic� P���'w�)�O��$�O�i�<�O�b�JB�����e�+;L�����?)���'r]�,*�L��!"���
5СI$ ��3J���Mu���I˟���V� ��I�O�у��o�nUaD�Ŷ���jD��O ��6���<�'�?�ʟ�ꚨqR\�!��fv��D�'�2�'��-��'E��~���?)�w����PJ�<ݮ%�v*׹D�:$S)O��Ļ<I���?�J~Γ#T��e��}���pG N�y�(��/�X���?������'���'��T8�x�Y�d�%�۾+��æ�O���?����'��Iޕc��� ���DHAf�����,��8�`H��'�rg|�>���O����O>�'����@��y�G퓻D��ұ�ܶe2����Ob��OʓO�I��b���O����\�c����oPD[�����A�������\�Oʓ�?!�'Մ�J��,J<xDpv��D�~�A+O*�e����K^t4ͧ�?���?A�C �VU�נ9y���熠�?	���?Q�Y���'��Q��̻yع`v�
/�"�8��'j�D��'[`��'bV���'��'���y��I*t4�䂅)^� �k#hĪLW�>a(Ol��<i���?���-ެ9#��V3	I�͂ᕷF*(�A,�<Qg�<���?����n��T(����(�t�^\T� �gi�?�)O���<���?��~�<���}�0'Â[���C�$�g#������?q��?����(�@$�O,�Δ���ɻeLց���g,U�[��'�����I� ��h`��O�� �gb�'0�d��Z�҅��'��'��1Z�'���~��?I�T E+S���7^����g�rTQ/O|�d�O��Н%��D�OB˓��DOF�e�b��
ץ����ׯ�?���<���&�'=b�'Vb-�>�!�E�'�y�ޢ�5�p���?1���?I�g��<aO>�)�(4����H���j�.�j �UK�>t�D�O�]m�ǟD��Ο�����D�<Yr��6^zAz�*_�>�P$c�N��?1�˂s~�Z���O��\��O"҉��8���3GH���U7��6��O6�D�O"�$ Q}2Q�����<Ib��$m�b�G*I 
�+֨��L�	ay�Ȍ��yҦ�����'�=��9K5��L�^1����/|�`�W�'���'�����D�O4��y��6Z��E�$?G��9��Ҏ�?��?4hΓH��ϓ�?I��?y+� �3v���(O�q�G�-b����O(��'�����'�R�'�R�L�q"9�"Ċ$f����	Ñ��	�'�R�9�'���'8r��� ��B�{N ��1`T7`�Q�',�؟��'-��'cҁ��y�"I�v,���Ț1�dZ��G��l9���'�"�'!B�O.哅����O^�)�(\�gJ���Ǜ0T�dtH�(�O �Ķ<���?	�`)28�'�$���}�QD�)26r�b�S�d1��'r��ؖ�y��'H��'�?���?����$���S�Qm�)r�d�����OD���O:�11����'���I�*p6�P�hK0�<�@T�)Li�ܷ�y��'s�6��O���O��dT}�ș�$�6�4%��#s�
(@�FB��'Rb�Y=�O�ʧ^12�Z�
ҪQp�����2P{�#߼�?1���V�'n"�'��/5�ɩM�̑`P�1G�������ɠd����	o�II�D�]��y�'1r<��.�y������2&���DCg�z�$�Ox���O���>9���yR≋�t��#�΋nnx���ͻ�?1I>�pd�<і���<����?����@��
k��i��[�Y�QC��?���j�'�r�'��'�(���&W��l���@�>e�|!pS�<s�f�0	r���������l�t H�q4&I�AG�{�)���?�p���O�O����O�T�ǈϮMJڼ"�
:l=NXQLA�=���MV�D�O���Oܒ������9=ą!��A#�Z��C�4�ؓO��d"���O��Ӫ�������<��l8nb�9u�R Z��} �2O��d�O~��&�)K[�T�'x��ۇ'ڑ?]��r抏X���j0�'|"�'R�I�Q�����v�G�	��H��˳-b�ͱ�H�O\��OB� �9O^���H��'���',H�86�L�4��f�@�6<td�0�|r�'=b�~�"�|"1�j8��\�1t��R�$�5^P,��'U0��'J�ne�Z���O��D�O*��'��B�R��Ȼ+V�}P�����?��Z>H|������IX:VO���PB��7ٚ�r�mޏS�&x����Ox�$�����ğ�	ןĩM<1����Y�1ò�c�����
�O��H�%�O��O�˧!�1��?ه����t�2��4L|��d٨���'^��'��1�$�O:�Dy�4���F�6�d�Hr�K�4�����Ob�O.��r5O����5O��D�O���3)��i�m->Y�Q)"�$���O��P�����}�0{�pĊdD�2���Je(�8h�'�L(��'��[�'���'���?�S5+@"jx T�.�e�D�!��O�)&�(��՟�'�,��՟\��`
��z���n�ujᣚ]�,��8n�	ꟸ�	�� &?Y���E%Dpt��AI��,
8��<���hO>ʓ�?�R,NrtG!�8����!=:�Γ�?����?!L~��[?1�I9/X4A%4_�dYQB�G�_!��	˟�'r�'-�`���y��'e��T�܌$�W����ǀer�'B���y��'4�ꧯ?i���?aḟc�x�8��P�o�	�2�L5����Ot�D�Od-�є��'M�S?`���vk�=��h0��ɦp7�I֡�y��'I�6��O*���O��$�S}�i^1/��3V�d�@��i@�4��'�^����<),��1����DY3�ؓ&cp��4HN�A�b�d�O0mZ���	̟��ɾ��D�<��(��#��e#g�ς6��#�JW/�?i7��<QK>!*�$]��3O���Z�����kp�J6���l��p�	����	����<����y2�G4|�0��I�(*&Z��H�?q����DǴ]���`��	�O,�$�O�� N�;Eˇ���:��-`����'���'x.듰��O���y��]�kd�1��c-�d-8@-B���!]\��
wf����O��$�O�9O�5)� ?�$�*5��+���"�O��'��	���'�2�'�R�F).����&��)q��x0%bE�J�T<�'E�d�P�'G�'��[>�	�ܓ��0cC��C�ꆹZ�R9�v���$������g����'H���샎0F��u�\�i}N4B�+��kz�S�'B�'�B��T��~*�R%2�U,g�d��C�ƕ(�$�����?�N>����OdM��|�$Q��	��al�pc�'�2�'a����'��f�~���?i�H�6�8��PO�|��A�/��qN>��0=��['��� iEsWP��C��B��s� �	��M3���?���?a"W�XH`D;>P�2��t�4���OD�$�Oqy��Q�4$�"@�Y��M2Gr���pg�5W�����'�hx�`�d�O\���O� '���I-9 D���5G�^,S�n�1����ɥ2�#<�*�hT�@1O����1X ) �	�ZcT�����<�����O���?a/O�ʓ�?�'����T ��h]��4L٢0�|#�G`�'[�TF�=�yr�'N��'��pQŹG9t]�!��7AX�L�0�'!��'��OHʧ�?�*OJ�!���,��p�-�)t����"�<��h��<ՁP�<����?A���B�OV���g`J�!R�<�dA�6,\!P����d�O��d�O�O��Di�0��%��}���	�`��\s���c��O��!0Ć'_����O����O���^=�@�@y8S@�(�OG(&T��?���䓰?��#q.���gi~ų�O~�$pTh�r��a	h���IΟ|�	G�S�����O��Z��xtΙ�p@��>:�('��O���>���O����(`gqO��i'�9Ea�E3g�W*��$��'B�'x�X�'����~����?	�e��14�R�G��y��	�AД�H>����?���^���TbW�|���lQ�jRE��$�?9Γ�<���4H�v�'"�'�i�<�%=@�I�$ݚc�A��I�ğ��I۟t��5��򩝠W�aȄƀ��(��F0<�@�	�O����O����O&���On�����s�$٠HNs�zlatM_�r�^ʓF�2�Ex�O�H�A�'RC��0*
-"%����O�n��6m�OD�$�O~�d�Z�	I��'Z��Ȅ��3T�}r��#$E�(`�$D����Nx���O���Oy�!��h/��9�$_�`,����O����O�˓����O��O�y���Ap�Y��Õ�1n�:�.�$JN�H�Q���w�ˎ*t4Y�G�	�<�ءB�Ǫ,Ę�"��
,p�+D�#�X�:ҁN<\5v'a��?I��?�����&����!$C��:�{v��x?��P��M��y���'R�'�'��	`�,�#��>�85�p,�/1�@̠�H?\�t�A�V��
)�b��t�|!c�"�H�J�.�%%�l�GM7v��R�9ㆰƈKU�,!�n�.{ը̣��0w�Д�4H=b�^9��7��P�G�NA�|��Z�z�Ǩ�ar:82��G�X���ؗ,�k�����$�,YL��	�w�
9PF��uZj���L�t�(�*�_ET�R�"j,�*�%4a�j���� !/o��Baעhl�s�(�c}$@2(~^��5 ܣM�ؼ�%`AR��9�b*��H���:�E�yh�Q4��%��̟T��gy��'"R;�X�oR8c��їM)������z�m�4m�n��(wx�,�w#�Z�Rl�!�̦DY�T��g�|�24�H?��+#]Ax��*4�lӎ@Q �	.�tH�fG܄Yɦ ��؟4D{��	0 {�9���+�ƬQ���5��C�ɾa�FM�7�_�0��h޺.kz�'ABꓢ�Y�s{���'qr�i�  ��K�4Av�9��Z�DTVq#Eɣ<Q���?Y�P�0�!�@"�� ��\�R�Zw�@�7Sje��E�Df��(����:�8 ���
�ΐ{``�?A�2�װK(�Eq��@85����.�"����	��X$>1 hX�3�b1ϛ�]a y�k0}��'� ��$U ^GZ�[�H��Tg�X��P)�� 	�~��I��{F��� c^�na�'e�9`�k�>����䧨?�ܴo��
�]g�4I'���\���'p�Ѕ�ދd�@q�bv}*�f�8:Pa�9p��#�5}_��#P�����CV�vq�����0|2�/�Q?�5�2	:i��QW�\F}���?�������4S�dj��_�~��E97	˅[��A� #D����%�?M���r�˦�F��0�	Ш��u��-"5 �e��s����R�O(��O�����M��U����PyB�i��	Di�Pj0C�n�	rᔌCS������9O2�(
V�R�3�	�.�8����
�b�piÑn���q��>�-Y|u��ǒ��}®A0l8��j�vܞ��o��~�0︡�I�,D{��'�Y)U��h���j����wt��ȓs��@�H�|��P�R/�}�L��:ő��'��L3��T90��&��mc6�Z8^�xQWH��1������	kyr�'��8�&5J�iP@�EG;`�*\R!��U������xmڱ'��s���yK0t�ã�!���$A�cK�� �i�$ꁰ��x��*)���X�KDH<y&�d�֐AW%#��p�e%^q�<�WeΑy)�����'�b�`uL�b�$�`�=^��#�i���'�f�U%T &�x%�K�+�*�1���	8�~��?���?y%���?��yZw��RS�`:�pR��Z?*r����DX�t!�>ӳ�A3@���CN�Y�2�2�c �6	���[�P�, c���
C��<����'�R��ȓj/T��2�X��L�A�޲` �i���7�~bf��e�� ��n� C����X���	�Q�Sݴ�?�����?q۴3�tqЀ��;t�t4�wF��Xؑ:s�'ȸ:t�I;\	��O�Y�S	b���a�,1���W.�;5f�LqV�qo%��S�O�B3��6(	�QI�d�D����O�EIp�'���' ��S���p��Ϩ^+�(9č3K�:�'���'2��r!':oHXYf�߉[l��@��$�W�O������ u�V�АɑFl�0��OT���O~dڔ ������,��Ky�iY�I�g�2Oz����HM_Ɣ
O<i���H؞�3p�B�r'�=y���g�n4am:��=�a{B���zm�׬�u=B�P�ȋ��&�z��ISX���&+��M��
�e�U�P���6D�����??�y���O*q�7���l����X9���tH�9�jyX���4�f��g�K��M����?�������O��n>�J�y�LM� �ʅ�9\�����$�a�����M� >K�b���W[.����Ey؟���a�쉚V��)wd��@�Ô�M>N�cc��kH<I�jô ��g@׉,�8����v�<�g�S�o��8��� {b�"�
�v���X�[���b#�ip�'ߛV��0T+:=�Nܙsu���	��g�˓�?I��?�G�ؑ�?A�yZw���2h]�W��M�����4bl���d��w��>5�ץ!b�鶪ڦ��z�	:�-����v�~*N!h䋁�+�d8k�Μ�[w��ȓY��țS-ҷ[<
좑i�4������~"D�%R���\�Iʞ����,b T1޴�?����'�?�ߴC�҉H��A	���F� �I:4�'��H���'`1O�3�$Y�zVn�;'����
�a�aܲ"'�	�c>#<E�@]��~�c�^2DsPHd�����3�r��M��y�^�H��Q8��K4�B��,8���v�J!Zk�U��(]I��>y�SF0�E͛�p������ZX�C䉾\4ls�JQ�{t>Tr�ŝ�CӦC��9xlz���j���+sʡ�7FF�xf��IQ��O����q���C9xq�͜%*{D] P�;D��:�O�.D9�!�<r<�i�D9D���M�Rl�$�p�U�����7D�d c��,T�����*��DE��2A)D�@Rs�۩=�X@ ���z�tep�'D��e��.0VQ ��J*u�8��6D����݅]��(�&�"��J5D��+��C�|�f]��&��R�qu�3D��#�"OT�qt���D�ǃ0D�ðț�X��J4�Z$�T
@b/D�Xk6��P\0ʇ>p���!&1D�IF�K�_V�`�dÛ,A�V�+'C:D�l���
��4m���b�Q��;D���5�:e�:�w��Hv� �#D��4i�4��Ed��6�V<��'D�$�$�=�Q��,.�ĚE�%D��1+Gt�⡈��������a'D�Xr�"\,[�@ԀEcBW��pl$D� St�%��U����V�ɉ!�D�i�~��%IE=l�0����!�d	PzeR'��Is����E�O�!�$I�m],�KM,	o`�l�ݏFe!�$��&��}#�O��y���2sG�?�!�Z{��p����0��[�E�}h!��  X'm)
c�Xŋ�X��S "O<�YV득~,�)�����3"O�ɢ�&�ihv�8.�Zo&�h�*O���� D�VӼ\�A'N�<cj]�'�J�9�� )/�A*�'F	1C̩��'�T՛���hmR��$��<:*�b�'��	Q�#N$Q��ptL��8�(�'�`Qf�$����&��C]J
�'?����͙�4�q	v���8��'zLPp���*"�̛%O�)�:R�'��!O�� �őt��j�|Uz�'7nQx�c�RЙ;�� |� �z�'�j�P�(X�*�0���I��,$�R�'g@!(W�V�K"L�����9q$ҁ��'��9����#���G���;�8�`�'0$)�1ԁU��ZټL^��''��2W�'5'\�BՈ�:^U�5�'�����~��DO�(�@�ȓ_ʴ-�q�[�~���X��r^��ȓ`�X1�G��-=���I�
vo����4%�]�g��<9i�ݩw�Z�"����ȓjJ��d��w���rB�S}�d��U��m#����<�´��:�مȓi�ޱPƍ�,���2wE�v'H��5�yv�ǔ���G�ۉ�$��+���&�#!��s�*UPT���ȓ6j��t�3@�*u��'�W�m��3�)
c+F!t���gVQv�,�ȓ\[�	�G��9L�J��e�R�GU�<I�&�d]p��qC��K��<�6 �U�<ѲC�c\-�Vʘ:,���)�K�<���R�w�\���F�b49x�_�<I��ܤ�p(2�
������Y�<�$��#�r�����a.��t��T�<1R�"H��#�X�ZN�:�\�<����Ji�u#��G�2[$(c�dZ�<��f� �*��t����:`Xs�<�%�D{��!W�ĬIe�Ā��Ei�<�!�}V�<3�n�+`G�<����k�<Fg�'$"��w� &^�I��ٟdsR��qO?aׯ�
pS`�r�&.�8�z�E�S�<هK
���x��! ��*E��W?	�gY��v4LOF�B񤞄@�xZؔ�f�K��'a�E��ƻf�N�Z���\	���5�
+
j����S����ē�Ќ��f�%uOx�R��Ť7_���>y��b�(DjcJ��g��5��4�vD���ģ:eV�#a��y�k��DwT���S�?��d�$��i�,x��;4��-Ɵ����Y�<j��B�N��xq"�
%a��\���/lOP�L��۱3;��E��!$5^}��9��+��^�H<��#�$�� �'����tԉ,NL�`2𠈑�{��zU�ز�]��2a��l�iA���U�n��T�1����瀌,G�U��J�IG!�dš:��	9񎏚d���q��Вn�X ��-�?A�/�G.9�)#?��-y�Nϛe���a\SI�aλV�VrreO�P�b@%�
=J|����P�r!�W83�L�Ч�̤tΐдb�%k�v�K��~��t�'LO(�Q���W90�X��'J̥���]�Tk3��,V�=�`jؖM�,�kG�&�jo�`�� 
2eB%�r)�z����t��#ѯG�^���ς�n��1Q':�lԃA�u�<�,��5Eb	�&���;Ћ�),��h���!�y�.���l����K�S��(B�Tf��CT�WR�27&#M�"��$��'+*Mi@��8\ܨC�j��J�0�s
�/�Y����h��l���2QTR%�Ra��q��JM����2)�m�`�5j��Hx`
�RR\ϻk�ά����& �јf��j�^M���5P�2l��&$0ꔅI"`�yjh�k��W��E�N�'�h ��%�^bu��%4����`H{�i�<yV�T.d���a�h��x��o�r�'�@��ET�:k �C��ݎ?��	��Sb�m30F^�I��x�A�\z�-#ƛ7 d��ʤ+M����g�3��O`�E��b�`�H13�`��>O�H�f�4T1�<S�耴i�d��O�B�(2,�#Ҽ�˥��V�? �ѫ�̈́�^F,���hZxd�5��?	�H��ɷg
xh�2$B%VnA�T�]w��TC���O \J��5L0� '	ȵch@��C'Wd]�4c� q���˒�<P�A'�kL� +��D�~�oQ�-N4:��'T�h�ڔ�]�8�H��A�"�L"e�F�O�ȍ�sOT�`H�	NA%Q�d��L?�|^B�BEDW�Az��� N�c��G~"�*#�.��ǔu^9�O��4SG��J�ڀ%B�K����i3tת}��,@ ].��D�-�џ,��j^g�xlQ�N�	�(����)�d\	�"����)�	� ���@�#��y��cE�"#��c`o�<N&�3�	�&>TB�	wN�h�,��Iv�3EGC�R�ba���Z�!�
��6���	�S�f�]�z f��BL�%IX���7�Y�2C�ɧ<���b�	�j%�-!�e ��t��J/3� ��v�>E��'�&9�� Ю��DR��� b<�=K�'.��y�E��(|��M�Z^�-3�'Z���� Ô�ּ��ɉ��X1pd�.��u�𫉷�D���\G�Yh���Mk�"��W�6���,p|��`#D�<�ב^ɚ1b `��K�ި�s.<�tz��Ĥ�- ���|*�NT3Q��!���Q����dCs�<9#GS�!������rX�tk#,�2v8�I�!;H��ҧ���� p����F�*
�t���MC=�!�D߫ ��)5�H,�t�
U�,��D�P���� ���p=�SJՔ���:�AI�f%B����Mt8���#�5��n�c�~��2A4�uH�� ��C�	8?r|д&�& �I�pI��ud�"=)�E;<�}���T�K}�����,i��q2�I�'O�2oYi�O-����2�"�%�$@t���'����EC����`k��uP�mhsKI�[1�3H>a���OZ���σC�L"	��H�2�*T"O��`*�|ꭉ��ψ
��m�X/� �"%�ym���1��4�%eۧ��yræ�@]����	7MhȜ(����`�b��D��uX"m�:g6	�a�����dZ<{w�d
ד*'V,8���C_���`M߇Me4��>����f��`�4��C�0�@�BK�����~l�p����sBB�	I��C'ܥn}��"#ĳU9�����>s�U�Ot�KA	��wq⌳L�쀟w��� �i�1V!�l�,X�A�'$���*��z*��3��-��p����a���H��ē2N퓒τ�{��Ov���dA4"��*�0,u�����'�h�P&�O�Z����</��T����aH	�1+N�%���F[n�h���Zt���V�Kv01 ��'ᠩ�� �/k�Oj8��!�Y�$�I��H���2�6)p�ě����hd,�	uZh,ۀ�)M���5>h�у��w7 0�j$��� C��<�'�@��!�h:p�%>��;C&ht{Ɗ@�H����8[�`0�ȓ/��� E�}r)�r���aq:�l>�Hc5��/g_�Ӻ� ��p���&�Ǉ���R�_5Cw������y��۲f}�Y�qe��V{`��a�\k�)�ɥR�R��֩�Ƚ𩟑��CE�9�t���4��&�"�O��(v B8V�t4@奖�~�h����-#  )���V[`���� �O�ib4�ٴ0PwD�aw��h���:~�Yk�cG�/
�9q�X��)�8��-���'H@;�l���Py&D�n�8X�g�2D1r����+�M���@����b��F�S���@eN,���rFe��]2t�wh��,������8D��9B+�J�ǈ��P)����LU�&����)�t�l�X5"(J�L�g�'��b�銺h�.M��W'Z��l ӓh��dh��S,UV. "��	m�d1	�g.f�#!b-$��%��א&u��	�Zy��L�lT���-Q�~7�%����&|2聡!T�.��9���
9�a�/���U�q��L�r�ό�Ԓ�"O�a#�Q�T��abQ�(�D��'���5)�%�0�؂��~��>E�vj���yG�ݱ~\q0���e�4�h�,ظΐxR,�/.`I�Ql*.W,�8� W�^7N��W6�ֹ�҅��b]�+$taG{R�w+nTHz$c 
TH �u��ذ<���F�� �Ԡ����K�}�Q#��:0�D�#u�-�n���4#pa~Bh�;_f�*'L�&FU�)�U�K$��L��03v+הN��Q�C�Y�a���
���S s@�+�H�%ZD8�)��<X�C䉂. ���M�:;n�b@��*wư�2G�� �����(6R�"��:�3�$��mͦ9����H���E'�6�!�$[r�? J<��S(5�|1� �{Ja�b�!z*����p>�V�T�NX��PfG�<fE����i�KX�<a�N7z˄�C��V?qw HY �ċ��̸:��ԑ@�E�<�sm��V�@���;��� �AF�;���(��A�?֑?�b���i���{��؊M�`��3J/D�p`,U�5Lz���B�m ���'<���-����&>�X���a��&q��aC�ƶ}^��ȓg�����V��Թ��f�u��l#l�JaN	-/��@I�W)��%�ȓF�� �!���^�x9��ˈ,�~���1� (K���d��ظ@g3	���ȓ0r�8��9<�^�@��H�Q����#R爭h7�8�Ȗ^�t�ȓA�h[޻E�>�rA�մ&�\,�� 'x#sFZ%��Qb�-̳]J�=��L�8ܨ�m��q,�1
Ƣ�>�U��%�rt�HE�xY�I� +�.\�ȓm�6�ړ�`hpL��Xu���� $,s�]�A@��Ѵ{^2��ȓ/����kU'z�X=��Iֱ@h���w-n�bѡ�t��x�f� 
ۂĆȓh��*%���jV�	��A�J�}��~�=�Ek��.�$ �%�9PՐ�ȓ�B��"
P�y�U+����[�&=��.nD������X����;���Y]b�q���	6F����֘)�ȓX�.4�(0K���҄��
#*=�ȓq>��JQN��	���0ҏS�>)���3*8�"���%��m.m&���F%����F�
L���x3���NU�1�ȓ gΝBB��)���(r��D7�ȓ!W��B��#?T����H�L܇ȓ	<��y�]���
�B,Ն�>�0"
��4@�&@�l�ȓ.֐e���A.b�6	>J-���*\�Q�C�%/rhqq�L`��h�\���[�Ҁ�oB�
0��w���a�R;�ѳ��ȥdN@�ȓ��i��٩VeN"��ݮ*l$����LBVF̟yD
�� `<B ���ȓw�������>gb��� o���r�<�2���7ެ��'e��j�p$Gm�<�fJq�0�J�(��Y���\�<��S'j3��1!�ri�y�����I� I�ƣL̽Rߓv��Z0��
2&�����)��ff���ğ\"`ƭ��i�����|�%9��Q�����Z:����g�t���L��mzj�I��[�K�D-�ȓ~���c�M�7%򹘂 3�ؐ��8�DI�B��8�`E��±a8`��ȓ\)�� �ƛ=l�v��GhA,-"�̆��xL�*ϹX�����(RYf��ȓ:{cl�� ��Ŭf�p|��gA�(�U���Atj@�DS4}	�A��}r|�cG�X����ڱc��(w긄ȓ|Nt4 5���J	b�i����U�܇��l����O�T��b�m�Խ�ȓDL�m)��	�q{�E1�,��j���ȓJ%Q�'喉�F�P��\���q�ȓn\l�rI%>�(#
G�E[� �ȓ%mh�A�V+	���p�o�h�\�ȓNx�$�敲p������Ll3������E��	��H ,��CF��ȓea��Ek
�RNFq�0
P�u�Jԇ�S�? ʙj�F�o�hIcKp]#g"O�!� I�J "ԣvfJj�j}�"O�\�GP��Z�{���%=��� ""O*x{$2X�&�2�a�(���"O�@	�D�� �e��ْZS�%��"O^+tiJ�\^�j�n��:L �8"O��)u��-!�MY�M�"q�����"O�����ުl�̰���U��	Xs"O��PQ��.\�6��2���,e�"ON �	$[s�`K7o@-L"J���"Oz��.��X�vN�1o9��]�<�w$_���Yj����=��0V�<a�C:=���`(�
P.`h��G�<�2ꇣaИ�P�K��z"`SE�<�CΏhj��1�n������K�<�E�7b�x�*�Ǖ�4�j���G�<�%	@��:�#�,�p���E�<is�*M'��`�Z�{������<���3kN�PwD�;bT��B��z�<!��	t8��j�l̴(@�:5g�w�<y��0T����%.�����Kt�<	�hÒC��E��\1��p��L�r�<a&-�m�*���4(�j<ZWj�w�<1������5��#@���x�<�OU�Z�V��!D� )��ٰx�<!Q&�"y���k��
̙��o�H�<A���-0����Oӈr5��C�~�<I��S�u�x���z͠ �Sy�<�"�G4�`���އWp���Xv�<a�-ϭ<�UG<5P>]`pn�H�<!�吺qè�Ҵ*�9-��0��L�<�Я�!>)P����/ &|\�6��@�<aa��H:S`㙢i$J�J%lW�<�v�C9"G��A����`�"��桀y�<�c�:j4���yR|:���P~��#�0>�#)G7qD4���҅z�Ir��v�����jZܟ�V �L�d�éD�`pkg:D���ը>M� I�p���J#��
����)��}$2m����:^�`�o*!�̦b�����HW�c ���'�[�h�d^��d�"~J�	
�0��ι/���rhZ�y�%�_���AG-E�>�4�J�(���[�u0���	b��`x���1.h�X�gʠ �a~�eQ�HGR�Ǭ#t���a��/��a����yr�C�tFX��H�O����i#��O*$��ӭg<� ���M�z�0Hgɾv�B�	���Q�$m�1e��Q�@B�	�-@������r�|�򈚲2��B�	�"B�C��M�����ؑ`N�B�ɀT� i�q�^�hnH�qD�2~�B�I�Q��x@
G�_���� oN�l�B�<(p
��¯ֈU$�P��!t�C�#z_�89fm�(o���J()�B�I�|�dh�@.R$@�w�G
N�����FJ���I�o��0�o�"-�8 3ӣ^0|B䉝o�UB���i*�y����vH��=9���r��Q�[�ys2$�A!Sqp�)"�"OSeC`q��	��f| �u�ij�A� �T�\�c�_�"~n�}��}+��QO�0Z��{��B䉛|�D�� H�.	J)���Y>T�ΓoB�X���
��@�-�[�'�^���d�Uk��|0����X��!F�Ɠ7ި��(��v�)�����n���8 L�yh��'W\��ǩ�p�b=3�cE�s�`�;��N��ܤ����#�<0՟�$��dM  숉sH��뚨�y
� ���&��T�,���%���	�,����K���/`nPAAv�"~�I4S�eI�hSKX�U8S�ݵ<�C�1e��!P��b] `Q"j^;p��	)b��+�	&Ebf� Ab"O� ��M�N�֝pu����،"��'n����L	�1�^B"-�0!�D-�1h[I��ZE� @h��D,��q!��F�,+�m"dt^�b�*�	�~�@�T˝&ؚ(�v��Fܧ~�b
.3�&�)� �Q�$�ȓ2��9��^������ր@��*ń�\.hd�6��!
^��Q��~�J�D�n�BQÙ�}Ha�"��?�yc�2G<�{�(C�pR6d٢��<����'�2���-�&��<�߶]Z��$�ӄO�����a8�����G�6D����a4oXq��I�Nڼ=Z�fN�=hVC�	0LvL�cf�.c��"e�56ʞ"=Q�(F��}�O�(D	W+X�@���ru�'R����'\��9��©d�iH6��Hq����'ި�yF���YR�{��W�;E���N��C��$5]��:�-CVD��TnљB3C�I�l�r������9Q�,HŠ��-�C�5V���ʗ�M�59��s��N�BΰB�ɗ=�(�2�Y%��k�kL�E��B�	fD�)�3� (
�:�J-e��C�	bL�݈�(n%�#�f�ڐ�R��Oh<�C�X9-� p�dDV�yo�1S�Z�H����d��(Za��U�T�$�;1n�@0��ȓ5G}�u ��ֱ����m�,�'/ʍ#���S�d���Eb��P[�9�A��3"7(C�I�$<��!V�yEte��L�	��c�D���M[x�8�*�eT�1����a�h�@t8�,x*�0<l�	���K�
!0� *I����ƓA���@:40������u��ȓ\�dA����V*�����I�l�:���Mt��ZC��0q"	�F Jf��ȓe9�M�ad�f� ٴ��h���ɤY`S��ٰ�M�fMǦHw��:�ℒP��{B��p�<�È���"	I�/@>��dIe�'1��d�3;z#}��gSm� 'ɔ�(�҉�f&�[�<iPa�8r�nq)@�F$��5��G��֭c���������ە'�F���̼kSL�:V+�'�!��O�~��؉�k�$��4�jחF��č�L�v�2OLq؞H!�߀o�<�ɓ�10�z�r��7�O��iV˔�C�4�l��[��!��I4' ��u#˯u�B�P*�#��	���BqΈ~X�"<C
)�tr��Ә!X�L�Ș%q|rᓭ�W�B�6�<q��?'{:�H��#��H����'��3J<E��'q� �#��+ 6�S�/@M��
�'�������7Vn��#iZ2L��`ʙ'x(8��?����� �:��!1u�ԐTP0Ȁ�( '{"�|�w��O�ß J�N���R%h!i�61LY[��5D���U��(ul�Xp|�Ո%	(D�l��&K�94�E��M�6˨�!N&D�t"�핀�ȵɌ!rl��E�<��۾X�&%�0ˈ����Հ~�<��,�W�j��S�:�;W��^�<�����K`����%�|u�3-�\�<9'��
А��̚7"�Ę0&�CW�<����(�1��ݵm�^D�K�<9�Ė�y�*�k��BH��]1VB��4k,P��h�#+��ؙqŁ#F�R"?ぃC+>yr$*R����+�@�U�����?D��*7�I�]�E� �CK�V��C�>��.]�O�>�B"�����qd����t�2D���%�Ӑ0����R�Qwg�U1��0��&�ތ��I!d�n����S,�1pJ[>x����F���(�MK�6z�e �ꅸI"\<;�IƆ��x
� ���fBs9�pɀ�U��Vt�R��Ǧ���n�%4j�����3=M±S4�u�Fa���%�!�dwUlhIԏǘ�~�1��"A�6�8�Ň�@�h�	�^�(��Y�l�KN5wb� �l�I��4lO�mc���~�"��ZY���Z�Z�&���M���T)OhT��K�&1Kaz���	B@a2���L�<\�qoZ��'_|���I@��F�G2�'<\0r BvuJ c5�0J��,ZF�<��N���"L3r@p�:@�x2�K�	�q�Z�M#����a�� ��_.{̺]�Ï	;V}�b2D��I��̶`L�LA2��+�F�h��s�
����H���>F��/.l�		�� ��G��n��0��
��$^�u�X|�@bբ<3��`!Ɛ?B�!��<'u���u�C�N&��2'�9�!�$��y�0�+VS��x���-�
F�!�d�Z��+�̍u�6p��V�!��\�v��ѸCÝ	��Y k+w�!�6�.�����n��)ɟ6�!��|�&���Ԡ|�`�AAC�G�!�$~LlPS�%C�J�s���)L�!�d3 bлP�٫=����EJ�!!���Q:�A�䋯t	z��)S$g!�$V�/�ft
�mS�Z�3��͡XX!�D�t֖�:%L<�*�#�JY~�!��(>�H�'�Wf�\�j�)�!�Djq��[i�4�k���4�!��ьk$�8YE䒷�8�z�n&�!�DD#�,yaAʱ��@�CQU:!�I�m�ޅ��ș�jw
��@�ת0!�$�%OX䉡0�>e�v8�F*��	!�yh`�u��y������̘wgPB�	��Ș�I�N0�q"�)`�:B�I�d&,�#o<�����@��PC䉟�AC��%Kʐ�1ӅӏW�*C�I�.�:x@����Zm��K^�r�C�-m�bP��� (Dta[�n]�ZuC��,p�Dzv �%��Ӣ�/��B������ۃ'�����*o��C�	 U�mb�ʟ=.�2��(�#�$C�	�b���Xl�V.A9�,�C䉔����(W��A���R���B�	6Fk�����v��m(�A�H��B�%G�Y�a�
$�X�yp�I�B�I
[��Cl�A�m��iٖ_��C�IZ$�	c悱2 ���`x�)Z�'ɪpoP T�� q����_�X��'��%�dn؏"{����ķH5�M��'7�ZOܘk��%�dEN/��!�'���Rh˟x
Z5yׯݷ!���'��D8��J6�^t�aA0b ��'�:��"��A��8k!A�o�x9�'���q�I9����h��y��T��'ѢYSA�Kܵpg�Ms�p��
�'uX�YrJ� zG�	�'�ܣ8�Q+�'�� R��e|T2�6H��P�'��u���H��1i�c�'��I��'�4�T&�7��Y�o�D��'�d-�a�L/^�X�R3N��t-	�'��Y*R+R>>Y�A3>�$Y��'�ƤK�Qr 5�G��5F�5�
�'>]�#��/�.�����,]�6��'�FQ ��#���䘪S��H��'��E���?����M@Gې��	�'� q�iC�H٘���ዸ>�.�)	�'1ZD���K�CW��*� Ǖ)p������ VD�� e������><�a�"O��G#�)p��ha�$N9&�x�"Obt��N�9E���0D"^`""O�@����Q"t C�w�(�"O�lR���K�Q��OS=P��2*O��`aW�(�×�s}Bu��'If�k�nˤ/T8U��Ț�o`0E��'{�h�wS	E�E��@͕3Y��	�'�P�����
x������'�H�a	�'���z��Cc�>��T`߮�Ν��'�m�׎Y���4I{���'�($��]t���y����>jJ���'�<)c���*zh�p���ny�$y�'���sI�Z�2�.e�,��	�'2F Y����!{ć(a�4��	�'x��CÊ0U�L��n��%��'h��/YO��0��U�l$�'��p�c�R&��(�n��&���'1� `(I5j<���C�nb��'�q������bN�\�{�'-�DzQ�X�A��}���+\�n���'��!�"ƈ*�D���OS3 �����'�ЛA� �9��ɳ�H�aD��@�'^d��+���L	V�"���'Ji�m� <��p�B�<I7iS�'@�(ۢQq�q�Q$��F��X��'�!�˃0mk4U�WhT-<����'�"�H2 M�Ln�Hw/>:/R��'����
�m	�ٶč�ϒeh�'�p���*&�&���`A����	�'r�|T���>�l(z ΍7�u�
�'���pL��R�:4q�T��C
�'t�P�W΃�B9(�a�jT*�H}��'�y9 ��O�ި.�! R�M��y�B#�Mʶ�ɠJz`��U��y�ӵ���`$g߷|ˀ�b郟�yB�����C�˪v���
�<�yR��2xU�
3�V�9�^m��˟��y�(M�V�^k�Û�fL���'�yB�M9]U�|!���4�`]PWJ�y"�W3�p�u��.�I o҇�yBI��m�@����#�إۀ�ʨ�y,�(�
M���Y��V��aP�y���t��*��̕�^�X6��&�y�����As�$���i�U�%�yr��cj�QED�(}�`��ƥ�yү I� �;!��n�4@��y"�E>�$H�Rnѿr���a���y"m�$ހ���L�n����p�M�yr�ߕ%�v��" �2]�5{��@$�y�@b{ ���&v�����yҍ� �����N�R�O�H-���]F��rMآg��%���-�ޝ��K���z3�#<���+��u��}�ȓx�m�t䙥^;���b��l����~IP�
V/ɢ)���Q�Y���ȓx ��:E���1����'�|��%��`��8G�Ǝ|�	�a�4e�	��$A��F�ܫ)dx��Ȇ6.��ȅ��XH�r�C/Zb���!�T�C�|<�ȓkv��KȦN�e��&��ȓ2r��Kp�M`�v|�&ᑈ:,t��}�t���5+t@��&�zB4q��=�`�P�"q"�R���|_lB�)� x8�ԃ�<M�.=�b���50a�''�DK�}��	6oЍPa�� �u!�Q�>j�Ȩ2\�|��5!���喁B����VT�jVX��!�d_�f��U�_T�����Ԯ�!��P����5j���!K��~�!�&I"`<� @�4R� 4/�!i!��Ֆ��փЁ_G��آ��#F!�D�#Xh�����5�(@"S�țH�!��{��P��C��D6�P��"O�E��3|Rrd� ~44X�"O8���5d��	y�Q�Yx�Y"O�ə�H��	�s �.��,�V"O���s$�
#0fCwES���a �"OV��u�G7Y�b����P�7���7"O����%�&x@rL+��V�,��X�"O�P��ÂM��8����,�`!�f"O��PG�X[r�A�A ��q�"O¡�G�@�|�Q�Q���t��p�B"O�P%g��~�`�*��$���3v"O�Ia�
�P��L��O�X�\i�A"O.���mCl,B �U8`axl�G"Ot��vA�'n����b��u&�D��"O>�DK�G���d�=jnUR�"O6���S9�$�['���>�4��"O�
�R(��!`�����E�!�$Mc�ܗ*m����׌̃l��`�'�P�3a�J�:%Zy3Fn�&o����'u�1��n&+ L���?7k�'TL�YoJ+
�Z���)���@�'K���A"h����(�h�0I[�'��!,�Jm�!�^����,D���BNY��Q��B��	�,|a�O D���`^*_�|#��F�V�Ju ��?D�82� ��\$Q*b�ɻy��q��M=D����b��,\t�#�`�����<D�4�H��3����&:��]�:D�d����&�n�*fcC�[Rl��-D��b�[�l����j�-��s%l-D�\`�y@�4����6|]<��2l,D��r�݆#��h��(~��(R�e>D�(H�O�~Δ�[3��J<�0HĦ:D�( F���E�9f|x�	-D��p��{����h	l\0Q*D����gD�r{R���OȔ_�����=D�` QJ�,��p���Ə_OؑA��;D��K��܍n`0ä���!�����7D�����~�Ju�֍n4n��ԫ"D�|zU�Y&�N)@�֦#�b�2� D�(�BG�Y �;�Ӷ}�t\��k D�(�5�xAz�AR42��:��+D�X���
�pV��� �e���0T�+D�(8�⋤1l�i����+ �����*O����oL*�}��9z'֌i�"O�!b�:@�L3&ّ[���("Or80�	����s�� ��(��"O�1��U�S�P�B���,�d=�D"O�HvY/{{p�3��)$iQa�"O��فL�
��y�� a"O�T����0��]S&׍Wӂ�j�"O0�p��F�1����ƞ�ĚI0"O��F�ق	��H��e��c���T"O�z��%& �16�_&[\���"O���M�� V	S��=�b"O� F���$��W;8z���9?�0�#r"O~��dL����ɧn݇j�t�Ҷ"O��[(��������Řq.	�"O`邒���fD������u��i"O�����v���C��rL��"O̱JB��i$�sgN%S�ą�W"O��G�"\kGX;(����"O�I����2v������=w��A"OR	�R�@��I�aȠN�\5	�"O��Q�
+�x쁢/�c{�e
"OzT�!�	p�^����\�?P`tI�"O��apdHu�#хL�Q��"O�9�K�0Vc:�s���\�t�"O�����r~<���7Vp�a
d"O�P�@���d0�E�f\a��"O*Ia���-&�� b�!���w"O��7�ߋF�!8��\).�̈0�"On�S��Rq>`ڦn�:�1K6"O��rj�d�X��lʟ18�Z$"O6P
�-�J���!��ɤ%4�	��"OZ j '�l���	�u����q"O�|4��v�J�瓔C�"Y"�"O0 S�͘ ��b6���s"O8G��]����s�M�&�8"O:�h�L�6:��aš ����"O�xK��-(��P&f��Xs�A×"O�L�w���L�`xc6NX�PUj`��"Of�ӵb�[�tA�T,�(	��0bB"O�嫥�_�������ŉ.!�!��		���8bcڷ�h�T��1"!�[0z1��ʳΐ6@ P�����B!�ٴn�BE�"j!�!`$�A�!�d]�Y&b�!�(�>	bE36���!�,4l|)��΂z��D�#cE�!�D�[�h	��-�f�ȉ����'�!�dBz���	7K�>p�phk+h�!�dώ����d�$aj�u��$A�<�!�$�z�����,�Y���N�Py"')%���h&b�)]md4c�P��y"��mVb�!E�K�I4
���啲�y���j��0*�lL?�L��Fˁ��yb���\v���%�%E B��K��y��]�]�n�r��Ik��;&&��y�žv�^=p&�JD�4����L��y�=gȵA�Kޤk*8I���&�yr�Ζq0U�`	]K�P�B���y��8����2�h�@���(3�y�ҍy��B��W
�Qr��K#�y�(I7`Y�Go�P����0�̶�y���NK$�"�a�25u(@K ,��y�JW=H�\	@��Ͼ,6���2(H�yrE8>�p訑%�2�i�qD	�y�� �o���K�OA�9�0�*+�yr��,��H�v�J�5N��g����yBѨ'�6Lk��Z���X�n�5�yB�AV�2ɂ�/]�Y���l��y2M� ``�h:�	���Ь��`V
�y�m�NJ��㫕�F�S�$��y2��?6�|b:.�aC�y�'Y2T��sC���H�*�E��y"��Z@��A��m��A���y���gy.��l�!;]H�	 �y�BT阝�B9Hք�DfĜ�yB�:I�I��Λ�G�ȕiW�D+�y
� ��S�JF�!)�Ѫa
�#�h��t"O&8C%ҭ'���{ei�O����a"O>��pA�%A� H����#@�v]`"O����]�B��I"�W�\����"O���n�=bF��!�%�#E��� t*O�2� ��K�0�*��9br=H�'i���D�V�Fw4<
r�O	i-���'����pDQʅ�˨0��+�y���*,��4�F з�f��GȚ�y�ťg�>�{���w}�x"��Q�y���@���u�ϏY8���@���ybD��n䰱�X�[�z����/�yi��g� e���(\�� ���ա�y�J0�L�� ��=<Nlh����y¦A��e%�-v��bɼ�yb��7 p�IV��(R>����yBm0
��تW�F��BQ���y��� �)�G�&����D7�y��S�7��:�*ǃ/m�sB���y"��fc�L���݆*��!"E��y��ܶ4���Q3C�,*����I��y�J�dP\-�#f]�s{p#F@ �y��
�u'��sgir�!�\��y��װ^�	eX17EJx̙�y�*�g@r�
�$C2X�
	㥋��yr-��3�X�+��[�G^|@5m��ybD� d4<�an�72�l��&Գ�y��D�� �$�R&�oc����'�n���M�6S�LPw�A����
�'�
!SR�B	?j1\	uF��'�����E�/O��Tf;�"(�ʓY��9�̀�,�*U2��P�=3"��ȓ�90��8RP�Yg �?h�N���DīG�Ղ55�|�gKX<����ȓ1(��ek7v�)�NS�_�8ل�(t��3צ"�x�I�i :m���1G�Taw�$_��5QU9ZT���x��$ڣ+t<E��I@�N��مȓ{�)["�:�He;So�'w��T��F�R=�� ��OvA�Cf�IA`M��j9�)J6�Z�\O�@E獬sk��ȓ)7����疹 �$(��A�0=<��{�:����ϩ �y���R�4q�ԇ�-[h�"�n�:#n�qc�ҟo�6�����=A�fĆT\��LO�v̈́ȓES�`c� p�> zt����D�ȓ	�@�3e⇑q������ռt38y��*C���q�Z�B@�3D�N�"	��x,-J�@��o�#�!�8���ȓeI,I�ƅ
;^��I"�ӟx�zH�ȓ2j̫��D�#<̤ao�nav��ʓ!/:q���*wY�h@�c؁GxjB䉭wr�k��"h{nl2&!�*
B䉅"�t�.֒0}�d�	 ��C�I�hK8��v�?;����$8kC��4��M�r�O$5�j]�1�Ȁp��B��-46d�3��.l��P��G�B�	�==���w�͓$� �X��W�C�IW���M+
��%Q�([��B䉜=�İZ�eBn�~�ڀ����B�Ƀ4Rr��4,�v|&�Y�� C��<X���j��'v��"B��|Q!�d�S��Tд��4pA2AA8!��O�ȴ-h�j��{�\�W��?8 !�� @�3�IO�[A�u�s�L� �0�U"O����� �vT�K��fŶ5J�"O��ɀ�6vl���i�@�<�I�"O�p��f2,f�f���w��!�"O��p5a0j?��(�?v���k@"O
�{�Ȁ�ܨ���B�J��`""Oڬ���H�%9�����PI���Ǟ>����A�g�^H*����7���@�c�/0��O~�=��|�a¯��������!'j�a4"OI�P-;4rp�K�d�6��""O�XZ�B�X y����c(=J7"Onp	��� 4Z�1�"�"O���ǁ�~�]�!f8=î�b�"O��J�,�`ؑ�e�*U�R5�V"O�qR��U��#��5��E�$"O�@����%,��m`���<����'"O 2���,���ܹ̺E8�"O
�bC@Q�J0�`m�0
�`�;�"O���1����,zQ�ú|�(7"O�Xc7ŗN`����,Ϭ+X�w"O�U*T"�>|�V|ᤋ��&D� �"O�5r��T%^���#��̣#��S5"O�89�c�(.b�(�d�X$3���J�"O()����56AZA	N�`"O���¡�?;&ERPO�~�h�c7"O�5A�[V�P���Uz���"O0�î�2)�dRP	p�ӗ"O��4�/-��SC�ݑcUzS"O�i��jĒe��%r��()�y�"O&��ä	4ݜe�1C\;I@D���"O���­�0T"Ɖ����w8,�bq"O�\�s㗑��"�F^�d��d��"O�)S���Daab+��ˊ��"OtuhC-�	������=��{"O"8'o�4z��Y��j��2d��"O��VBH�*� �����"O����� u�R��p�t����'"O~]�`�߶6 i�� ^0�1�"Oʐ����=@�u�H�)A��RE"Oȉ��.�*�*�۳u(��C��'Aw� ����$���t,= M�C�ɦʖ=��e� *`�`WM�.�C䉑�t�(�@Lly��bƻ8q���d�>YtȚk��T�2�C��\�2e��<�$�km�@�`�XEe��#��A�<q���V\���l˥e�F�S,�z�<I�	gN��2!��M����E��r�<aPh�Iz�2��Ł����nr�<т�M��y+�R�K~�1���Cj�<����>՞��RKؠ)�(D��*Vf�<YF�ΕL��p�c�^�F��Ad�<!k�.g��8�U��hS��R1H�f�<�ц��5+�U��֒p�b��W�e�<A�g_�B�<��͙=<N!I��d�<!r�Y� 5-C�!�: i�B��]�<I���\G�7�L91��dkEC�y�eV�{{�� ���$��5�s�6�y��Y�Y�vE���b|3kؚ�y��P:�̘7�P����R���>��O~��b��s���b�U�`x���"O���"��@D�����7YVp�BT"O��!�eK �
�Ӛ9,�"O&�s��%N�x���i�6���"Op5���g!�����/ `�`"O� Xq
�$��X�ThY��9R�:�aT"O!dƄD�|�&��"�"OP����	��t�[ �w����"O��`'�	��Bf%N�#���#"O-�v�8�`!H�AX;r¹�"O |��l��(�q�L�;H�4c�"O>}�GMY�~�*]��GֽZFnh�$"O�!�gG%hs��Yc�Ԉh;2��"O��7��~:r�(  �{2Z0BU"O2�g�tؚ����"|���"On��N\A\�Ȓ�`�	�E`"O4ٵ��\��@��Z����R�'��)&�HJc��\�.�ucFl@�($D��SW��dѢ}ô��o��+E� b��<�O{��ЀgOL]@�p�#�"W48$��'���@���)3͈�ە�G"V�Z�C�/�S��?�t͗�`�,-�`�ޒ]��Pj�C�<�"
R���g�*(���Lx�<��L�m�@"�S/j�r2E�Gq�<1խ05i��z��X?s�|�yᩔW�<!��Zqݺ��!�7nr��qAGR�<	�@�<o'6�p*DP��@��SR�<!�F�$��=k�!�a�x��M�<��ǄW�b]9�o[i`�����F�<�����`���TmL5��EL�<YP�
7U������}�N�U�WE�<Q��K!&Ёf�ܷx|�'EK�<! �S�W4dd2�L���Ͳ��En�<14 L3f��s����l��-i��Uj�<���Pe��0A�@)0��� �L�<!P@�/IVe+���1w�EF�<��],1Ƣ9ۗ�
�:�lZ�C�<��o�\�6��-�+"�x��!{�<��Τ(�h��j��&��9 �@x�<�G��O��"beKQ�0q�O�<�,Ŧ&�rQۇ_*i��	A@�C�<9�#R��Z�[�f���Q$�\'�y�l�=}"T@a#��-ݶ��6�Z�yb�
�u��L�d��h�Ʈ���yr'�0r�~03��OE~�8�霾�ybƀ4.�bQ !��U�hu� B���y�%PT�D�p�ۦ�qI+	�y2�Ml���w��!
Į-bpD8�y�j�m�@�X�P�@T�2F��y�k��m`����2��EZ�R��y2�	+g���@v��
��A4���yBkK�J1���������]*�y"H�5����X������y�O�����˴8͞0{���6�y��@-vb�UO�#2|���n��y�gA)yئ�SE�6j�:�������y� 
���(�hW�8�8��%I���yb��3k���n�
1`�4�L<�yR+ �sPL2|�r���y��	w��`� Ӻ�h8��T��y�,��^^(��R��ŨcK��y�j� �x	��"��<�m��� �y2��]�LY�`�G�n$��G����yBd˲����Ph/m�VT�7d׊�yƣW���ɓg��*8��I�y���:m�Dm�5�B m��aFF��y�ϓ\Hl�:(�/���2�C��yb��?�[s.�����ª�y���崡K�&�� p$���D[,�y
� �� 4*WTM Hƭ�0�$"OjU��,�N��`p�S�9g���"O�l�uo���
��Dc�?U��x"O�D��#�6zCP�;ޤ=2��"O��I���ίX&
�A�"O��(���J/:����2m
]q�"O앒`˛�<��Pxʌ���"O&]���P�	�P�q��k9v(��"O��z� .J��(U(G���e"O������8r͉i��'��pa"O
��u`�JL����[;aT���"O��hϞQ�\=Zd��
<La�"O�Y V�R�S��p���U��Z�"O����"�M(X����9����W"Of�����M�S�@ 0�5Q%"O��)ׁY������ڱy�<���"OnE!,߭
"XA!��ʒB�ؘ�yR�m��1�W�s��q��畜�y��]�H�ڱ呖]Y�\����y$�Wmf� r�>!/j]%bX��y��U��:W"!A´ӃhA��y«K�'�(��E� 1��83�B8�yb%C�*��5q�E��x�v�GP�y���<���[QZ<`z���]��yr��MǸ,k��9n�����i�<�y"J�cB��i٢�:�O��y�DˊaΤ�!��N�9�K�0�yR�+3^�ԛ��^�(lx�º�y�I�*�<��f��\X�+�E��y"�U�hR�;��ÉTҼ���+��yr�Jg��S��KlRyȣ�0�y��Y i��(���W������y�C�%! ��qĐ CI$�f �!�y�!)�ޝ��� ����+L��yr C#k��QaAB	�v��p ����yJ� �8�o��f/�aV#Ր�yƞ+����T(��1���O��yB��
.���݉!�d����ߒ�y�愋vȾ��fL	�Ⱥt&��y���2�D%�7�rt+N'�y�I?.H`�'�­���A��y�ϋ��	���o��۵ K��y�Ƌ���zP�E	���ar��"�y�4-YLq���N>��`\2�y�˟g�Z`ɗ�F�F�J��"�yrL�n4��"�B,o��0a4l��y��nv��C�eM� l��C�
��y�I��[D �0Cӆ�t��@V��y"�͙��GI������(��yX0+BuaW�J8$�p��V ��y�U�(BR�q�f��&lܨ�y�	 �3_L��dL�&a�@Q�%ϓ/�y2m�3
�HQ��	U��X�6l?�y�ê�2�1х��If�	ض'N%�y��ѷ$4��j:*~�#��yRc]/4C� sdՕ˪q#R�X��ym�,08�Cu��2��*6���y'�8lT)3q�Q�ta�qv%���y�CH:�4)RqEΏ!�Xd��a�)�yr�
Q�m��B׷�с)U��yE�6���Y��K����O͌�y��)/�j������ l�yr=n��]
W	�YC�$K@�U��y�!PI��I���S`:�ŊX��y
� LШ��4�m��F���5(f"Ol�*�@N+GT@bǦ�,u��Ӕ"O����D�4��Is�C_,,s�sV"O 0���0":P�K���[��8�"Od�kB���[�GR<ST��J"O��B�(��"��܀Q�Q�X_.\ʡ"O��`��R�2�dā�+^S��s "O}�E-އ�, S%D�p�P"OJ�Sթ"I.r����M�;�� 9�"ON��&�O @�!kUD�$5���[C"Oʀ��B�b6���碘�`�Y"Of!�Fo� m�8y��M&f��@p!"O(D)�� (6� �ύ"k�L(�"O(9�%���eX���nV�4j  �2"O�H(gI�I0\�!cV�:��ey�"O�4)�;JÌ���Ώk��U�U"O��K�OՀWҤ�@�(����A"On����Md{1C�fP1�"O�k!eʔY`��!�!��l��"O@h+�MN�b�A�5"����"O����F��d�T�`�~�<E��"O�)W�P<{A�͚��̱s"O�����	��*�M�sĹ��4�(�x�eA"�J$�B)�-1���T��M) 嘪W	���,�h4�ȓ[i���%A���Խj��|"��ȓZ�r�
��G���ԩ��U� $JՆȓI�a%N[�����21@b=��#߈�jQ%�0 T.q��O�=�,Ʉ�D=��8�`P�-�.���e�8���OZ���D��-mˢ���
���3a�?,��k�L�9��	��VT�]�դW�5�������.���ȓ|Ɖ`�l͹o�)����̈́ȓ����a["m�6���PǺ���7Z�@�f�*ʪy��NA�Aڜ��ȓS���S&�0��柖>����h,�*�PH�])&��2'nu�ȓiJ+�Bԓy$u�'5��h�ȓ+� �4-W�'X��ui
�5��-�ȓZB"��K�;W�<PG��7�y�ȓJ��9��bLy{��'�'22��ȓXɌ�;&i�:8�<��$U=/U Ą�558(t��\�k�Q�Z���ȓtBr��V �&�T�+m�5g�9�ȓJ�"�9�f�4`@�k����Bżȇ�5e�౔�å6/�m�/ה#���Ҳ�A�#Z&V��z�O5y"̇�]� �IW �|Y��*b:e뎀��a��,�K�D:�O��`�ȓR���恌.o�f����M �~A��oUb	 �G-<�!��o�6؈�ȓKV��vOȣ�XP�%F�\�$$��.�ށ��Q3����&¢yk 1�ȓy�LhB��+�Y�ӊߠ*D>��8���a�ѣ(��i�;�~��ȓ)���0��)}a�(ك��u�T���k��\9$��)Ԥ���YU�ņ���;�	� ������"����ȓd�X�"4�o����5���Ȕ��
S̙��Ib���Rɘ�.���hآ�ɕA�"(�2*N�\@��ȓT]0�"eeY/ �T���+$%����\/��!�*:.S���BW�9��S�? \a2�H�!+`�եE;/�p�"O�pK�/K#.�µ�Aō�+��BA"O�� V˝&�,�$�eb-��"O}s��E�F�,N�>��;$"O<�KV〸X����d�{��"O$����x��'�W~r�"O��Y�F��0����aE�_2d"O|�':��y�dF�MNp���"O�� ��|r�HA���0d}�`"OD��P<yD�i�㏈-�"O҉�2�N-���U�V-G����"O��%@'!�:E�0�F�#/V�@f"O�aja\�aڸj�o,4��"O���Fe�jlz�;a��P��h�"O6,!��	�����'�1D8�Ä"O������&hej�"(�&�<x�3"O�ث�⅓<��s��I��]I�"O<��&�>U��
E�Ҳ3{J%a�"O��Y���
��9b�;�|�A"O~�(R�h��e0K�;o�$�"O������p�9�gׁw^�AZU"Oz�)�`�qipA�Y'c��!)�"O�uз	�:���y[؉3a�E�o�!�צ|��8��Spd���[�Q�!�͂Iڴ�C#A�6~|0����V�!�$@�x��bs�$J[`��fb
�5�!���n|�R�^�7^ʵh�L�!��Κ้ŋ	!�G��4�!�d�rZ`�oYԜ���Q�r�!�ح/��t�a�*I_6�@��<�!򤃛�$W��(��W�X�S�b��r�~$�W�D�GW�5�ƥ�	\e�ȓ~ڜa@��0[3&���W��݅ȓ1�vI	jۯ7�:�б������i� E��OD3lv4���[�zU�ȓVV��:c�ϫ"�J�R�Bي$�r��ȓk� |�pO��c��}z�U6��$�ȓ/H
U"Ga4�����ܭh0T���o$�A�@��0f(�2�ω#����hʶ-H�R?O��%Bg�Xc�؅�B����p�W,����K:]�vB��+:������$a4ř�O�#|�pB�	 F1`eLC0�����H�;ΨC�	7Z��<ٔ��%A�B�T�G�GP�B䉫�l�)��^[D��BB�M{�C�I�)d�&e*�,R�a
�i��C�	
$t�{"CD�"\�׀�;^/@B䉶'(�y�N�A�41'ҧ'�RB䉳�0 ��^XT,��AQ}�B�ɐ<��H��҇g��]�7��&RB䉻r�t�5�ܴa�>%��&<��C��c��yzU��  �9i����b�>C���<hQ���h.R��v���PB�	R���A�ʟE�Y��bB�ɀs��h
�͙e:�0��-�C�Ir��\����	f�����.�B��*�����c�2j8���F_�^B�	�1��#@�����F�%�TB�<;p~�s�o���cs�D8&B䉠0~8e�g'/#���F�f�C��$���I�ҷ�\XA�W4=��C�	:Z�D�pa��&ߘ�x6n�>��C�I'0oPM�G�FUO�!��/��X~B�	G�~d�7JTm)�(�� ,(�|B�)� &�qDo��$E�U�c�T�wE�Tj�"O (�� �@�p�b�
9V� "OE�Lv�~\�R�V.�U	�"O�@X H�?���
ƠVE��L�0"O`�K�b�-{��R��
�$��)��',�Od��B���o���M^�I�dpQ "O� K6��'#d��+��ɞ�6	�'"O̠yhG<-�(��M�`
<i3�"O�ݳ%D�3v�!àF�hPJ Ip"O�!:D��N����MΒs�tm��"Oމ��=�JX���0�`�U"OjLQ�T:q�`X��
��OC��"O����aTlF��6��2B
;�"O�TP��E�myfL��J���;"O����D�g�d����	����5D�h�ǈ%?n2��F��4!~���2D��r���L��`�C.]�!�5��A/D��ˆ�ǁF0ԝ8����.@�s�1D����}If!��Z�M�،)Q�/D�t�U�#����3GԤ����Eo/D��[���*4�Z	 �źfuV(i�%/D�L��S޾��@�C\���Sv/D�L��l�BY��&�S��'8D��iq�&#�f䅧o�.��'4D�TC��}��Y�+��vt�x׍=D��;�E�vY�MB��45i��sg��s��ryʟ4�����;�'�� v�3&��C�!�$V�qr��X\@��Z��1�!�Ɔz�z�{����!*��G�	�{L!�ԊU�H3�R�,~��!�!�ƕO["��L�^��{�O�6Q�!����)�KÔr��Vo�9g+!��n��EJ�NN!4�(���̂l
!�D�#?A�iA��?R��l�l�g!���g�A�um�9(��hՂe3!��	��T#�/c!����(!�ы.l���X5,B��Rh	�]t!�DQm.L����ׇRF:�1-ΪAb!��nLRc��'$�QA�T;QP!���K�lA�
Б4�`b NC�]�!�� �R$��-�jal�K7_a�!�$M��I���EB ���lʦ4�!��:G���w�J�'�Q���'!�$�p�<h�J�5Rm3��ǐ!�!򤘭P�{�#�6+<չԋH
�!�$�7`�2�(�	�R�[PJA�;�!��߬/�m���ΩOxv�W�V�fL�:�S�O�x�rf'XS�"tEʩ9� 8�
�'�rLbB��s0��p��U\]X��
�'�nQ"�h�t�	� P�v�	�'�Ĉ
Ո�u�^]*�B�4Xs���'�i�� ̈́))|���gB��qb�'�<��F.�JY�až=�s�'��Y����/9%���u�X?°is�'��8�A�G�4�hH��J��R�	�'t8��$.e|���bsȋ�"OR��B�(�HSd�;T��)�"O��h�3�(!�FJ4��"O^�X��jU�P�Y�R�V%A.!�ڛ������)VD-���.!�P�7�(�y虻,6��W��i%ax��'��O��A���y��a �J�ʌ2�'��O�����7s�������U!���"O�)��j�?)%����F�?�]�U"O� <�z&�ɮ02n��1%S�I�"OT�A c?�:<k��VQJx��"O�0b���\i�]P4?JYB	�4"O�X"3�M��iaRC̿��@V�-�Ş(��ݺ�Cү=��a�+H�F|����9r�� ��Y"�,��#��3�C䉮1�htu�V�C�$`R#oܯwG�B������U�)>���i��B�ɴ|�(�:R&�>p���d��8��B�ɦ
�L����юѢ灇U��B��j��%�a��찤)��3�"<����?�AФH�R�V��v��O����7�"LO⟼�Tmr���AӠȿCGpL���<D����!� n�8�b�@UJ؂�:D�����P�{���E�< I��%D�6�کO(���#�&���3b�^�<)�(�0jcg[�h'���q�<Y�o̳{�ZIwl�;S|�2D�R�<Q3��6Q|9��3��Ҷ��Q�<!����^D8p���f��+OI�<�d_<,�48'"Lg�� (a�Nk�<�����!��!펏C�R��5iGk�<	�E�h�m�m�ʒ3'��DC�� �2�$cׁ{�Th�UG�2�B��o��[+�o�,�R�a�i�hC�9p�]
��ܮN
���e��w,2C�		��;5FK�	·e�J7�B�/�y[ǉ�.Ajޜ��=P�|C�@X*DP��]�T"
m�q��tUvC�I"?�����aڅhr�LYd� ^C�	�d��1J�W[�)Ec�)y�LC�-u���r�M��Uܩ�č�9��#<9ϓ%fpɢ��#';���*ƹ,�$��,LPG�ʘBt�av	�_ND�ȓ~�b��I��N�0EI�JR�FZцȓpM◂�9�� u"N���\��1�V@�te���� wo���jņȓvEp� ч!�x��	,�ʽ�ȓIp^�� l̇7��p"W�g4^��ȓ'0��R!�{��A:6Fšc�Gx��)Z�(�,HoT���n��\�=�p�Om�<�S��C�^4���υܔ�*&ng�<i@��*��U�[ބ:Q	~�<!Nܢ:R���G�0u;NZS��R�<�d$̼s�0y�H,*��pá�Q�<1A!��@tvm��L�G����,�N�<1��6�Tp������thr��R�<��Z�cPF0{U%�@��mPr�<��Ε/�Ⰲ��4�Z	�s�LW�<i�M�H^������a�eS�ɀj�<�OҤP�d��ƪh�jl9�#�o�<1�a��bܾ4��)��%6.HQ�
�o��$�'�H�@u�� �Ht�J\2p��+�'Z��h�
0�Z<hBe��h�1�'��p��LM=������?rs~���'�t)����8�Q)��ӱ_�@`��'[�8�aʲ0!��K��l=}3q�<D��¤�k���@�Bw��}�0�-D��s�gS�{ì����N�ڀ馅1��hO���l�� A��[ p������n{�C�IH%\<�`�I Z@5��5N@B䉁f����)�5H��T��\�4B�I�o�$M	�鄩jv��AT�[�N1�C�	.:� UX�̡MX�(�EY
��C�)�  XZ�b�j��`
��1|���"O���oM�(�)#g� D(S��Q�O�,��ukD'��)�e�zG����'��w��Q}|��%H�u:����'��0`X,J�6ii�o48=:�p�'��x)�PGw"��#@�5�J\�':R��Ԣ�Q_��#sE��,�f��	�'��B��E�)RII���	�<m+
�'6R�j�Ւwb\|/L�x��I���'ўb>�v��R����B�^�bD(�r��t���I� ��C�_/�ƍ�j�3�RC�Ɏ+��	S��C;V�q��M�Yk���d^���'�84��s�0��J���<��'��v6Yo�AB,8Aӎ؂�'��KއFXn ���UlP�����y2j���$Pq�E��(�!���_���M�)§��Ӏ>��-(7���/�
U�׫ ���HE{ʟ��*#萰_-|�+�L�75R����"O ��4�#�6�Q�N@���')�O��@��i;4d�P�O�B$�A�"O0�S�h�=)$Tݢ&
E�d�е�V"Oj���(ьx�t5٤HA8ʪ鱶"O.Q���[��}����"y�a"OL��	X)FԠ��fƷL�F�A"O8�Ra������|�~4z1"Ot"fB�	X���V��=ps�7�Ş	U�� ݏ&��+�9zx�ȓi�$�S4(
�h�r���%�XA�ȓD���[��Y_c#
6�E�ȓV  ��J�!��
"��e�	�ȓ:}B�ʓ΋+TC�8
���=�p�ȓ��{f�ԁol��I���u�x�ȓ72�
� O�$����Ń�GfՅȓ8 �P7 �>�� ¨<(�4�ȓ9b0�����0���ĊL�o��Ňȓz�tze�;P�X< W�� 7�FP�ȓ ���`�AH���a��I��l�ȓY�p
�e�.tW�y�A	N�0,�Gx��'9d����ZB��e�^� �Ρ��'�NL��%�*w�8;���%O��[�'�X�&U�"��X�3� E-<�C�'>��������M:g�a�'���� $�H�vn�/,��'�0��i��N���+�`G�.� �I�'8����/���Ҽ��cH�"82q�
�'�ʘ�W#�Lt��uDU!����	�'��Iբ��[_�يŬՐ�,4��'�����.W+N����� jyt$X�'/���Á2OEԽ�*�f�F��'ƒ8R�!�m�YY1��[����'0�!c�:�j]ȁ/��LPЉ�	�'��d�$AI�}&,(qa�@�=b���'x6mhfW4 ��Z�' �<��5�'
���T1R���oH�!!6=(�'� $�V���?g�Ē���fF*L�'�݋P�����$��d���'��HdC�&�T�K�$�R���',��y�K)U��!���X M�T��'n��V�S�kC��RjF2X���O��d?|Ore�SB�+��D󪀹\'x��e"O:�ٓKSp��YtHCW/4��w"O*����YJ����@�q��"O�UzU�>s����GgP�1��"O,����('i�X��ŋ�'y����"O� ��L�Gb��
� qH�ѻ�"O:������/C.�� Ȟ -\<;�"O���P,P7GL�����+h��P"O�`�e`�z�B�[e�W)0ғ�|F{���Zh6��QV��`Wz쫳cU�6�!�M6 ���������8Rc�y�!���i��tsc��8�T���D�	{�!�d�!*�DɂE��5���:!#����'ўb>��PKи3nq�� HK4[A�3���<�'�,h��26"� J X�S-NZ�<1U�/,,��s�3!�ѓ`�T�<��A�W݆QK� �z�nQK��O�<�(L�g���,�w]b�
��I�<����W��[5ÍvG��Q�^�<�P�Y�n[�@�E.��sv��<����ӵ���{g���>s4�r�
=A�B�ɝu��j���9iء��`��B�	�X�f,x�N&D�҅�Z�T��B�	�7ȑ��O�hӰ�j���'	DpB�	=$,\ !�N���wA�~��C�	:*� F��_5��@���3��B�	�/�8"��ӥHtU��j��9��B��ퟠ��A��ଃVo��J��A�#D���խ�z��U��W0\  M��"&D�4�&g�/-�a�� �+X���:D��2�%4�8їm�.�
���-D��Ԅ��h�l ���J���H��y"iD5���� ��8#�$~��
�'��9Ђ�\1
~�I#��3=P ��
�'�Dh�RЋ��L# �+b`�O�%	�`�7�
���N �1�"O A���� ��� ��B���"O�a��	��)�֩���֧*ǆ�+F"O&�P���ھ�;��,I�>���"Ov�br�G-@��(C��jB�"O�%���� .����ϋ��4@"O�ᢅ�0u�<�1p.ƒ|���3"O���i�4����K Z�*�"O�1�䨊T���ѐ(�9���JV"O,�S��?N,��$�3��e"OnH���L�u�8cǓo�Di��"O����=찊�#C�&��)�"O~�p4��1#�aMַ�X�0�"O��[��%;�3�E�4���pQ"O>]Y���R�$���0A�h���"O�A��/K�Bd���D_&Z�����"Ol�1́	c���P�F3Bx��"ObU!��߀s�rɲ�#�	o�p)�"O�}�'�)�!p���9e�]!�"ON	�	ՈwhPa4@A�G
�  �7��|���ȯ"��H9͂�dtѲ�C,6B�8��	�DUP��@#�����Y/A�B��#B2�0�ѪSQ��}�#�lB�ɑW�"���y��1)���2�RB�	�A7T<r��:�����ę�
� B�ɫZ���e��h�>`C�-�0T8PC�	�K�r���( ��Iؕi�BC���,*pL�)�D��ӎx?
y��2D�\������+� i�L��-D� @u��U�(�Æ(O�9Y�D���+D�0��/��^��݀�(ʱ@}�$*R�(�O��c"��`k�,p�Y�h�cѼ��ȓy���[�#VA�ą6�p@��E�|����	5����D]?=X��D|��'$�>� H�yv'H�F"b����{�<`�"OH����o�4I���u��iR&"ONY#s�L>m:~d�@�� �~��q"O���#��>����)X�����O��$ɸ;����
�c���r�!򄃏k&�!��Ðk�:���#�9%�!�䚏n<p;S-Z7�P��L�����6s>Y�D
gG(�E����yBH�K��#�隲aZ��I�m��y"��5�=s�Kӭa���h
1�y��2\9��{T�Y�^�����y�%���,�C8"�� &�
�y��G7iü�����'��Q���
�y��=�*d��;i�4kGƸ�y2K2%�� �̆7Y}���mޙ�y��tW����'<�L�����y�b�z����D�:��#�Ƀ���'>ўb>! G�Bz���1(��Z�ցp��=D�0!��6kne�NZ8F�`�)!�7D� ���VVpƮV��8��5D�����ǫy�4�S�T',fXhB.�O�ʓ��	
&ğ�#��ٗA\�em,���!Iz!�3�!l������YL���#���!��@���
�ҨK�>��ȓ���'��� |1J��rx ��~n�1I�H�V�<MIq� �fX ��%eI�0R��D�7
� ����<uɺ��8}��h��A6fL��	Ay"�'<����ߩ}����(0Kq�	�'��������"s@�q$Y$��y�'�ȅ��b�~�:�7o ����'#���L�"�Ղ���~9~k�'~D|��@Lzcډ����w����'|1����0|4��rF�v�j�'{R@چ#�Jt��yv�M�C�h�H��?���?AƁ�7p�0�H���"8����UC�'rў�'Z0�Ĥ�|���娄d�Ja�ȓ1����B�Z�k��
-� Ex��i>��	�S�"x i�!QtPջ�ðj��B�Iw6V��q͑�9z:q!dݏϞC�	j����g��R�����Y��C�I�4���P2���wZΈ�E&:`H�C�v5T@�l�d�h��jC䉮:i�7ߵ �P����8opz����4��P�mX6�j�dI���)�.*�O��/���3U�2D��m�%:��܄�*���H�ˆ2Xz���CdM$O�x�ȓ_@�Җ�� ଜ �bG7���������΀1+����F�t��4��e�Z�p�@ ��dc���/ly�؇�C�wS�d#`�q��Հ��
�o���qbH�[�F9]��$mĺN��T�<	���i��A�B��S�9XE��I��LZ�!�D
/D(䅲��?BT��U�51!���Y��}I�D(=̱1рl�!��G�18P2#Ι�V9|esR��jU!�P�f\� Bw���0|���EB�p�!�!��m�ቁ~fЬ��o�!�_Jl�(��-|֜�$M1}�!���+\ɪ��p#ބ8_|�%�6!�ć)pJ�����hFr03���N�!�DB!+\�H����I?��:eo�9s�!��J<uܝ����:"h1@��_ ,~!�DI-d@N}:����*H�u��O�� Hp��.�/5x�	��1w����"O*�	�,Φ:t�KW�� o�U"O`����S,Zq�GJ];���"OƸ "��-�Hx��ȩ
�?�y"�$F*D�R	���7���y�I�!��us��=X��)R'���yr�R*!�>9X��-�
��q�"�0=����6}l���4�M�zT�j�@��y���+>� ��qO���c���$ �O���#Δu�}����JOf�h"O6����v��q����_F�)�"O�v��C�d"d
�Pa� ��"O�����C�؍�F`�0oX���"O8s� {Rn���
D��ȳ�"O"(��ŷ9�=d�ͨn��`#F( ��|�����'����Q�'b�t��GC_dTI
Ó�hO�i���o���(nK�6�x-@d"O���2�V�D�\��CGW8	VH�e"O�ق��RDfᘄ��5T�u{�"O��%�.t<aw�X[��88�"Ob%�3D�s�����3pZr� "O��2Q	�H�`����RK�}ʅ�'T�O��	DƎ�vX��D55��5"O�`ș�>�*b���/&}#��"|O"yy�d$f�qC/�;t�=��"O(-���'IZ,�t�#D��y��"O��*�E@�j�T����+n�>I;7��l�'��	
9�0�B�Чh��횄�\�0	�pD{�T�8�ʄ/�v���A֮�2��iu@��<9���ӶQ
<�IqO��W�f�����C�`"<a���?��7 �Gy|����������b�!D��`��<���!�O��ԡ#	!D���ЌD"'�Z���^1��=D� �@F؊G�H+�&2uR i>���	�mb�m��Ym�����O8i�����(�I+9�i�
YzР˷kL�0nC�	�p���d���:���g	�bP��	~��xxr(;������	�0�p�W x����	;{���#�kR:`�jL��Gů&�C�ɺeoV��g�!��*Ŗ7P��B��(W�@0KDbC:r���k��S���B������˃�*�5��<v��	{����N���F\c ���Ḳ��!a0"O>��de||4�P�&ɬ�r�"O��6`L�|T�j�b� zR?O���DB"
>��"JӠD��$�����
�'>��"1b�X��@q��ܧre }�	�',f���@K��9t���V��	�'�xz��65o��ul@�JJ��'�,-h'�o����t�	��)!�'<h��A��%Pb�,\*p%�L��y��)�S�08˕�R9$�K"l�?�2��e�I_y���YV$���0�>f܍�����!�T�6"&�#38��W*��!�DZ����x��P��	gK�!���l�4}�s��	./��2��`�!�[R����v��/Q#��[U�^(�f�=E��'Ɍ-�@95-�<��M�.5>�`
�'z���R�K� �Ѝ���F.�0�K��d3<OZ$r���_,X���k6ʥ"O��ѓj�1jJ���ᘍM�2r�"O��r̞�[tL���MؙSs����	x�'~:M �Ϝz� �4㏣%u>	�'��3ǁM�I��U���ߕ ���y�y��� �Tb&	�Nl�X�!A�3$�PК�ć��P�0Z���!=F�0�� v FC��"h��O-�XA�[y�NE+�'Bb���>+�@m�$	��_ ��'��x&��/���ιd � @�'�r�8#�Z�c.���I
��!�'�����12�Z��@���8M���)��<���<q�`�R4NօrE�0Çi�R��F{b�L7.�*��Ȗ�0݀�P��6�x�'D�$xQ�C+x��%- XJ���'����M�$%�T�WQ@H��'��d�Bb�X@�$fܹҒ�I�'��jF
�/w�ȃ3��3	}�3	���xU��J�C��h qf�P*l"Vчȓ+�tX�l��LIj��Z'e߆��'�}���??kt4�Tm�R@���4�yB��R�� V*�-b+�I��bG�y�!�*+Wl� o�Tu]A�$��y���<1gDTZ�G�H�F�ϵ�y�nR���5)��-S2d���^�0>9I>	0�'��@s `-"����<�I>�
�Mм
4jGF���mН>!v���h�r��Cl�1�����O�t`��ȓvk�ȵG%Lkr/	�~����.`8���"]�D�Z�h��U;1��]ʕ:e��&��##��p؈���V��$0򏝛\$���陨����	s��UU�Wꛌ_X61KǤT�O�x��y�IXLD�3�O_���`[2a�#q���d'��(_�R8�A�z;�xYg��w���|�IE����'>�A��,_0�j�seZ�!�䀣�'MD<�	Y+ z��F�|��Z�'�H���C�W�v��D	W�El��
�'a\U�GX��i��K%U �(z
�'66�J�%t�T�b�c�4#9�M��� �S���FiN5x����.ǚ���,�y�DiJ)`S�1+�z�[�%�3��'��{�kQ�;0ܡjP�M�BM D���yR�F	sԢp�gL�y�D��)S��y��S�t��5J%�p��q����1�0>iO>�r&Œ-���8sO�6�d��B��q�<�H�	?�]{uI�3yj
�Pҋ�n̓�hO�����)uf��֮B\�Ċ5��<	�*��+��-�d��:��P𒀘n�<��%҉2���e�z�.̓��o�<1��* �`�,����A��h�<�tI�mx��cCg�|*��d�<��Ӛk ��5M�|��u1Q��b�<aЩ��ؤ0b �0��y���d�<�Sd�{�Ġ���Zc��p�����x�jѓ�N�"f����(!��yB�6�d�qG�s�x=�ߔt�!���Z�aZ4�	�%��d�sυ�e�!�D[�u\�����Al ���4|�!�''�S�K��p��h�v�9!�$��PCr�\ ej����wa~�X���T�C�2u�s��,�"�;D��)���) ���\r� ��F/��蟾���e^�� �W� ��=(R"O�8{cT	fv���a��j�j�"OH�``�3f�89��K�/1�%��"O��ف�
���Nk&��"O��4��8����'
՝iall"""OR�1t����P�I%Y�f���"O� h8E�Y��p`�=��!�"O��xP&��}R�}�R�E3��dh�"O��3�OD�5��Rc��%S�F���"O�-�CcRh�p@I���C�|�@"OJ0e)��k����Ά��8p"O��XD��V]z���õ���a�"O|ȣU�ͭQV�(�L�.ϰ)*�"O\�G	?aL
7�OeHX*�"O�j"�.U�B�A�Z2����"O�	pѤ4QOY��蚀v�TU�S"O(-�@�T4�9#��W�3�v� �"O��%��8Խ�F���*�pȀ	�'��D���@W�ܫ���S3���' �\+�	'5�Ȅ�b�	���QJ�'	,�1�����X��=B02�'��Y�SH�?x9r��q��Ezhh�
�'i, KRhl�(\ ah�+f�l�3
�'D.a��g��7�^�S@�;d�.�a	�'E��
7�*Q���b
!+)�r�'�<t�P-�.
	;��_O���'���
J99�u��fR,І�rd̜§�#ɢY2B�ɱxS(���l��<��O�U�0�"�� vF4��E�Da�o�D.H�"�!u^���D�N �A�a�Д�4���_M�x��S��=qW�_5���k�G����Fj����*Ǯ!:�(����NU�Ѕ�zl��*����C�n% ��K�ͅ�=Ɯ����\��ѻ��t����"' �3�M�	D�,i��
mD�D��\����ʀ>2u�����np>���8�^�!�S2����HR= �ȓ*��Y�F�O$&�t��c�'\�=��N�P�;�V	3���t
S%Z�>��v�����L74O�)����9T�����	�ȁ��S�k^r�瘹v�����2�����Ͽ.Ѷ��1��6���ȓu�@�� �L����'�.����)&�x����${#�t���t䄇��b4R��c��̀�S�s>�ȓ؂ThFX�4"���D�h�����{�ܣ`�HL���M &���$�0��*�UCj-�.	;Lp��?�@x���Ch��b@�J�4L����0�le�3ǄN�^U��똀y@6a�ȓ P��䃝�4��Q�$й�^T�ȓP�^]��K�+>���Q��4cT`���9�8h�c��T��)��b�,g��؇ȓ_h�L�m�[ߚ����HEg����2p`t��%K�)����
��%��1��F=��37�4$��)���΁#10��	�=cc�K�b��B!�:M�i�ȓf8
U@@���k�<�4A3����}8ȵ�b��2�A��'M�BJ�`����"0&��eJ�#ѵdC���rV��!��oi�8ZR&�o��ՇȓE����D
$H�y�Ŏ1T ��T��L��ǟ5j���!� �-c��L���>q�Θ	���%�G�q<�=�ȓ?DAD�ћT�r��� �V���W.����]�d�!+W��J�dl�ȓwgl �p)��'���R�/]�Ml}��}pE��J���V ��<����ȓuB���7�WtjZq��R+JR���S�? �)feB"TDy@!�л��1ʅ"O�(�V��dl�d�ցYh/� a�"OZ��E�:���@@�K��('"O*x��ѡJ�E/��
�d���"O,E�e��4	��{�B�\0B�"Od$���Y�b4d�����V���U"OA�D�J&a2l��)��i�"O�5@啯/��(���O:���P�"O��0 ĉ$�^9SU'�M�|P7"O�	�%o�;�J�jBGB�A~�-p�"Oh��Ӄ�^�V�i 畼3����"O��x#
T���Cf]��F��"O�z?B���0�]k^��"O����d�t�\�T�I��txJ�"O�Xӕ��S�� �5�ߩh�h��"O�<���B2u	�`9 @�F�He�3"O,�ZaдJ��!��,�&ɲ"O�R����6���0��1�0���"O���t� �$#l)�CF6�Qt"O��C"�c܂���OT86�޹��"O �*��-EwP�y�(�1*�8@q�"O*� �o�!���!���R.p"�"O0ɐG���]����
��@ʡ"O��x�Č9�`�3�>v��`W"O|hQ2H��G���������5[%"O�h�&�#Y

Q�B��6��i�"O�����C�{ t}������jL�w"ONY�,Z<O��	���P�n4~��@"O���$%]r����fN�cN��u"O��@F�V�DT��o,3��[�"O�X�Ɂ�_�l��ՌO0�{T"O�h���ƬR��x��p�	>�y���S��ŀ%ʦW�xBwgI�yb�F9x:��`�RI���c"��yr(�ppi���#=� �"&��ybNY�LG,8�iǽ_i���f˒�y�HI#@O^�*��X�mI�]� �M��y"ċO����̅hUΝ����yRd�m�|�{�l�x�����ۋ�y"� |^�TP��N:WBl"�lX?�y��Ƙ_�(���9���J�I��y�NX�~$�Q[��E&*�(ɡ�c���y2`�  �l�a𠁡$5��26J[�yRD�2T���A��jY%CO��yb/��;�(��3V�Xg� DmG?�yR �,��	'�A^<p,�sc
�yR#$��I�d�ԛT���q�B��y¨�+$�8��DN�LҜds"���y"�� 8D�S&��
Bz�������yRW��a�@�R�L�:���y�+B�tQ��"��3G0@и֠�$�y�(A�f�m)�g��:/����A�!�y��ؗV�p�I��Ո/Vޠ:��V/�yblZ�L�aqFAT�HBg�^�<ye��>��0�f]�Z9^a��k�<A�`��/1 �`� ��'��;V�Q�<�r냘��	8�"�-cqJ�O�<w�)p�j(p��G�����O�<q� ����B�`
 ="��6��H�<9B�]|��`�cK� Ә(C@��K�<�TC�Y���Y�[�4�j��I�<ٰH�I�d� G������H�Y�<��GQ!j��p3���c�H0� R�<t�Q15M|�{d,#�6�Ham\O�<� �A���� ��*G�D9Yo$� �"O��@�	C�D���V�.0Te��"OVI$�J�=�$ �gF.#8��Q"O�U@`���$����%�Z>3E{�"O>����<wLE�'Ś(p�C "O�ٲI �%�� �#�ޫXmNYqR"Op�kI�c�>��v˘g�E�F"O8�'��?)�H���	d|I�"O�Py��޴�BC�4n��u�"O���''G��a�Ί-���!�"O����1R���%#��~��`U"O"�C%�҉@Ш	�A@�S���"O���%F�.�xq�g���z�c"O�m#w�	6J��t07 H/M�0dA"O��Yҁ	$� VL�Q|���p"O�����X�71��zV��c�Q�"O�E˂����U��;
c�ș#"OtX�SLײn��Ѷҩ
V$Y07"O.0*&(D$U���!�VN�qF"O�9�����8�OF�v���JE"O��p�� C�R�r�@ˣS�ĜS�"O❰���$Z^���s�x-��"O"XS�
) ��@���{[��'"O^��2A�:Q'��QEL]Oyp"OVdB�tA�4�!��*=�E�"O�y���=?�a��
�6��H�"O�9s��q���riA^'јv"O\�{����&5���!Q�5��8'"O�`
s�÷]0bw!YZ�9"O*=��蝲�(��Q�B�%�T�"�"O6y
��ʙ���#!��ڈq�"O���%P�-�z�rGk��Z�6`s"O��C1����U�7A�9K�05��"Oz��g�T ���h&��u�d0�E"O�<�SlI�*���)�߱���r�"O^E��:&��1��k�@��"O<T҆ŶQ|�(���Ů�3q"O��Mƞ%O�u���E��p��G"O�0��O�)���6�� Q�5�"O�E��mV�4�e��-H6��Q"O���t�^%V"�A���: G�<��"O*�#��L g��TP���,��Kw"O��0�'�kD<� !U�4)SE"O�Y�4��<-���B�o�H���s"O�qC�NQ�>���R�k@�Q�,iJ�"O�p�DƑ%��(8���?ofX��"O^q��Csm���D�U)P�,s�"Oܱ[U��	n���IG]0���b"O � ��A�МYR�^ \{$"O�$��T6tI���(����"O�Y ���wP��Pl�8D���""O�����A'$�ZdQFM�;Anfšs"O�������~�4�1Ё�.lf\��""O Y�ъ����-!�� |U��"O摲E��>)�� ��C���D"O ���"�0lL�9Z�f�q��B�"O��xB&V�=�����-d��{�"O��A"휛I
�"���6E� "OU��F�XИ��зv�B$�4"O��A��^cl0�[����B��x�"O���&�;%Ά����Z��m��"O���ȟ�7�z�!@;*��Q{�"O�M�pe�	(`D���	�/��EYd"O�17'~��r����I�F$s�"O� �	�O�_M�չG�ܫN�ܡ�"OV �g�(j���l�x�� �R"OT�a��,8�KA�R�`{�"O��ƀ�V�96�ՎdD���"O~y��a��kݠ��`�<v��� �"O& W��n�2�p�e�T�b�1�"Ovx�S=���0D�2ҲQb�"Oz����2=ެ�2���b`x�5"OЈ�獺P"$pu�P�M��"O
��䟓�4i@iG?f�K�"O�wOب=�T��'VVyp�"OQɷo)nx(��i��[R�y��"O��briJ')e(�&Jh[��+�"O���a�Ĥ|����P5$��&"Oq嬓��is���j��S"O>)c!�B�|���JO����B�"O���Ő)�(��7�Șxj`{ "O�]Y7-�)( ǈ�z[�`��"O~�sp"T�U�(`*U�W}V6�i�"ON�a�ق?�-��kN�:��@""O��`-ݞ+4xc� ݆%&b�C�"O�y��	�0P6E�ůBE�P�r"O��f�A5o��j7��U;&��q"O��	6��l�tUz�M�&,$�,��"O��q��OQHE��#�� "Or�@��,f�VIB�j�/d^ZEx"OH�٧.D0mmVM��^-\Ndܻ�"O6��U��r	�)HB�Fg����t"OV,��KY�Np6���f��
�"OF(�i?7~6�a�Ȑ07E D�'"Ox�!�T�*�"wN�\�2t�v"O�m�����r�tMQSσ1��)�v"O��	��D�[1.����U�<�.�r"O:��TGI5l4��"�
�6~8$��"O�̨VDS�q�]��Ƙ3z6�1�"Ol�0�k��=�d��Y{� Q�"Ox�yg�M�\��kRD�Eu��"�"O(Xzr�۟�Hi���̎tYZLx"OLh���ݏ:�|���!�{FT��"O��#_$��DPӂ�G\b���"O�ً�˃"~�2�k���+3cJ��V"O�T��+ �(D:�ŗrIx<("O��0���:=(���nQ�JLr��B"O��/����"��ía=�`�"OVX:4���f^Q�f�ƅ(�}@�"O� ���d��'W�"+^h��"Od��S�6��#�#�.E���H"OB�
�"�<(��(ǂJ7��I)`"O�ARu�E�B�QH0t��p*@"O�1 E�y�$XX��O�G��0�"OąA��W��a{�덬J?*=:�"O8��Ca�L�p媥
�'P��Y"OdPK�	ֿ?�� �
׍Bdz�"O�y�D��*�F�P�IڡZ�h���"O��	A8U�lp�Pg�;s��pju"O�#0���% E�y����"On��j̆�FuZS�T�ߒ�"O*��aP��V��1��U"O���U!r�`m���+}�
5�7"O^�Ԯ� N ��H|��S���y �&7+��8��ڐ9����'��yRF״��(#ԫ�24��Q�R��&�y�c���p�#���0p��e�R��y��E�kq�����U�"�� %E���y
� .yk �%0p0�t"J=��H��"OT9�S�=}��BQ�V[Q�`k�"O�H��L��]� ]8<̃V"O�0ٴ�W�mVf�Ή�}�F8��"Oy�!	�^$.q���/�F�0�"O<4��C�xE�I��4T��"O�����Ͱ4Q���ː2>���"OLE��ė��8H�)E/F����'"O$��<����G�@ؠ��"OT@Pbl�'{��Q��f�'��A"O4�F�|�v�k��
��%��"O��������VCQ��&��\Jd"OΡh�b�L<��޺p�4C"O��p��Ⱦw�1��� ��t�@"O��􏋨Y��X8q��"��Q�g"O���d�k��K�N%�ڡ�"O�X�V�X��y���F$C�j)3"O��KL�mw�l�បU#�q#R"O�a���D�gM�8�#D=pQ�"O�����ZB�|+&�N0_�ƨ� "OF��L�@���q�*ó?�ڵrD"O�1Btl��h��h��kӜ-R@"Oؘb�H	{��Uʱ�� +�m�A"Oh�@ <�D��o�a���"O��1��]�$�
A3�
�]�f�@B"O&,��)�*]�ځ���C�X���CW"O��CT'M�0�2��Dӕ*c��"O��x�G�_�j�9Q��{vr=��"O��9B��>
lP|2��+Z�P:#"O��
4^_��� r-R�q"OTQj���X�s���H�R`i�<�#"��`��	{�%"�����i�<�F�5t�H�e���,��Gc�o�<y7㕸i���b$�<���GPd�<i!�5q��lpE��b�X����k�<A�,ʂS�|�	B�B�&ƞd���j�<Q��O�h�Z����"���b�<q3D��*����<g�Ę��_�<%m�/R�p݃��@
9�v�PЈ�X�<�'⇠�j]�Rh�MA�Ux�SU�<Y����#$l<�)�N�<)�mʦ-PpS�M]N�]���d�<9���bΈ����D�D
<�"�_�<ie&�$�Ѡ5L�	k��$,]�<�B/ԘX+F=A*Ū	j]��$�X�<�a��iI�t��ҩ?�x!��k|�<�'ގ 8PHJ�k�$2R.�#S�M�<�&*�j�؇�_�E1����(Sd�<�`�"O�L]%���r��̐���d�<	���mV�I�7��wĀ��"	�`�<�B��<������9t�r���_�<9CDI.���:'n�Hȩ�#jI]�<!'o�=[�de�'�Q,��0�[�<I��B�nV$����h�V��K�m�<	� ��'�����Z��P	ԡBc�<A��"N�څڅ�9	��a�a�<Ip�������+- �M��R_�<���Ҍ1�`C�F�Rה�*�C�o�<!�" ���@*�Bɿ:����b�<q�%�������9d���+&�_�<�C��;R��t���ܵ;�@h�Du�<��iܟ:��t.E/x��|xLUX�<�U�P�f��x���M+y��T�]M�<ѳi�6=����]� �HIF�<� ����Ib5&X¥O&����"O�i:5�BI(�kH�r�0K"O��y���D�u��V9sё!"O`�H��)R[����Uw�5�`"O^�9f��&N��A��o4}�"O�%Ѡ�J!{+蔑���T�8�"OP�ks�V�)�e;Ge��EV,�v"O�����5siN������k�``�"O� �tIQ�DaPt�S�N�^���"Ox��的~��ePw���<�l("O�t:�.͜:��A۲A�oÎ	@�"O9��@�5:H���O���L�`"O.1�%��~>��O���N��6"O��u�ˋ:G�)�N��X�9�*Ot�A�'���)P)�-T��D;�'�"Q���h~���2�T�`$�t��'��Z��Սn7&e�3���D�����'�򱂇���c��Mj�T�/%8,��'t����A,u�1�2C�{0Tؠ
�'n�eCJ�����B��yL�h	
�'g�1IB0H��K�yqJ�	�'F�K�OF�Q����s���	�'2Hd���	][���-g$�9�'h"}�4�ݬE�T8�ph���!��'@���-�Z�2h���ϰ-��	�'dt�j�$�>sPR)0�Ω,����'`�,���<T^�����'A2���'p.�����L������<���A�'�m1��0{R�a
٭D���'�,�g \_<����&OM��pr	�'yV�󴊁g=���!�&JA��k	�'^�i1���)8rD�s�C!;�F���'��I ���?�>Z2��@�>�"�'-���0��a��)2��5���i�'6΍0d��-p������.��Mp
�'d�Dg�/:�t�`#]��z	�'><9a�B-p�~�y ˂�t��'�P�b�\YP�����i~^$y�'3:���\8Ŷc�'ج
%Ua�'�R����:% t���Lܨn�B��'G"ݒ��<@����7!�T�!
�'�T��R5f׊�`rAM�=�hl�	�'�l�8-ڭ&`8���-��&��
�'���JPN�� _�M��L�#9�1�'p.x��K���e����XJ
�'�P�viX�<�
���G� *�!	�'�z�V�J>HH�C��>T���''4`�4M������e� H��'�tY�1�>�5p��ΰ~�r�'+���i&�%���b,��'l����Ԓ�`+�B�X� �;
�'~���!�͓.���A7ȝ~��
�'i��;" �3'$N,ʁ��
yw~��	�'��$qR�W+_�j������nH�UJ	�'�<0�ηWڢ�js�C1s�P��'�:���k�s4La��7d��	�' 䜩�`�1/]�jE��s��+�'�*)e��Φ��Ĭ��rGdp��'�,���B�#&R�- �lڄm�$d�
�'�����G
N�K�R�h��P��i�<9�l@CD��o�a4@�Z��i�<�2��KT�Uv�;\؁�iHd�<�w������ɾp �U'�\�Ii���OyF=��딇.����?������ .�w�B �Z��FfQ�k[�j��	_��x�iV����L_�p�S ��y���>?�zMQ��߷% P�:��#2�X���'�a}2+'[����� �8�"��-�y��C����!�A	z� ��+L�y�cU�dT*!�X�1�
��TI��hO�'�"%��mh�H
A�3cU��0C�	K�"��Fk�����B��Q5n�,C�Ɋ\��2d��d�d(7aq�����n���J�$Bs��@�Ȕ�9^ �'�ld��	�/	BLse햓?�>ZƉ� �^��=}� (<�eK1��10W0qs5�е�yR�[a�|�fe�1sH�r$ݔ�y�ț�ڹ�v�K(m�x�X��E�yBJ��m&����`W�x�̈��y���L� ��E�"]ٰ�
�Bۆ��>O����	^L��4�Թa0=���+D�ԋ�
� �X�go�,����
*lO�����DW?8j�8�ͤ_ʥb�)'D�K5�Qsl�i�� wQ�rp'&�	J���'�^��U������OJ9��.�p���( ;�$) �M0u�h��ē�0=� �#������v�T=.԰���Cs �sG�������@\"!�X�ȓC�X1@X����E�S�|�Fx��)Z!aŎo:�	` Q�FJ���l�<I�OH�g��Lj�ɕ=M˾a�V%�M�<i��!E���I^e���3�E�<��@4:n�-�Ԏ�".��(���F�'Hў�'TZ�4��-3'6�j��hfC䉣8�R��E"υN;��30��@��hO�>2ɷ)Ӵ���mX��hQ �2��l�l�� �! E�/&`��˒�C7O���D��OIjty����XcdU=r!��@tL���󄒪`c�����]2W!�DU
 �1���؎CF��IW�בl��OȢ=�OP��[�o�:;�L�!���(	��:�"O���M	� wکq �(1CB�9�"O��AeYp>��V�6��p[r"O��u�5^�J� �+�9QdD,��"O���O�J�i�JL�M$�qC�-�S��y�-]'O��!�'b@'8RqR�Q?�yr�P�K�"���gR�^(���@/С�y2�.�Of�7cރu~�`Hr��F�6t��'��,�O|�
0ς
Z �U�F�\���ᕟ���)�O>��`"�O���q͘�.5���W�	`�'7��� �I���2X���A��oրB�ɜ{�xСE&�T��(��֌C�ɚv��Iqai��9Ӷ�p#�	6��B�I�f3����EU*��$1V/�L؆��ľ>���ҕJ	�l��ㅵ`��|�jLL�<E��6�HM�7%7e��b�F�<��iF�:��J�
Y2���f��wx��Dx"�ʚP�i.�
Ղ������*�S�O"d*�߀�&d�튞�t K>1����S�\=�s@�Ә*��bc��2��4}�΂`yJ|&���Ԭ�Ta�$ ��C��:$�̪�˪L�D�T &.Xv@���ѕo��$�,x��ᯙ)�L�b�|�Z�����#<��&��`Q�*�!��܃=�R�(�	�;*�� BV�	&�!�$�<`0�㊋S�~̈R@�k�!�D�"e���B�]�9�8�W�^�p�!�$ԙq���Ҁ�+����MT��Bx�� l�K6B�+U"��{׎hrD�'����<� hJ� �6o�Z)1� M d B�	�Y�$��s���5�*��I@�Qj�#=AQ.2}r��̞YJ6eB"G�!�h�26�9�!�d�tx��f�+� �Z�KL�0��)�'P��g��A@��c3e8�%�
�'ar	��G�q�c�5Y?|D�N��D{����ם+�B`ƄX�Qh�N���>��O�9���O�����-a�&0)�V�D��ڰ=����G�=����P�
E��jYx���I�<�2�ƹXO���1��9)�P� ��Q�<��lU�z�IDk�5�\=�O�H�<���5�ԑG��o����,�{�<�d����5�B,��"C*ࡓU~��(�S��G�0H���T?n�Ȑ1@��L�L��9���Y���/9)����ϝ�NlX!�=	ۓ��ٓV��w�*��kI�]Xj���x t�t�F3Ʀ��6i�����hO�>�ȇFEr<U( ��-O�L���J"������;��P3�@�@��Mˡ@������v�&�J���ȴ�ޖ&��i��h�,`��'a� �Crh�(�R��"O����G�zb���MU�^�
4�"O4h�Q�Y{��l,ƗY-�T�Q�$���F�D�B�9�"�a�04d�3we�-��D?��b8�;+:S�D�Ҋ��B��+b��O��d����OnU�,��'���f��7=�\`:�}4(@��TX�ܳ"�X2c�mp�K�'0*���'�:D�� ���6n,�@�'�"i�4�:S!8D�����֠:�9{6�^�\Y��1��Y��(O�b��bǡ��4����܇N���0�O��'q�)Cv*���P����Dwf�2��)�t`����2�%ׇ\����C�\���'K�M���"}:��	aK�x�!�@j�BD�gg�<�g�O	f�HU
F�T��*$��Y}2�'����,	)  �,ɶ��
&u���
�'H���b_�eeF�!(��K�١	�'�(�� ��/����-�.�d1��'=�dI�.ˆ.����k߆r��1�'������8t�4�
���WO�@��'8���g�ə*E�`9����M���:�'}@8qP*��J�RI��9S"�@�'&�
��G 5XPcs�&z�(�'���Faԥd�t�ӥNH�8���'�8�i�W $ɤ0�b3h��q��'Ųx����+|��rS�O���i�'~(��F�
I2 l�wjK�~�M��'���Kb�6'i��kB�Ӽw��d��'�6��@ګ*IB�����)w��}��'N��ه�ӭhɖ�CZ>|�l��'Sح�W!�&z.��0u����x��'����s�4-T�7��-P�-@�'�Ԅ���	;�X�@�/luP$��'�-r1'ڞl�X����f�n��',���D�
���4D߇J���'�Z�q�m��Kv��>�-H�'�BU9�'�oc�S�� +���A�'��ذ��O�x��е�'D|E�'k�	9�C�3��hҴ�P��fԘ�'s��qB��|�%����8Ċh��'���	1�8i�]A����e+�y8�'J`� 6L뺅ؓmD�]lhe�
�'��Y�&T�k�V0VB��&����	�'9�`9҅�r�'B�,�e�	��� 4u@��T�jSj�3���Qt�"�"O ���\*Q�XC[�ud���3"O��Xe����p�� >4���R"O������U�.`�F�2 FԹd"O�р&$ީ�JUb��X���"O�pK�8g<8�篅+lL�T"O����IC5D� 1�2-� k�"OFX(4���C���D��%g��C"O� ·O�"[)��)*�xl�Q"Of)J!��HА�1I�T+�"O�(���Ƚ\ľdc��=	f�h�"OZ躒�N�)/R�Jp��Н(�"Od���V
y�P۵���S�"O����=R��(wX&�Q�"O�50c FY��Q��T�^�Ҕ`�"O��˒���;� эQ���s��^?+��!��? ��d��"L�%ҷ�)b�庆�F0$(!�[�n�LI�-��j��M���� !�D�9�ݡ@eD��M��gд^!�D�;��ce��@h�I�� �!�$ݥ!IP�u���mW�����@�	K!�dЧ�Bh���ԬDQ�b�\!�$��8!�G�<i����E�>!�$W�*��l(��@�3i�CPo($U!�DS�&�BXi�F̯TB �5�+=N!�dO�:v8z���s�rd�����!��)I��rG�L�A!TS����!�$�?gDQI�hL�g0k7���!�D٭B�<��ә8&�Ȫ*�>5�!��1o8eY�DT+xG���*�
9J!�d��j>jeh j�<*(�&H��24!򤗉�U�ь��|?"ŋ�B��~'!���3L��#��O ��2��
=�!�d(-�P#���Z��y��@i�!�DO�q�j��T�j6���8�!���\J��Q�A 2�6ܺ�ڌU�!�DU������-��tp����ю;!�dʎ,G
�U&׷xd�VG�<<!�D�+�2���懆Fd��a��b*!�=yS ���A��1&���M58!�䊚F�|Y��Y�l�	���T!�[#��e�ૃ�#� ]�a"��8�!��84�q��G|�
��RI�!�ć1uY"�����&���×.M�!�DK�Vw>@� #��C�d�1EL�<�!�$K�YҊy11
�����RA�3X�!��8�[e].k~���ҫ�\p!�ʔ,��HȤ������7z!�dϳG�5�uc�7���'#�PZ!�$�����1׉]�$���aDۉp�!��		�0�p���h�<,ä%���!�$�/.:�x��dΆb��]��d
�E�!�$�o7����	j!NMZU Q!�DM:Fh�l2���&G�X1E ]=No!�D۠@�4X�SgDv�P�xw@\�FJ!��I�֦�Q5 V+v�!�/!�G�Pef<9ӳ9~`,*�+��<!��1�%��MIQ����&�!�DI	�
��@�Ή,Y�4XF�^;}!�ĎO�@�*WN�P z4��J�H!�F�B��ӅkYDF�[�	Oj!�$.U��B��ɩ^9�"g� !�dZ+7���R�(He�,�e��i!���6*���+��LS�(j
�HZ!�� T*S$�++ [��h�Tt1�"OD�ڄgM�^�:aZ�C�G�j�{�"Oz��q�Z3W�<�ib��8v�(��"O�9�3c�-_��]� 	P)n
"O=�a�E�`���j`� ��RQ�"O4�6O��^h���؍v� ��"O���E��l��
����t%��"O,`�X�_�T���&�'Ws���"O:a["�$BA�W�>s��{u"O��㌎�$���w���[���V"O��QKi�kq!Y;iQpՃ"O����Ʌ�x��&�ZK  �D"O�Y!傲` ����+���"O���B�,Xyz��"%lPD�"O�����S	p�ң����S"O�pXf�ۃ*��6m@w���J�%�O�}s@�֞�����������U�������.D�xAb U&�f�
�qz�y֬������BV>�k��'tѻ7��l����	�������$��N}rݫ7�D�b���b�b��})�iJ [�LB�2.�Dq� ���Sw7t�Tc���m��Wϲ�:�M�=%jh�}R�e�t� �*6�8. $����g�<�� F�c�4:"���x9�&��hƪ� �T�H���O�uF��O�a��çBŎ���ǣs���*��'�D�hT��~y��L����3����Eb�E�d��B�?ۨ ��-ޥT\"�I��"�`"ˉ�aS($�($]4��=Q4�ү�(�.O�\hp��)L�|�s@��+z��gF��:G�ԧF�xU3�"	�x�X�024O��_u���&H�>��}��eK���eg�l�.i�c��R�
T��_v���6��y�V@��|�0%N>N�<���-�'�p?��� 	YL%�VD������@�@�,�f]�mJ��
p�@�>�I"�̒<d�-�6D�����П��aPj!qL�ǵ6�TI<�C ��0)���0vf�"oMR�
��=q
�i%*�ZYz0!�+;���T垽	J�\�RO��J��bC��L]�ͻ�D.�!�J�8��.@�Y8�T��̓RL��R�o�� :�I��Ş�"�N�S�x�& �qn
-�T8���E !Y���D/N�ԕ�d�4B6:ҥ�K����@HF+v��	�%�FU:dȀh��px�BR]�%�EB���Ђ��G�.|���[�@Y.x��(m޵PU	>rJ�W�<�h1�Ot�;(D�L~���Ύ)�.�"fJ��Z�:DƇ�i����rM�/f�0�����Aap��KO�,�"�2�O|�I)	�q��
�/�����r�#>�p�A=h0�t�cD�9��(�`n�?�Ѥ�!Q=PQΰМ̊TCL)b	*��Q��$k�MȯM2�E�홇H��%� ��x2J�;"�ȥ�y��3��W�=$ޘ@��͹|�֤ލQ��lc��
�b<�1f��<�m�s)��!�"�"�cf����I�p	�G`J8%0�0����`3F%������CR��z�@y�U�`)ʇ�;!2�$��oe?^�W�"}
1iZ�9�n<�D�!D�"��$Q�JV}��H�Ѻ};����k����N�3{�|]y�M�7r{���v�
�d=��H��۪eח~�'W��	2�g
JT�6�Q�5�䠢��$ΐx��4{0B�7:���-��kS�T6� 	!s�ӱJ@~(;�O:6�Ji��Б0R4�t3q��?fÃZ7l��D��(N�\1�Do�ɔ)J�H�Do�(L�LѤD�c26���Y�m�,�8�b�U0Iaᆞ<u�1���(F:}j��� &raM؏�
��B�3�� 4V�hʄ]� N�(���ͻKF�j7i��X���	�̉�=�(Q�ȓSS12a�/r��a�$��$�P�(ue1%��ba�9}��9O��Ą՟4��{`ń�}Զ���"O�젤�V�i���b�*� )�=Oj���� X��דA��g��%�� �	W��@)��)N�6=x�
!d��(T �Lϸ�fσjR��� )D�D�0�� $ �S��6B`0R�&�G�L���IL�|j2`ފ}%���iY:+4$Z�D`�<�V��l����`S;%��YDc�4h1`���n�>	2ӧ����	`��t�Í�B�D���FԋX�!�dE6�X��ԾiN|�RQ�:���S-D�d���=�
R:b���wu�T��K?�O���i�./:7m�?H)�%0�˧,>�e��f��b�!�$�C�vɸ�`�@?�9�Ȭӑ�p��!a��>���#�kP<�
�g�-/���y� $9m����'�g�? Q�(�~�^�2s$�5n�r0��"Ol	R�gQ�b8�i�P��w�<!����w|�9��|��d8�# DO*� �'�3V�bM)n5D�T9�`�!EXq�4�� ep�DdA��(��I(ߓgS��[s�l�����L�Z�6���i�b��_�:�i��`Jl�c//X���{1&Йz�5�'�����"`��,���@L�\�V�x�+R�?�	��d�w��9M�O=����)v��V��&�;�G^&i��г"O@��ǟ�~�Z�GIW�ʼ���T:\~���gA>}�'[�r���Ç/B|�D���;bą�R�nHI0 hL��t��N�<�`V�]z���Κ�xh��"��Ɵ`#�e=��&���&�J,p�E�5�|"a�7G�`�c�gɊ$Lh��#з��=I�D	^�f$�6�O�� ��ޛL�4Qz��d<�S�lR��Ӱ&s����'�ZQ�GN�� ��� XY���}2@t�6-Z�^U�@-/�`MtjB<m%8��HC�'J�`p&�~����'�<#4���&�����W���P�O�@V�bJ<��n�f�� ��8�i}޹�W(_�x��)�1��;t�|ա�f'D�`�GHq�Cw��.��d�i���� ��g��m�K��s�Sg���4 ���"��67��)ӪZK��ȓ%I�Ui���ũ��ۧj3�5K��O2���O�i�u���s����H�O��A���jX����/7��}�F�5��$�4 :[��GC�cC��EL$����eP�Pya~B��KB��x�JH�d����hO�ѥbґt:ֽ"bb3�4��O6D)�ݖ!]4���Nw���'z�y���g�|x�I��D�\\���, ��a��
�4V���r	/�禅�C�FS�X[׃����h`e�4D��8pd� R�1d����k'�Ԉ@l U@�"E\�kA�ͼs�T�g�'Y��i��&�>�Q�ā^��	�A�� iH.U湨"��!T6ˀ�H� Tr������s��+�h٤��ex��j��[�a��� �/��Y.�����#� �[+��˱kïS���cj[
�ɕ"Jz����-50> ���,s=��R�N�y�i�00-yDU�jNrp@7-WF�xE0scБLL��$�p�nay����:k��,�;Z`dH��(��l��4��2'Y0���`�P�m��QC��pe#�T]����'V�B��pI�$R<��UEZ(|l� --�s��aD� o^xM�#��)�>L��I�B٨���ǉ�Vba�n�=5���(�E�T[��@�Y�AB
��#� \,�C��. 2��H	`���l!�:�%�$�gؿE<4EC�BC2		!l^"x��ɧ���N̢g[��k7��k~�4��"O���P��$9(��}U��x�c�<o�1[���B��)�E�!3���'|�X�پ��l2�K"/��'(�]��
<Uو�:b@�w$x"�)Z$��5�Y�!�|�^7V���`�H��C��+9�ay��#~�Hy��^�Vs���m^�I��ILoDB���7�!�M4qr��B$N����A�b]M��'���i���O��@G��)
��u�DH��`�^��y��Ù@z���EӫN7��נ[q�8���|�������3J^8%`�(sP|�'�vB�	�b�"\��玦L~l�D$ֆ h�C�	�p�(���\�0*�Ԫ�B�vB䉡�쨒w픈��QW"!.TB��:>�\h�7�_>o�d�	�%�*kxC�	�g�tV�u��@�Q�^�J���"ObQA��	�U[KL�T�D�P����yr���
� Ѐ�m>L��2�6�yBʄ_VR:��$ip�:�&�%�y���5]�8�`��7�H����y��C.Vu�X7!BY�]XT��(�yr�X'8
��Qe��\�8#c��y���F�N�b��*��Â��y2fP4.u�D�a��l�b4`i��y��Ǔ&s ��'�X�0Z�JԘ�y��>�,�{���X��[B�"�yb�ڊD�P�1�C��i6�U�p����y�{`%{!kP3eqę{U�:�y
� ���ٚ�he�R�^(�(��"O`�c��ԟ5�xaF�P�6����"O�(��h
#�T���N�=���"O|�:���Q8���FW��MP"O�`fW�=�*L/k8|)v��)�y�_55`�P���pgH�[f�L=�y��0Iq�ͳ$�=v�FC�ؚ�yR	�N���wk�;��[a�=�yB@L	!�� G�sFM��V#�y��+�=����o2��cn$�y�ɏ/�% �G��g�Rx9S%-�y!�M��J�>G{X8���y�o.n�YZT��;rPhj�MA��yB`�>��Y9�jNXh��k��0�yr	FO4����#"5� �V��y2a�	Q�B��!�y5.!2A��:�yR�,"|�h��vY0){T�ϵ�y#� ~T�A��.e��!�����Py� �%`�ڨR G��3��+�^m�<���(,���T�Q�J�V�ȀB�<���U�F!��aN��|X�[U�<9hT�W�d]zQ �f�>�
fM�Q�<9t@�n������ĹGٛ#��P�<Y����6�>�L\h(Fe�<���)\nP�q�\�4�@4�1l�j�<�R+p4�􎒣~Z4�c�[f�<����/R�@X�vE�99ʨs�![E�<��eYUt2��%�ސ@�l-Z�Ė@�<1�dݧNa�FXǰ�9�nGC�<��#��V�Τ؇䖵�L��B�x�<�7��[�V0`s慩?^hVOw�<1WO�M��@�K,tW���l�<I���c���
�H0,��C`�LR�<���V�x��ʐ:J�3a�L�<є�Z;�]��H�=�|�#���r�<QaC,)��O= ���R�$�:�'�f�
C N�}XK�n4��]�	�'�T��7���Kͼh�àԼ [�4!	�'����LM1M��!�C'L9
_`=��'��)Y�J�0:�� �be�+*0y��'fn�q�Ϳ;�x��FS�D٠�'/4���a�G_���r.�8���q�'8���$�V�w�ɂ�)�5(�|���'c���֤	O�`b@�Qq�81��'� ��g�Z��e�gm�&n�a �'B�ѱ%���I���~l܉��'.Xat������9�hh"�'��u���X\mX`yƅ��3e����'H�Rn[�Q���ȅ5)����'�*�FH�Lۆ����=dH��'h�0�ᜏ�����Z�Y�*���'uf�y���:�2Q0���oJd(�'�D��a�1=��,��mg�M��'�� �텳0��1���Ax1�'�~My'��ayzi�w��T{�T��';^�(%��=�A#�)N$\���'� PhE�Y:RJ�2��-O�ʕ2�'VV@(���U6����C�8��Z�'�5��k��)c�*>�0�q�'$���2e@6J�BH�����`�'�\�Bu蔔�t��vA�y�y
�'���Fdά]�@ׁ}�"���'�dY��?~R�Z`$S waA)�'�"�K � �v����;1ޱ)
��� �%����8��J)�B��"O�UH��C�Z^ D��d� ��(�$"Op�e�J{����Ab�6H�9�""O�9)��D:J��<�����M>���6"O{a�H�d�du)�ؓs.���"O�C��XVfh�%�߷` �(�U"O�m@Fa
�,4�<(�J�Դ:�"OF!S�� _����Ɠ%�03�"Ox� u�Fki�骄f]�8?<���"O��IvdD}��-#d%Ю7�A�"On���)U ]��2 0e"�"O\��g��2K��80�"�$2Mu"O�dk3��&@䭺�AU>A�ذA"O�Jv�W6@�z�pǃ��N�qr"Ofs�����\��@��
`�0Ӂ"Of�'D��l����/֋fP&ى""O:�Y!�)^tk$�D�n�˦"O�;4�5�ؙ���	�^l` �"O�d�4�ҴVܢP��ҚFs2X��"O*I�뚑�θ�be )Kzn��"O�Y!��Y5b�HhÆ�?��I�"O��Q LϰU'>��M
�d٣t"O��6��$0\�-��a��"O"���n��_�H��q�p�H(�"O�(A�X"e�%
Hb�U"O>D�B��N�`
�W5l���"O�@ch�]b���a�'T��W"O\�;�J�=B���"�1+vhÐ�'T�&�Ny��7fd���ȃ%E�g���y"�
C��YZ���(F���L�޸'
vI,*(r�@��IȄ�4�iҤ%�z1��}�!� �-0��1���j@!��`���b���?�&As�\9)����}�A� ��%24�@���.�p?�KZ�cE�A��-=X���M��}�RaئkB6l��q�T�J��|R�U.e���J�C�A,��A��@��O��ŬלX�Va�>"� ��Op�����e��0#T�Q��NP�yB�ѩ�JT��I�D[�O$N������^� �ɴW��l�DH����0�%N��}>E��O�TM���T�8 ��2&���-h��Z<9���I�^��dS�/[�ݳ C�% t��D��.{H8�rX�6>���[�,B�+��L��ҧ5�n�
JD`�I�R"�%;��4�0?a���r\Lx��޶U�|�� #�Z@3�2��E�ˆ�	>�:�`5��	ql��}�&����b΅M�~��UJL�'�n	�C�^�P�։�cIV��D�'}�~�b ^
k8��y��M�����O�XA��ΘH1x��I|�>��jY!C�bL*�FD�*�!�cL��<!��Ʀ7eP���	ѡ<̺	���6!5JS�#�+&�	ംV|�p��ɉ-6���B�'ؚ�ٷ��2D�����F�\�e�@���͏:B]`8I��\��u���b�]��.�W��Ʈ�Ge'	�L4pt�}�s��'�h����*�V��!ɸ��g��՛B�
d���;̚�x.ԠAH�,��))�	:V���6!���EN }ꑟ�X�P��H�1�,��.s��`����P�B|�⢂)M\�+����7���TQ��ƹY�џL+s/!%h$hx� s8$A	0�3���q=.U)�3��9��0�)Zy,�y���1
�ld�5Z @6|��P*��<n!�����%*��BG^���R 6ܸ�rCƚU��u36
Ԁ|���� 4�n(8�x 2��#J�agf�|(!��H=��� 3���F6�ͻD[�8�����
7��yL�"~Γ���e��k
y���3IH�ȓ��m��#��c@B��@ǌ�j4`ϓ>�qZƤũq���D�{�Ġ�r��9�0䳷��a|��_�� �UJ=S�< ���5`���v��4H��`�']H��U$�n^��x���
A�����dH0��K'�(��m� �w�(դ�;q������u�<�D!S�!hd@�T�i�l�G�ƱJ>EH"�`Jӧ����w���B��Ƅ�� �/�y"�	w&|M뒪ط[,��憣�yr���-��a��A��� ���d/S���a��Z%ApdyP6�'� ѹ��٩'#�fŝ]T�|8��ْg6 � �$�y��P�Njڴ�!� �|H��#=1�hߡ�֢}j�-֚Y6���mү`�p4�][�'�>�{��l�O�<dAK fuJ�:ԩ��G8���'�VYq �LS�!�(֍<�H5�2�Քz�L>���O�d���2�Q�=&P)�b"OR��2�W����I$vKh�i��iX��:��6P��5��C]�M���+�p!;p��60�����/���44��Q�IT�(�s4�G��z���� B���:���	1\O�1��(Z�**�ɗ@�X*q��d�IV��g ���'��A�ADrl#Bj{�Fl�j�f���	-�yB��i��:��gČ�I����X������!aJ�~�b�#Q��8CŒ�'�h睻c�. ��1E@b-��@Ƙ|��B��&�"�+dس`�p���j�x�B�B�cG�%�-7��qϚ<��[/��_>�K�+�t �@	�)�z<��	B8) ��ݎ,҈��}xV����@8������.?u�T��"I���<���F��EM�]�RTvNQ����#��n��'+ k�G�<�2���T�g��1�0Ɂ5b�zR��hh<���G�nEi2 �94mv��'�	?{"$PT�T�	#{�` 0h,*O�O%��ʴ�@���-�vN�ӧl��EI!�dȜ�B�XC��,�@!*��J"�����c���%�H���@�Hc�I����E�qAW�m�vY7�&O�(��vK"D��HTǗm�VL2�ǫ��	[WLC�E��+�% �ȐJ��ݰt�0�g�'ӈ�(LϠ1<\� �M�7kc<E��ka4Q�g�c�R�1�>faс�^��G���Q��k�3��MQ6g�:T��Kϩ+jqG{ҭL�hV��q���%���Sʪ|��/K�Ly�$ڮ1t9k�r�<Y��H�T�)��R s,N�zD�L�9�
�s�]: �D�P�X�)��s�P��!��&.Q��/�9�D�b"O$Y�ō���AN@Z���U�s�yЕb�8L�!��K�8x�r�g�'��,"��6^�Sw��h��Pӓ����H�j�~kE䐳+l����@��9��Ԡ��O�'EXl�b�J}��cႭq���kF�5�QMM`p%�0���Ojd��и�Ƥ\ ���,�d�b3��556T!2�u�8#c"O���!�6P(�(P2 _7~�d�T�IcE�#	��(cǑ�{B��>��CHO<�y��ٷ��h`�	|�`yX�߬��x�mC�\ؼ�C��UU�1����P|йu�J:A#����1}r�ıp%ǜXҨ�G{�dغnqbh��B %,���-Қ��<���H�F�RhzGE�%6.�c�M�0O���&�!	0H��u�(��d��qla~��n�X�1��(fS/���Q7,�PV��	 ��)ؒMZ�;���cB���ӚeX�q�'���
�i�%�*h�2"O�49���"F�i�F��-V����&"H�e���0B��l�X�r���k.���'"�i^�8A�e�q��8��Аx"'�0Ġ��@.YF�: J��M>�K�L˹dd��E�'�X!U�� ��!3� �w��m�˓%B21�3���e����'�h���AɟaOةؒ̍�8v����'Œ�kw�"y^����=0��msO>��S�2��ySw9�,�z#V�5*�(P��$� �ȓ-�$pr4-)y�&�)ъ�
4 ���
����4��E��O�lUO�� ~�5�s��07X� "O��h��M���1J�
H�"O���ծ=7dm0��$E�:\Y�"O\hC��Gt�A" �@���"O�%��x���`�B�!��A��"O�=J�	ИNM�0�$
� �NUh�"O���t��
���K��h�����"OP�)oL:h��@&�B���]��"O�%!��q��s���i�d�w"O�l� ���iwp �箚4C��;�"O��2����k1.���M�;���$"Oi�E�J&>�� b B��bL�Yt"Ov�����u�\!r�V^�İp"O���H� 8��`����/K.吠"O� t������(J�L1�D@�@Ob���"Od���ճbFe�1!#�YE"O�P�w+[�&�y�ؘ����t"O���KV�n�DA3͞	���I�"OHmp�D�Mf�͙�K�:a��m��"O��X��Mv�h�p�Glp|,�u"O�LR� � �>��È�sq�f"OV)"��&x�$���gը4t���S"O�)
!���!�ѡP{0�X�"On�BA�<p��.�?J}|�"On�FA�4h�0��^�d�B"O��y���/D5re�ȫ���!"OF����F�Z��U�'m�����"OiaTm��cr1��+��qks"O��@���|0,XK�ˆ
!���U"O���5_4Dl�I�W�\�܁(B"O����Nۣ14�0��uu|i�"OaZ���=0���%�o�t�"O��c�O�|k�=��N��D��q�"O"R�9�P᠗�^ XD�ʵ"OH�m�xӂ|�+V�
��@v"O60�C�I��P��v��k�"O�U�5B��*b^�@�/���� "Oi����ކ͛p&9�|��u�P%����?h��$��b���c���@aVx��� W!�ĀI9�dY�לp�>��?oB!����eK��Y��0PD�C!��Y�
Z�+��A�gr"E�_�g!�ċ��@`�£� a^�t�D#K�|V!�d�%��<�G,ľ9R�MA!,�+kE!��J����7CC�c�\�ڑ�K�s�!򤚧�X� �^���y�c���'��#<�����i:��<�c���W�Δp��:)���P']�<Y�lL5F��J>E��bW�90Ԏ�q�8� 4W)~e��A�1O�?�pb�7xL�2��׏� A��Œ%��b�P��E2�'����	�ҹK ���O�i��̕J��b�p 3%2�S�S�f، �IچE:�H4�&���O���u�lzC��9Y)�ɳgƂy��B�	�.���,D& Z@�*E?)<�B�Ƀ˾q��	�,2�>���H0f
zB�D[�#p�1C$z�)��[jR�C��4���*J9,p&/^:�!�dLT�d��CZND�qKP,V5aB!��9�p�v'�0/�>��V*�+:!�dR�>�J�A`�I�y�i����1~!���W��0�N;w^�i� Ch!�IO�����׊Zm�m`� �n!��(3j�-�;:]D�s  �!�䓍^�T��m��sN�\(��#,�!�d7���c��6�T��3�]w�!�d��`R����M�N�i)���PW!򄐐x�]�W�Ңx�$$��XbT!�ܒm���7���D0A��:g!��З)_~�����3:�b�AЂ�g!���*4GN`3�D�"E�\pKs"8M!��߸gz^���G�S��d��"Ov ���q���q��(�tHh�"O����% L�yH�c�j�܀e"O�1��M Y�,��P�̌�"O����L/ �1���J�$�d*O��eO�c�PA�]9iP^���'C�i�sj� >*���u*�r���'6p}��'ZF�0� ��L�d�>�Z	�'<\��.ˣg�6��m�X��ؒ��� ��Y�mܲ\9�������jp"O�ZVė�gN^<3����G�����"OT�y�����,���-Ǽs��v"Oz�;`��:H���,P�#��="OLY������P�	.۬�c"O�0�N�C���w�]�-cyYW"O�Xp��ε+O���$'K> ^h5�V"O���"�[�q��,:q�ŗP&E٦"O�2睘�>Xx��W26�,Q�"O
D %,�N\�Voȟ� ��"O� P2�XZ�����+\�b(�'"O`Ԑ�I�x���`J�
��d
�"O���n�/O>�q�<�\!e"O���у-b� ��[6w��K3"O��ZUcV�]:���P��"hh�*�"O�A:ǣR�A@�@�E6��"O
%��oM1?c��z���#�l8��"O�,���Q�^ř5Q0ݢ	JE"O�Ѣ�n:[�ҤpաV	,��`�"O����D�9���v�1"B��"O,1�B,ٹ]nn)��˔/6d��"O�z�,R��q��к"�f	�T"Ox\�sǒ�~��C��(�(�"O��w�ƪU^谰��%���B"Oxu����Lr��R�

t�*�B�"O��4.\���\���
:	�N���"O�4I#(����ĥC ^"�D"O�xCZ-���IՆ�jLr �"OX�����Y�4ܚ��^�vg���"Oބk��Y"vE!#Q�_]�l��"OJ�2�	A�b+�(v�n��#"OZ ɴg9u��"�� ����"OxQ�@�l�>s� N��@|��"Or�aa�^u��)�Ԑoʈ#0"O �е��//��Q3�9R^E@�"O�Q�D��6�bQ+��	6� �"O d2b�&1|�IA��>��a`�'��@���	l�֭��@W0��'M�#�лf:Ik�d�<(p�(C�'W4���ƃY�[W��Wt}��'�>��g_�#(�y��AR�����'�@ 2�h�a�|Φ���'��|�b���~�QY�hI#n��'��A*��Vd�B���Ε;�'_jE�d&ك]�
 ��Jx L1�'=�\)����F�I*Kz�F��'˖TC��M��œ�������'�4�ŬI�G�x�����c�`���&\� r�d�[�ސ��,W�~��ȓ<�����
[na�Lv�ӨQ��h��S���`'	~�\A���0$8�T��yz|�gh��$>�Yqրű�vņ�"Aр��q���Ё�ȓ#���R�b��?;�I`��r�Z��ȓT&��q`ɶ#-�xa��<-4.��ȓm��K(g��)��Ҽ
�	�ȓ�d��d�ϷR���ٴ*�ܝ��/�`��Ġ�� �J��b��n4�)�ȓFd*T�_��DЄ�͢^�� �ȓ3+\� �!B
��b�R$�z��ȓNg@�T̼);�����P�hD:ԅ�&���(��_ct�)�G�ZI���ȓ.�|���h�z�J�3���T4��q��!H�M�����/�����S�? �i �N��h��!�L�&���"O�����`��ܶeڔ�Q"O"��q�2d��M�o�BEE�"Oj�2d�;M"���H�D[^ h�"Ofػ�X8Ȝ;f�y\�4��"O��Ҕ��Qz*ĻD`'��*�"O*�y��%^oĴkЀ��hzj�"�"O��7
L�Mq�P L�fhZd�a"O qň[�m��z�/ū���°"O ��o[�$+*��.	�K�y�"OY3� )Zv\-�LF+N� �q"OB�S��M�1���2`Ԓnل���"O�]��O�ut\�(w�]�r��tQ"O֑��7�8�3�ʚ/x��;s"Of�	S�S�`p>�Ai�!ib���"O��Ò/�7K����	4��"O���%T��p5��fZ�g ����"O����C	����S���r�j��Q"O8�p��@�K�����ρ�D�(�0"Or|@�ɑ�g"�Sb�O�N��Ek1"O|e@�"Y/H��Dȯ�<��"O�
�.@�T���i�ݱJ�t0��"O�)��-Q|�hR�e@:-Q4��"O�(�.�;z?��8��V�X:�H�r"O���$됈����S6D%@u"O�5��)��G�l��d�'��c"O���b�ܝvQ��"$��
����yBO��9����ꀈ9h�I�/�y҉�&Ȯe��OCD�����h���y���&�>$`������@��yR����x8Wb�?y-.��dh�y҉N���B���n�Ɓ��;�yb텩	c �Bw���^����`��yB�D�HX��#ސ)[VHĢF*�y��GZ�"��F-�V�L�v/߸�y���a.@ 0bӆB�Ե���y2��s�T�Ң7���R�y�� j`Y3�.�6���C��W��yb��1hp�8#%�+�8���J���y�D���� đ�5ĬY�0���y��8s�:H�C���7ϴ�1���:�yr�K�{��;�%Y2t��D���yB��${��$���+A�5� ��y҃��&�F1�M%pzZi.��yb"W�wS���`Ѵ�����y�	H'략y�f�2!���`�L��y���<W@ahv#܌Y<��CG,��yr�Ty�t:�O�d�!�y�ʈ9W�\a�AI�0�F1� ��y�X�k�T� �J�whuf͎�y��ݴ(9��QQ�=�\�[�!F�ym)W]0���E䤽�A\��y"�7'��$ǬH�1"��QW�	*�y2��6ut�ؑi�4�`���K!�yRڃ/C|�v ���"+^�yR�в)��|��"L�9t�B2�T=�yb �l��#��w=E�$C���yr�C߈�A�"ʫZ���Ɂ��y2�ѐJP��ӍDQ��y	5�yR(P-��H��;8^֕�!�Ǌ�yR�$`V�	k �0,�"T
1�͵�y�ݨ���C�
�T����#�y���$�0�I��޽N���R��K�y���W�>�6ѩJ��Ћ6�=�y
� �qH��;sFH�%�� �RQk"O�Ŋ��S?g��i�w��-�04�"O���	_�@2�͔*���"O���.��ԁ͂��<P�"OLU3v��)�.؈��O9�"B�"O\ȷŮa�$q�g�9m��ҷ"O�(��(+|(r��/s�9��"OpH�&�/~��qz���T����P"O���ؔA�`�#Ӆ[�3�2�"O���7�V�+A��I6�&e]AA"O4��&nɑS����/AS\[�"OD�:�l � ]<i���M6oZ�6"O���o�g%���r ��a��3&"O��)U.�)�r�����GV0C�"O8Ac��"C����	4-���W"O��ь�o����D�9R�@�"O0q;C�M�'�P��M�� ��̑�"O5�T�>lQ�8�bT���"O��MY�C��8)�?B� �� "O Ń�[�B�t���$��4�"O�7JI8y� ��be&�T��t"OYQ��Z.���`���x�{@"O�q*V ���r��o&E� T"O"�!H8.���t�\�6{�z1"O�Y���?=�>����6^��8�"O�ةV��
1b�� L"t�D!�"Op%)����o���� ����S�"O�=8�M�n�����N��Sy6|�"O�u�k*v�3N��:PQ�"O.�)4l�`���i��g}��9"O�j�fס&�����+j�SW"O
|����@�܄
��U�[c Lu"O:�����N��<;�I�>~S:��#"O�E�G��_�:U"��O�����"O�A�́/5��9w
��~�=�"O*��ٻH"V��צOMeБ�6"O\`�qJ����Q��eҙMOƙ�S"O�h��ɞ� �C�v8�$j�"O�����(@�Qz��j>�I��"Oҍ��lW�
�b)�&d�
C�.$Hc"OE1��E�L�硋6~��"O��[�i�&Nv��b���l��1"O�I��d�z���p�zxc�"O�i�����v�pQ��;I�R"O؉��,�p˾�k'#P�o���"On9��M�&^�����H�>7r="O����(BP`4�&˧X�UcT"O��4��j�YFߚ�4"O\�ha��BoA�5�Z�y�l	�A�!�dN�vR~ȁ�@͓-�n��h��t#!�D�sL*�JGAȫ|������T�!�$���4X5�N4_z��&��"�!��I+��d�uK\4Bu�5��AԆq5�������M��OH����O��$iӨ�{�n�+@|M����%ibX����g������|f��{rx{Aчf�r�U��dlI�U'ɮg���i�nB����ɰ��N� v�čz�؆=D-z ��?1��I剀MCt#|����u ѧ�!LLXC�k"�Ҁ�a��ğ,&���ID�'��-�d&M<	�̴�u癮Em���{�,u�����O��oY�D�'ٛ�%݌O��8*� �]&i8�Q��~�Mљ6`�6�O�$�O��O�	}�JY�$+��L,!�*��i�J���%cڜ����p>y�a v۬�]5���E���Xi:١aP*��u���ևIP�(ư���E|���~��R� En.��AOD�s�ֈ�Q/�O���轢��[y��'��'��ia-B-:!��c,��!@��)�{"�'� H���x�z��#nҰ(q�m�!	��q%��`ش�*)O)Z��A?� ���RmZ�~JZ1�Q��=J������	g�i>��I�:�������#c�Ηh�p�$�M:+qj�ӶH8lO�u0�c�o�ԕ���(���]-E��qAQ*]�lRe��ɳ.(,�D�O6˛*U��.Up<�rG��y���ĩ<�����S'X9�Q�S6J�h�x�oZ�w��C���v ��A��l�A�t��6L>�7�lӐ}lZnyr�Ԗ�6��O�c?��CC�dx���>T�q+�M����I쟴���5�	쟰%>�x'(^�)Ŝ���a�,nu�epT�:���Vi\�`�:J�j����)VHu�yՆ�<d�)������O$��7�'��5�I�~�&F�������.�@��e�X5n=�O���<QB��5d�z���X�|�浓�'x?q��I��M��i��4b�����ƛ�jg�}`Rə�u�MS� �;b�v�'|�)����?Y��M�㝿w�p��%Z�y�0�Se-I6ykE�>�*���>�O��)@�J%j���l�Q���iC
��8$(������D�Yv�i>�#}�'�X�i6⋿x�|E�B$�$?����DO�Ov���Ԧ���9��>��BJ��a����ү[�!��i��ub�	m�'�j̋u�Fl�8p���U��\я{�N`��Ym�M���rڴ'��b�ǒ��h8�E�Ȝd?,���+	��ĳi���'tr�|�O�fI[)A�8S��Ԅ)��-��Pv���7*�j��P#c 	45@�G�1A�����k`ӈ��E�N�N�J�u�'�^����*_PS��S�^h����T�
�����O�lZ퟼�'��Z��n��
����PJ�.I0��ќZ��B�ɲ �ޝQ��J�<$R��T�T�ls�,K���d���'B�'��;J�`�� @�?�   �  A  �  k  v)  �4  {?  	K  pV  �a  �k  �t  ={  ��  ��  ͓   �  ��  ˦  �  P�  ��  ��  V�  ��  (�  ��  �  V�  ��  ��  ��  G  � 5 � � ' �/ �6  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A��!'��E�L��OL����A�*C�DZ6:��ga�3�a~Rk�>rk�;]\M�`��]����aC`�<9,�mj�pV�L���0+t. _�'"�?�w�M3s�r�k�$ޘU><�E D�"C��	��9��]U8��<D��"E K�Q�R�S�]�kg�ݳ�N9D�$B�f�$^ʄ�@��:)�M�d�<���S�!���D���<J07F>|9B䉢.����+�A'� QȀ�x>�C�	<,|@��Y�{�T�s��/F�dC�	�epA�`OE�5��ē�T�C�I�G8aS��+s�Ԩ䎇�jـ"=��T?y��HP�.�k@MP� "D��2��^�&�|��GM�/b<�eA?D���kM�ai�A�$
�x�l�At0D�(�ꊝWf艫f�H3nj��V�0D��"t� .Ş�a �o�Ppp�0|Onc�,�%T�J|�u��-UN�zc�;D��*��ň^�X'MD
4D8��9D���$瞶#^=���>��}I`<D��Z�Q;�Αel�pJ���&D��s0lʚc�@�� /^Ҩ��"D�8�`�+sP���Q��!x�����L D��Xe���@P��XS@����9�g2D��s"�Ð^��lQ���\(�X��o-D��
��������7��k�`�'�)D���ӊG�h����#�(hP�|�g�)D�@�P�P��l��+Ԧ  �dS$d&D�d��*y9xi@o�alx�2u�6D���J�Y�J��5-2PJ��5A8D��� ��R���-\Hr6F(D�\�0,Ke���Rρ�V�ڱ�%�%D���s�:Uy3�_\H9�*���y��ԥM�쭰tgI�v�<l@T���y�����0��|l0�C�a],�Py2 ĂF2$�ʑI�<��[E�B�<p��)dJ���U�)�<4{��E�<Iv`@�{^̀�nM�L��q+��DC�<��b֢	�0<;�CO�1�V�ƨ�Y�<r�]C�����7�h�+c�}�<1����*:֭X1Q�ܡ�l�h7!���V`�wa�6K&-h�_;&!򄟫q@��Ч���%��.W�iI�':��"�*�?@	�!Iq�U=8�k�'4|EB�H�$*�2�ʀ%�9 �d�P�'9X���Ry��@(���	|��!3�'=�5R�m6y�xE�VM
>t�{�C�2n�0����-�-x�ڦs�(B�7qrBEF)�:�h�C��\�0^�C��7a�m�'3p�p����YxP�>Ɏ{Ғ?������P���>��MȦ=D�� Bi���C�[�ZP�!�G
_�*�X���F>"�d^6RyF���
�&0|A�P�7D��e��(�X`4N�q\1�lwӂ ��ڸ���	��8 �`���B�̜S3�I	�p��DvӠ����%�	Xp&lYW�!͆0��'�Ƀh?U��w�_�e��'k�s��.Z���+V��! ����'�5�GU�����ڿ&D�ڟ'��	o�S�O�L<�EAW7��ĪŋW>o�RJ�'1�U�b`J@�H2�D�8�0P��"�'��ubԕv->M��+L�q�=�
��ē���KR�.iX�f��"�F��ȓ9��b#�D�,�Ĝsf��2m�F��ȓv&��y�e�#p<��%�	���ȓi�d�����S`Tqs���
[:��=��'��>��.@�i�S6O��L�%�]�qN�C�I<0h�I�,�'K���!N����O�х�ICa��G�S~8٥��� /�B䉀a��)��:Мɐo��b 
�'�D����I�&�*0�V�YEኈ�4�/lA� �?���iG퓳Ķ܇�\Ğ|R`�z��@��c�ssṄ��Ҽ �&K$�&Ib��c
�ȓO�*�c&�%����Q�M<ޱ���	e����v�DO`l�!�:��s77�O��Ŧ1��H�q�&Ce�֧�xap�Vrh<��F �b-H��wS�*U&�<SC�Fa���,�$Ǭ)��gT�<1k�~�d���*ƋyW\y(r.Le�<��ӆX$��*d�MM�,l� _d�<)�D�� ����K
��qP���d�<�C`�aW�T�b�1/��r�E[U�<0��! 
P��&��Dfa4��Q�<Q'nץx�@�u(�K!�0��D�<y7�K�W�����J��^�Y�Mv�<��L�LLI����%����#K{�<���O�l6*�"q��CSZ�*e�u�<!t�TuB�HP$�S�;4VȪ��Y�<�����r�fx	��1q�,ʕ��U�<15�̯x��XtiB/Pz>܉P(�K�<R��.]V�3e ��$�e�BE�<a�	�����+N=JN�[����<!c�$)p�B�ٸL
AS�O]t�<��G���]Bi4B�.c&a�q�<ɒ!	�]�l�a���-#��ct�c�<�r��c~���5!�j���l�_�<�޿�d�c �WBdL��E�U�<�s�%�P�"!U�(����X�<���V�t%nP��G+'�ث��W�<Y����w~pb��^q�DX��h�L�<!�d�%rx��Ԓ.`���R
L�<V�Z�"�]��bGt�$��fL�<)�S�.�t�qo�K��ёp]�<a/��w��������h������X�<�nJA�|���LҨ4R5Z���_�<���5�����L2��B�<i�$N�yj}cP�ϐX
"q1SOIz�<��Z�C�B��ǩK�����U��o�<I�㈤Z���qP�;����En�<)�N�-5i��b�"��ԑ�$�ZP�<���ʬ68�F�U�L���R�O�<�b�_��e��F�?T�e"#��N�<a6.� y�\���Ž�¤*�/BN�<�%�Q6^( p3�ǻp�
�Pc Q�<� "�OWC��	9unŌ�b`�"OfyÀ��Uђu�Ҍ�;�b��2"O��sU�<���[�=w�<�P"O��ɠ8�`�Z��)X���W"O���cG��;�0ti��X�.�4 T�'#B�'���'b�'�r�'���'-��
���-=>�ӂ� ipIe�''��'�"�'�"�'(��'-"�')^����ϓghrQ��M�,W�X� �'`r�'�"�'SR�'^��'���'n�0s�DݭW�P�s�*��{r.y��'R�'�r�'0��'���'x��'�E[���3��IJT6>ޱR!�'m�'�2�'�2�'���'��'Ht��fB
ju�0q���? �%���'Y��'6R�'X��'H�'2�'b�����ixH����V	}Q��Ҡ�'�b�'���'y��'��'2�'�^��A�#~=D���
*LZ� v�'��'3��'���'d2�'Vr�'�.���̟s���qW*�(C
6�d�'���'^��'b�'c2�' ��'��%���G��!8��� z,`��'7��'p��'�"�'���'p��'9*�ʃ�]�*g	`�'@"Jr �F�'���'@r�'�"�'Q��'x��'��X�P ŎM�-6���A�9Eo��'�b�'��'*��';"�'e�ݠl���dj@6Y>
u����@���'�R�'YR�'���'�7��Of���Le���u��7`��,ڵ�8�@T�'��X�b>�r���mZ9�@@c�,�mQ�a�!�y�\���ߴ��'���?�Vh��h��Ti��\1PБ/�:�?!��WQX\��4��y>W�R�O�"y�E�֌�f B��԰)��y��'��I]�O<�b�iId�j�ڵK�3!A�����>.O���#�+�Mϻzav���@�{ʬ���MV���?�'��)�S�
�Xn�<�E�O@��auF\�� �H��<��'f����hO���O��ڤmݔ4v)#�($-,���;O����mm����D^���ⵄդtj�Rr$�U��㟰ȫO:���O@��^}�	\�w� &���$DفA퐗����O��QG#ۡ/k1���Y�/k:�D��>ʠ���4d(l}yp 3za�˓��$�O?�	�fH���@�a�BP�V	���L��	�����<i`�iQ�O��<0Z6�g�S������[b5�d�O���Oz��5'k�4���$����hi�M��h`Q�In���@��������@e2����@U,A�C�W��I ����Or���Ot�?=y1�B)�@�4AD� ���(����O�&���05���H�1[T(2S��+ip�
���+LT���I���O�0I>a)OX�e��0�,34�G�c: ,i�'��?��j�3~nJ�r��
z��M�H��?�P�i$�O��'�R�'<� ş; �"��W]eZ���[=
ǜ����i��I�o�(`P��O��@'?%�>J��P!V�}��*B�lb��Ij����rf�`�Q	�C�Nj4x&�ٟ��I֟��O�S.�MK>�/7+��s�M��v�����䓶?���|�c剨�M��O�n�WMp��d�)��q���������O��J>�-O����O���O��S�^4S}�P $�f�&DR��O��$�<�V�,�	ןt��F�$GX� �X�F��	+t�
��[��$�O}��'��|ʟ Cv�Tq\����� 
�T�sw 0DGp���!b�~����
�|?iH>	���A��9a�@I��`�?a��?����?�|�.O`m1q�<�e�ʒ.�Pt���+3�n�	Cy�ks�Z�D��O�䟘q	�S�I��y�t�6i�&~�d�O��ᱧmӦ�A�yj������O�6 �Wo?E�}Y�m�:B����'�����@�I����Iӟp��p��&ѐ�J�����3^�a��NZn��?����?IK~���%<��w<�:p�A5DM�8�G��-I��[D�'�R�|����9>+��4OzE9����8$�A��?����'8O�(q��~�|2Q���@{�	�f�vqJ�D���Dl�O���I럌�	kyk�>��?i��.�&�Ye��L]�A�"/A��������>Y��?�J>Aw�^�ZE���1��h�84i�d~c�$_�!��nR���OR�1�ɐ)����sHx��[&TN1�gD��'|�'VR�ៀѡ*Iր��1]��(i��	۟1�O��$�O�lS�ӼSub�7Fet���%D�?�9�0��<a���?��{�2���4����_N�	�O��
B�L�)�X ٖC��p�t�sӚ|�S���I�	ȟ��I�l��g���r��i�/�~�RՃOjy"��>�-O���=�i�Ov��B=�&�٢�\�������Y}2�'��|���K�6:��* ÖI��di$�9Qw�h�����dh��<�Y�b�O��/!�x�Uc��
 �h+1L!Hzp���?����?q��|�,O`4�'[��
�P��G(�h�6�!�N�����M�r�>!���?��?\Vt[3�0�R�y����W2�+�R��M�O\1�"OM��������� ʸ` �Ӳ��]���ږ.���>O8���O��Od���O@�?q�� Z>|
���������I֟x�Iɟ���O���M�M>����3|xX�e��O4��@n_����?���|�p�U	�M��O�zrF�iM:p�B�d�^)Y6��=H��'�'�ǟ���ޟt��-@ u�Zg���Ԡ�)PYD�����X�'�<��?����?-�z�(R�eަQj ��+���%>O����g}b�'���|ʟ�}s�h&���c�#��a6L�7j�U���ϻE�f��|�t�O��I>I&�V6&HU�1�9J>N�·C�.�?���?��?�|r,O�1n>G�1���.i�5%�[��	������M�I>�'5��	ޟ���ܱW?l�Zs"�*�
I`FGY�\��)��tlZ�<)�c��0�F��(On!��E�>�����3CG�a+5;O&˓�?����?���?�����)�m�XH���[�>��Xzm�9ME�T�'���'������'�7=�.1x�#/C�L����R��U�P��O��5��iY�y�
7�p�h0`�\/n�P]j��@"i�� ��fa����&_�$1��<ͧ�?q�D�9-D���E� �3,E=�?I���?�����D}2�'0"�'Ό9a�R�TX,צ^�0� ��$@}��'�|2�8,�fU
�(ϚY��M���җ���Q������Oh���'?]c��O��ʯtERAxgA�T��ɸ2�̝[s����O����O���,ڧ�?	�?:�$�h�i��gx��谏X$�?�_�,��ǟ0(ܴ���yG��<gH��e I�mF�}	�!�=�yr�'��I.n�@nZn~r�Y�`��S�<RЩZS�A?�U3���_�6����|�R�h��ǟ��	ܟ@�I���[2�'w�\jwjH;Hl����Bjybj�>1��?����'�?�Q�I�x��aPt�Y�M�4���ۂi���ʟ��?�|
��(>Z�Ct!ːxN�ٸ"#�9D������Ċ��}���V2�O˓{B��xs�Ǯ[�I��ˁ�޽���?!��?���|�+On �'��B�y�v�+���=�x�E@�#.�fӒ�۩O����OX�D�wT^K�b��de�A�`��u(��i�q���
7`�0� ��ơH~���V3�TR�C��\���K4n�(�N�̓�?��?Y��?����O�\��]&1���e�D�L����'���'�0��|z�vN�v�|r�[$5���ੂ�K{�Ta����';����m�$��v����VJ�K�ꐪ�~3�<� ��Qk. ���'��$������'�R�'L�8;F�=<f@ЊNg�D���'p�Q�XѪO����OL��|:�B�	�pq�V��<T*��H���\~�í>I���?qH>�OE�@�OQ�o�(���i�.Z�bBD� 4j*���i��i>����O4�O�EH!だ!#J�o3_w��C��O��D�Oz��O1��ʓq/�f�ʬ/KF���ѝs���@SS��y�T���4��'����?9�J	�j����!8u�x��FK��?��b��9K޴���:��q���Ԥ  d%�fW�`z�a5ɑ6�y2P���I���Iҟ��I̟P�O�^p�u�;
,��A�U���T/�>)���?�����'�?�u��y�ΜV2�`1*�%��h���Q�MPb��iҖ�K^��y��M"j'(� n,1�
�ж��yb�B������m�'��������9\?d05�ĭG�x�#F
X�T[\e�Iן ����0�'l:��?Y��?A �^��� ��fI������A*��'U���?�����r���
F=w�����	vuz��'�mca)��ܢÞ�tN����S�'�&a+��LAz@I�1����LT@��'�b�'���'��>E��&7b�3-�.e5t�/�D ]�I����O:��N٦��?�;4��]U��"��(C-�6u����?)���?� D��M��O�n�6��i�5c=��`A��Jm�a�[4c9��yN>�)O��D�O��D�O:��O�B���lM�"!Ν������<��[��I럨�IY�'e� ����*DZ��K�(K�l9Y� �I��`$�b>5�0K������-|�Pr��5���nZ'�򤒋?��-��'��'��Ip�� ��%�
j��|@�I����	ǟ�����$�i>a�'7lꓶyr�S%o��1�ui��8Hv�)����?i��i��'Z2M�>����?�;D3��auDK�
E�]{d��>��*��ی�M��O� �D�S����#�I��(љ4�Z�6�|��d��L����0O���O����OF�$�O�?�)�H!�^����ssm�ڟ��˟8��O�ʓgꛖ�|�2��P����Z���<i��'������-Ǭӛ�����Ã����+e<;���F%��y�l P�O�O��?����?���{d@q䁉!v���Y�����?�+Of��'8��ן�O�Y:�R�?3
U����0�����O�9�'w��'ɧ�)W�^O�c׊*�0��'M�pK���	�ܐ1�����- �B�]�I�Pi��;2n�1|����Y�)w�T�I�L���T�)��ky�sӤЁd (%���wcU�h�( �0O��d�O��nZD�S���������D���p��3�6(�e蟜�	��bLl�V~Zw���`��O�6%��� ��Y�AW!h���u&�i��\��<O~��?���?)���?�����i< ��"j�>f9=�3�0�$��'���'sR��4�'�v6=�r�����	0@����N<-B1#�O��D4��ݶ�7m~�TI�oںU��p���?g���dw�����f���A\��Oy�'O�Cܞh�n	
�f�5�Ą8� k����?	��?)O,%�'�B�'B�Q�e��d����T�����6U�O���'��'��'�ƨ���>\�h��<iغ��O��q��K��uY��I��?	��O@�.BmD�r���l_^�"�I��odR�'Cr�'���s�	
!��^P���N؆!,\��ƌ���O2���Oިl�N�Ӽ��I]=-�x��g�Mp��1�!��<���?!��
q6��ش���(C�\��'p�8yT���_=t��T���q�P@��#��<�'�?��?���?T�ںL̪يg�:�\m��a]6��n}�'�R�'��O���_�J��#ā��y�'%/5���?����Ş�v�x`�Ǩn�$�	!>:,�$�Fn��'.4YE	��Ý|BU�P��;�`=�ਜ਼�kL1��Tܟ��	ڟl�����Gy�.�>��bh��Q��їE�*�$�F�{u6�9�1����N}R�'WR�'�:PQu��e�����%D�,�h93�D_�L�����0�EɌ�S��k�c�S���Ö+Ű>�
$���ʎ9Bje���k�����������I�����%�	��K�CRc�������?���?�'_��ş��ٴ��=��A{7+8dB=���&*Ɔ��<����?A��Rh�ڴ�yB�'{�m�����	�x���L2���{Do�Pʌ��Z)�'�	ʟ���T��=p����ݣ*of��ơ�$�0���Οx�'[�ꓜ?���?+�b�a��Q�6]�'��y7��@����O��$�O�O�ӻ.n)��B��%���R�ƴ��ֵ�쌙��'?�'c������Yj��ԅp������$+z�!��?���?1�S�'��dզ�:f$�'�rx �b�<`fx=kQ�}�0�IǟLX޴��'����?Q�a��J��݁�cO,6�����,�?��O�8(�ڴ����`�!���R+Od�;�h�x����Ä5gÚ��9OD˓�?����?����?����I�D{ x��:V�:5+��/e��'���'R����'�z7=�LٲK�R�N1��,�/�2�b�%�O���5��	r�Z7�s���A�_��c�Y�TH
��Q�|�ܰGع6���'�D�<�'�?���T�j�������%�@M��?���?����d�n}r�'�B�'��u���( TT
5C!��\ƛ|��'#���?���'�*�	W�s�YĨ �?#ք�'�`��[�	F�	��������	�'���ufSN�!���g+Ɓ�6�'Yb�'���'��>�	2�B�
C4�dI�@l�1�I%��D�<i��i��O��N��[����
��Nې���O����O
M	�)n� ��,��&$�,˖,�:e3�eH4�B�G�L�q�G)����4�����O\�d�O����ܚQ��O]p��-{p���Pʓm�	ɟ����'?牘C�-�b�XZ�	e��"(=b�Ot�D�O��O1���JĨ.�专�ݍS����ѨͺJtt7�=?�"B�3�,�IT�Xy�냺Ta�,�7��N�d��D�0>�FW���I,��}�F옜�։���7U����/�MË"�>���?q��R_�ydD�6�� :�e�B��IPh��M��OBu&V����%���� �`kƼA�(�憲�F���5Od���O��O��$�O^�?�b���s�&-{0��2F���ڡ�
my�'�d��|�����|r�T75��΍~�|�T�pU�b����jy2ǅH�֚�X2�NF�DU$�+���*���o�|��XZ�'�@-%�L�'J��'��'�ر��#]7HY���A?v��L��'q�P�Ы�O���?A.��A0��.G��=�4�Yf�� ��D �O��d�O,�O�S�g���[��2n1���s���<���yV�L�jC���\y�OC��Iz�'���j�cI�or"����!>����'q��'�����O��ɬ�M+�H�]��qs�K��X	�j��<����?���ic�Oz��'�r�ЮR{���b�8-��kBb�6v7��'�t�ӳi��I��v��e�O��-�,J�̺`���f֏>�������O��D�O���O����|"�I�?��h���� E�� ����
��ϟ,�I⟠$?!�I��M�; z����
0�)��/L0x������?K>�|��P>�M˙'�<�[$�@�M�p"�"���\�A�'�L�$K�០{��|r[�������х��i�m� A����qiU͟��Iן���ny���>���?���X�(Pʷ�N��v�A���;-����r+�>����?QK>����u�d�{s�
zLs��Yb~��6ĠQ4�A�$��O
���ɳ$���@]���(M�}I~�ksm�I�2�'�r�'�R�s�u��"Н�N0a	��U
A�Nԟ<�Ov�$�O�yl�Q�	���F��i���S�.t��b ��qɮ�ޟ��	���x�f���̓�?ŀN��)�|�? 0Y�����ld���k� D�����#3��<ͧ�?���?���?1�-�-#hl�3Ƶ�r0���<VJHʓ{b�I��Iӟ4'?��Ɍ�敺�(�X����U�x��O��$6�)擧$n���,F.q�5f����	�S�ܿ!���'�R�b��ğ("�|�T��2VE/kPzС��P��BM�������x�	��S~y�>�� '��Di��o,8|Г�Z�R�X���;����De}��'���'�6�J�F�e�Ȱ� {���*��ß3.����̺v�1M�Q>9�ݜmƐ��3T7v��s��(`>��������I͟���f��g�:��I\�t��K%!O8#��Y���?!�O,�i>i���M�L>AR�\!!��`�� �p6��9�-�䓐?9��|��E��MC�O��W!@�r���8"ܨ0�t`�*�|q����O��kJ>�,O����O����O
�᠙�
��aE\�0&p}"���O����<IZ���	ɟ��	l��A9�����l�KF�2 �����N}�'�ҙ|ʟ>T�!�WE7h\)���k�����C�3�I;��Εx�i>��&�'�P$�t��A	
q$|x��O,\����ڟ���ʟ@�I؟b>9�'l6V�`U���w!L�qt$� ԋ�a��D�O���NͦQ�?��S���ɍ{	��Զ����E�{�~��IßC+����'D�E�eܧB0�!�ˈ�G\�	�f�6v�Γ��$�OT���O��d�O�$�|�4d��\9�i�(����R}��ß��I�L&?�ɗ�Mϻ�J�:<[j��P�"a�����?�K>�|r�a��M�'���i�"L��\�f�
�9���'-¬ʁ�[?9H>�-O���O�i
V!������3k�!���O��D�O��Ľ<Y"V��I����ɠ,��K��ՒS�h`�V�I�Q���?!�Z�����p'��i/߄�xG�$+���.I��ɏw��`�	�]��b>�hG�'����I�o��8��� +�͋��6��֟��	���Ib�O��«H����ι-�� j����S�h�>����?���i��O���(
7�a�CmM�a���>"��d�O0���O�4�|���{�R��<�J܈#[&D��J�&#�JQ D��&�䓣�4���D�O����O>���(z�8l�U�ܤQg�a�� �{�˓j���� ��ş�'?)���U��ۀ����T؇��M�On���O��O1�i�����6C��4�Z�����=�b6�.?aEg;Hm���`��dy�H��!���脔i�����4���'��',�O��I��D�O��ö!/�q��A�������O��m�U�Qp�	�ĕ'~��:�J]�x���)aADŲ��Wd����� u�
�f��At������!�l����Jպ0ZTe�p/m���	��H�Iß�Iٟ�R�1;���z��2:�1��Z�?���?ɒR��ܟ��4��R���h�f��d�`&[�F�:H>����?ͧ/A�0ݴ�������rL�Kt����HV��T ��i	�&���$�	������O����O��C�ԮE*bJ%�2�l"1?����O��q���dyb�'�响A�ڱ��A� ��h�@L9\��{�IџX�?�Oֶ�`����#KF���h��O��k�20Yv�Q�4F6�+)O�IX��?��%��@ �!4O�!ή\3�ط-D����O����O��i�<�1�ixXy-Õ-�B�T��*$)���'�r�'�6%������O�۵�B�e�ł��]�,<r3��<q�e��M[�Ox0�Aۖ��ȣ<QB���v(5�S�=���Sh��<y(O��d�O:���O��$�ONʧ%1�aB�C2��ze��|%"��P��'�2����'\6=�L!��aڽ82�`���đ+�.����O&��/��Ɇ���6-d���6��@X�(;E�9��c�z��	$@�W��A}�wyB�'f�%�~���Ga	rz(�W7e��'Q��'��:����O���O
���-"߾,y�b]�i�$ ��1��O�-�'X��'��'ɜ��vI@�dP$uɥ�G����O�HꐋG�:s�7MTp�.q��O�]Е��6q��C*�b�HJ���O��d�O��d�O��}���0� �9���,6��3⥛�#K9k�hF�Iџ�	#�M���w�;6�(O>�����x%��'���'�bf��J�v���C� ��/����X�
;��R�X2{�$�C��(J: %�����4�'���'�"�'Il��$nU/�~qTGB� V\C�P��
�O�ʓ�?�L~z������L@	�|Z$�L�C0	Z�H��B�Ş
"����5lb
�x%ҢD"�'�9�dQ�.OM8�B��?�E!;�$�<�Ԫ@1&�P�z4��"XV�`x��1�?���?���?�'��Z}��'f!��}U�+�͜�xx��'�x7M*�I���$�O��/_`���l)O��-:&A&oN��Я^�M#�O�9�A�J���F�2�	���)X��	�"R�\z\b�2O��D�O��d�O:�D�O�?���Ȃ�$ur���H�-e��D1�mCiyr�'����|�W�v�|B��J����Q��6�T1������'�����ԨD�F���zì2� �=)�/��A,T胶n<2������?I�b%��<�'�?I��?I4J	�*�"��9^|��ӓ-!�?I���d�y}��'�r�'�-V����@���!��R���b��	�`�?�O���a�)� Q[�M	T��8�� +B�MV�>�� �� m�i>E� �'S��%�d�&
"%԰H�MD #{� ;f�I̟ �	��$�	��b>��'(�7m���n}���V2u��e��gR��On��¦��?Q0P�,�	���*���!!�����:�̰�I�0ЫXʦ�'��m�CI�?ɤ��	��� �.I:���&����2O��?���?q��?!�����	>|5�`q7�Ʉm�-�g*Cu��'H��'����'��6=��[�a�8 �����H߼�����/�O���?��	��o�f6mg��9�-"9�p�D���'���pGr��"��
3N���&��<����?Q0�I}���Q'ʠ$�T�a���?����?1����PL}R�'j�'���
$oP�I��d�d 	�#\�U�$V|}"�'l�| ����2LH�<nȡRF
����D��8yjdp@-,�1�p`P�)� ���T6|��!�܃���KD.�	� �$�OP�d�O(�D3ڧ�?�F-��v���CēeX�a'2�?A _�8������޴���y�Y#��ғ��o',����y"�'�R�'M8L���i��		D��h�ݟP����J)�J��g	"r*-+�"4�$�<���?A��?����?��ׅe\�}���4����,��D]}b�';r�'U�O?��T:>l���
	*{h�b�;W�X��?�����S�'Q�\`��H<&��q #�HI�I����M�Q�DJBHB�Xl�$#�d�<��υ�3Ŭ����]�	x0�[���$�?���?1���?ͧ���Q}r�'�b�Y�ͭG�D �	��'k�@��'��6>�	���OV���O�c���!%�2����9d��y b�1h�L7-$?��#��	(���Q+u���b�M�4
A�Q���KC�~�,���@�	�$��؟8�"SA�9�t����P�8����� ��?i��?1�[���˟���4��B��t�g��2jp>���bY>I��bL>���?�'1�<kܴ���P?#��R�S�<��
*g?:�zf��nZ+m��'z�i>��	�H�I8+��Ĺ�l�g�`ӐΆ9/J�I֟`�'�ꓮ��O�˧2vi�fRH�����_�V(h��'I�ꓖ?����S����7���a7�[!x
���^�/o>�yC�E�mv�=��Q��S��R�D�	;
�Xhf�/��u��K$,��0�Iʟ���П��)�S_y�MeӜ8�)�u�U�Q���@D���5O����O�4oZh�H����ˠ#ˋ<�40d� �䕉Q������ɭ]��ul�L~Zw�d @�O�䵕'���CF��\$FQ �o� 6�Q�'��I�����럌��ڟ���[��!�,g��y���#=�10 ���/�듬?���?�H~Γ>���w��8�G��!Kµ�t�Q�s����v�'���|��D*H�Z���1O�\x�,ݫ
������R�u7Oнڣ����~��|"^�,�	ҟ :�o�&=�ŋfG�]�%Cd*���������IzyRD�>����?y�%�9�_*�! ��=B�
��DS�.��	֟���F�	^���v��e�F��+�ު�"�N�`�H�:�U�|���O�U���c":����%*K
eV�Fe�P�����?1��?���h���$��gL1�ġ$1�T; 
��	iJ�$�l}��'QB,p�.����@�C����r�d��k� �	ٟ��I�<Hq�ɦ��'�\l�d��?I��^,���V G�n�CġB|9�'��i>���ğ(�Iџ0�ɯd4����$��8����kѺ��'m���?9���?�J~2��X0�	ŀ4D !��%q��A�S���	�'�b>�S��@�`8B�Ȇ�#���Q��9�X�[��+?i�蕣sZ������d�!x��A!�ψr��E�@�������OR�D�Od�4�t˓Y���� �c уD�PEjջFyʭ�à�⟤�4��'듧?Y,O��X���!lމK$�?K�t}+"G#'�7�5?��m��{0\�����'������`�\ŋgH�"K���aen��<���?���?���?َ����#R/���9Bb8�
�O��X>p��O��d�g}�O*�}�Z�OXe`���A�(1�����L:Ӆ4���OL�4���*��V����"ܲ O�x ���=98���^V>��Q��ilFI����f�P@�&d�()X�9�熕g���W��u~n}R�aG$��a�ak)�����6ct���c*oe�����:y2�hʧDM�!�@QI7ET�_�2��+)�aR'��`*�������R��� {|�����I(����'�&�isE�r8d��P'<�B�*���[�@�+�ZN0t��ɵ��Pfi�z��&�N2 ղ,k ��o�np�1�h�� ��te�i�'昍t�@B&&ʗo�@�+�NҝM=n�t�N9_R�(E�ˠ]�R�vӀ��Oj���OZܚ�%��"md�b Hƃ23��p�
b��̟ ��7!�Ld��m��TrV�V�7DQ�%@����$�ߦ!� ������M���?���?�R�$���? zź���J���@Gϣ�M���?�2��?QL>�/��p���iD�-��`�q�މ��$ �}ڴ�?��i\b�'��'_����D�t8H�G�E�c4p��Am9s�ZXnZ,�6��?�(��h
�2O:��T�? ��zdK�^D�J�Ѳh͠����i���'��'W4����O��	%W�D\�l�52a20��!#b��q�Bǟ8��q�D��ȟ��	," ��Co*|X��\�,I��ش�?A�Ot�	Xy��'�ɧ5��"B�|��B�B/R�b������C��
��,yi�D�Ox��O\�O���4�D
��M��Z�)ߴ2��Ihy��'F�'���'�ٹ .�?���C��V�z0����+�b�B��y��'��'��O���S- vY�.�Wd�
1��<�7��<�����?����̙�'F�t킢BЄM3Fl|�����B8�y��'�R�'���v�O����8s	��b
�7Th�:��1;��6M�O�O��d�O��	�@*�	9L2u 2�Q��`�N�$�r6M�O��N�S!�D�OHi�Ot��'�&�M�v���Pz���"@��<O���O������c���
�2�r�ё�[J�r�;�KJĦ���in���ɲ�M��?����?�_����)Ůa�e맢޸5�$���%��M���?Q����'���(`�7��J�DҀ�ƅ3y�E��m����V�'$r�'���'%rP����ǟ�"� h><�cJ�7&l�*��	��M{������	Ĭp��$�OR@�ff����y&C�Z ��z��ݦ��	�l�	�<�K<�OL�D�?-f����<30F�{�+��H\�V�'B�'�H��yB�'f��'Z���G(�`	2 	�:,�fK��g�8��O�$���O=�� ��&�؀s��2��Ea֐x��'�ʼp�Obʧ�j�'nJ�Z�픷a�>�7NߎF0(Y�ش���OX��*�I˟X��<�t��/\�4Cd�R%eA�lZ)'��m4?i���?ͧ��?iw$h��8�#�jY$i��`�Z���O��|��xyB_.�MS��Wz�ɑ'HQ�<���$Z�z0��ݟ����u�S� �O4�C�.?��C��r�p�3gFX�>6�/������'��H<�!!�+3�yj�n��0��9z�̃Ϧm���0H��Nwy�T>Y����x�i���t ʷl�Զfi�4c"���#"���OF�|�@�DxZw���ц`:��xI$�Y:&�\��4G%�Q�(OH���O(���O<���<��g��[pB@�\�`4��{�NlZ���'"H%8��4��탑�i͂I�5g	A�:%3�O#VU���4�?��i���'�'?O�ӻ>=:E"�N[�yK�A����7��O����Oz�O�V�\��	�N���cI�D�U&�������ش�?*O���<�O��d.�	�σ|]��O�<��г�	��u�O�yb�'c��'���BŞ&�(}U��"�`Ӡ��Or�&��S����xyR�^�a������7969C�%�5ho 6��<���G�R���|����?��'�~���H6qh�bF�K��z��_��M�+O���O8㟰�Ig?�`Fo�H��3�Pq���	F��=���6 ���ӟ���矔$?a��OV��gӼ,4,��$��%���(�O����O2�O���|�����x�U�V��0XX�t���
�^�<a���?���O�Oc��'�?q���.2-Q��:s��]s��.z���'���˟ԗ����'�e� I��D� zB�큱�҅'\�1lZ��Bψ�I�����6�$�O
����@A��Zq���̵Y$<d�i���ȟ��	�����s�S��Xvi.8!�K�.}��ه���ֆ6��X[���Or0mZ��X�I���I���1l.ޔbū �F�����㔫	C��]�8�����J|r,������i�f�c��ݼ~�t���[��J�4�?a�i���'���'��듺��	w�!��^�O�� ���DEo�-%$����|�'��|��vl�(ya*D�aA��9rP�׵i�'�B�'�����O8�Ɂ
z����^p¨ѕ�=@��'/�	�/��I!z�D�Sҟ���ݟ�Y�F�'�1�gV5"����!ԙ�M[��?I�V���'��Y���i���ʽV����L�#u�A�Eκ>��E�<i��]�<����?�����Ӥ{\ ����O��l�a	�aPv7��`}�Y����my��'��'G�lʧ�`���j��/h(1�2��y�IP�p��'�R�'e��Z>-��O�$$eL>n�ؠ�%>J촸ڴ��d�O��?��?Ѥa��<2�܄��S�Y�u�����`T*u�0�s��?q���?���ʧ��ǟ��Y���w	�$M+F�jb%`�f6m�O˓�?)��?q7(I�<����~�̙�CB�)�d6���(�-%�Ms��?Q5�L�<i�Q�����I�v�v�����).PQ˳$��b��x�OL���OV��A�)�$4�D�?�`���b̤0Ӵ��,�R�s�!o�D	z�3O�Ăʦ�I�4�I���K�O�nC�bK��h _=K��i��8?o�F�'O����<�,�A"g��e��)~L,��K:w�\@b�i�"�oӜ���O�$�Ot��'��	*0G��6@3pHdT�ō�6H�8e�ߴTc8��?�.O��'HF��'�?���9���j&Fk��ĺ���$����'�b�'�˾>i.O,�D��\8�fL�)3r	r��<�İCm~��ʓ�?Ƀ)��<����<���?��5c�X�o�&}W`��,K�:���遾i��'l�듚�d�O���?��{d�;����I�Ȃ�^;����'D��Y�'$�K�'���'k�~� >���J� ���cF�@�)�:��g�i�\����O�˓�?���?!'$̑Z�戈U�H��[1m�[ ��%�p�����?����?��'�����|�"�ɱ�
��r
f�<#'F���'��P��	��@�ɞg	,������ҌG[�`P#��+Q3��C�d�OZ�$�O�D��.�8m�O""l�h������#�Ԑxt*���7��O���?���?�b�EY~��Me&�D�|�sr�(;8��&�����ID�R�x���I���)�O:���O�((w�[/��k��<Un�P5�%�������TbTK+�������� ���;�l5��)��M�f���<Q��x��V�'�2�'���6?�U#�L\Dx7B�5Md��U�⦡��˟T����ݟ�$�̗O�� Q޴6��PU��E-6�`ԣ(!�n�؟`�ߴ�?��?���O�Ԩ����\�C�}���xքȦ�p�et��&���OW� �'	BH�<M~�Q�Ѓ@*d�Gi���:6�O����O��D�G�IПT��R?���'��A ԵxS6l�(ڦ'��3���@�}����ݟ\���;B�r y@�e�U)V"@�
�4�?��0��O�.��Ǝ����،�%QŤL�Y�n fS���!Ee�8ق����Iʟ��	l�i�+T�������CJf	:��<&��7�IƟ%���	Ɵ(; 
	$�^�q���F����8�
��I�`�T������ß'?���O�v!#ܓ ���b'Bk��j�O����O8�O����O�3���O������%1��[���2�i 1��Q����O��$�O��'>]�����D�%�A��B)숀���*cr�o��$�����D�`��ݟ��O~�r�I&$�⹡Ga�(��1�ռiuR�'
�q[�'�b�~Z��?���T0���M��
t��L�wOB$�s�x��'��/�/��|�ן�9&�~�p�&S5(E��ҺiY>Y�'�B�h�:��O����O��'����C��4�� ��I!޴�?���5&��p�������5���FR�#Ur)aQ�.3(HP1��6�M���]/���'��'�2�%�D�O�	�]8�X�q0�ٙRR�!JΦ)p"�t�$'���O00ii�'EB*�(O@�`���*e���&%+�'�?Y���?���n)�'���'��d���(���%.D��+�0�V�|�_��y���>�yr�'?��'&x��_���}�����%�����	c�Z�d�O 1$������@&��X�,�֐�����n�=�w#�V*b�~�a���f~�H��?����?�I?�)_�e�6���έ S��{�Ec�p�'�H��G�'�dW�\Z
�P��<[cn`�'�"��v�'� k�'���'������u>E[��Ռ�����6�z����t��ʓ�?Q-O���O ���Z�$L�B���Ч���J?�]��+	#x�]�[�b�'��'7�֝T�䀪~���)*X,8�
*s�h�sv�թN�$�p�iFR_�p��Ɵ�I�_�H��|n��bGC��2e�c�	�:�I3�iK��'&�Q��'S��~j���?���;4������mR\ ��@�X��R�\�I����	�n�B����?�`���
Bʥ��%S7�,�(n�\�k�>O��D�ڦ���ɟ���(H�O뎈
L��\���%�F��eD� }���'���yr�|�T>���zӊ���!0[��4�o6+*I���i�R�w�����O*�d�O��'l剨���L�W�|��
�y
�iCڴx�`�ϓ�?I.O@�'��Χ�?a$��<�ʵ�U�i\��-ReX���'�2�'�"c�>�-O�$����E��1l�t{F��o�"��c�n�`�D�<ɒ���<Y�(��|���?)��t*�8䂄�N����A�0H%�Ӹi���'X�����O�ʓ�?��C@V��d�� ^H$���O�nyoZ�8���k�,��ퟠ�	՟��	m�\c۴�
e�F�j\�)�f��u��IPٴ�?���?i���?)M>a��~ �����c���4i0f���M�A�
���̓�?	���?YO~��<��c�l��0u��� "ɪ����T����ߟL$����_�.kBD�G%58t8r�Ů Z�E9O��$�O��d
d�4��I�ODDʔ��Bm~H�����7�n4 ���ܦ=��K�	�8E}��).jɨQ*�3-���T��/�M����?�QN��<�'_�S̟��������D��u��0SH�tA �q����ē�?������Fx2ݟ`�H*ݏNq��B��y��%˒�iw�X �'� p�<���O2���O��'�щ���=��T: �9?n���ݴ�?���)q|DxbY>}Q"oe��̀fo\�l�p�����v}p����i�R�'f�^����yy�^�@��cP���%����~xt�d�1����G;��S:���	���j ��/iWPI���ž}b"4��Z��M{���?����?i�x�_>u��;i�t#�!�͔Xyp��B�.IЎ}ڏ�y"b�9�yr�'P2�'�H舆a �P
b|��-A&u�2�P Iz�:�D�O��K���t'�d�F��U�&��/9��X� IP7�� �PJ��M�<i���?�������3�2)� D�&�ecZ_����i>4Ol��O\�On�$�O�(��Z�>ZF,#��Y no�iY� �(n������O���OD�����'Ĥ����R�zt|!���$P�e�'���'��'���'m�y��O*M3'��.lN���HۤmIH�IfF�<����?q����O��'�?)'� 2u҅"M4�F�HE'5��RƷi���|��'�b�>��'��x��� �*�y4�Օmʜp��4�?���^p�A��?��Q?��	՟����m��=d�V��N�2Ӛ,hK<����?�!N~���i]��6����|�ӄ��S- iT��'S"�'�r�'*T�@ (G7B�+!��	
�T���Z��M�����20+��.}�7�ܬ|�x�S#I\  �̑aw��Y��f�'�"7��O��$�OL���d�l��c�� ��pY���`Э��ᦽk梐[��|�-�~���?�&V�ahl���Bt/��R���t�f�']��'<2R�d�O]2�O�� 6�W�8\hy��3�t��o�u�'���n@���#c�0\���P{#��h���M��v
5*��d�Ѝ@ܲ9z5Ȇ�u{�P� ׄZz"������Y�D���<m��	�ݗt�b��Ɍ4{xBF�
B>�{��˙^���/J:D��Gm;3�� �dN�TN�y��8@��`q���"6fAT`lL��E�U��|p�J�4]tt�G0J���
�ۜ�rv�HT��`B�i���qL�.ic���B��'&�aIp�G�xmPPI�КK��آ��
�P���HQ��ypb��Of����&���0�*^#?P`!�W�>�ED �~<��д�����iy��'�b8���揳06�kf�L�I�6�+k:��qtBV�9.��gZ���x�"ܔm��d��D[��|�i��HQ�u/���(�3<n�q�ǓS�=�	�p�'xE��V�>l�1 !+ݟ1F�芈y�'�&�y�CR	?��P@Ā:AS��2�'R�6�C*���ƤŲwXXtBDiU\s�D�<��J�4U���럤%?=�	�������C�jͤ��vKC�G����	�d*$�ĦZ�t\H�D&"�j���S��W>U
,�4�F�;��������*}r��LBsB��x�X�U�S+�V�!F��/u�b4q��0���'���h��?�����O�\�J�e�,jG���?�8�P�"OZ�ڡH�x���5���V| T�'��#=9Q�T,x�Jӡ1XN����[+%��ٟ �I!�����	����'�b��1�ȴ���e�����g�8P��'3:�F	Q�̘��-�L��ႃ���I�  
d��Ǝ�/q��d���&7�3����0	0��;Qc燃�1�|�D5?����Ο�g�'樸��Q��i+G�H=F��y��'62���O��i��}p�`�>7�.	9�O�`Dzʟ�[�8jwm8q� ��w��(Y5R�iE<vW�&�'���'������I�|zF��25�P���]��\5�̪�*�~@a���'U��i�MH
-���Dc�}�6�R��	�X$�ǟ�|Z����֋�ʉ;pH@$#*&�C6��zu�V1a�R�'ў`�?Y���9W��m�1	��ɓ&_m�<��%�� r8�eœ-E ,s1'�h̓o��	ay�᜜y�v6��O��O0oXF�bR�ԧU�X�˦ML3���d�<9��?)�O�F����FB�(2,B�^�����v&I��	!4��8�"�-#���ԤY�R-�B�j0O��J�jӎ�OH�x��P.�z�Q�L�7�����"O��A,G�N�"��ĊI�llA`�O"mZ�b���d�U�=9�W���c�t�d��M���?iJ~��7��eSt���GC��!6f�"lˊ�#��?�D ��?Ɏy*��I;��ݠ��?A|����ǋ�[=��'�&����	ޅj�L�c�ԛ4����G��4m��	N�S��R�����ωW���1�I�6����@#JqȐL�)�bD�P�{�2��9�HO������ z�h� �=6d@���ئ��I���5A���؟P�	̟�'����f��"���C�w�䁣S�/�dI)@����|��	+Ip��AǄ@![�m���7p�O.͒�L
�����_�u��m)���y���W�B�'�B!�8���,OV�D�8tԌ�`l�%	��9¢E�G��B�	;��H�ï�2 "РbD�߶ys&�����'���M�8<��'��|��P����=&w��R��˦U��ܟ��sy��'x22���DN�w"�I�Ī�B��USA-�'8+!𤆓Ah��`a<)�S�J�<D\j4Ox���A�䁛A�'f���Y� <:��'��<��cR�2mH�ط| v0��'=�����L"���!$$��@��P�y��>��
p����4�?Q�E��H0�ɉ�y��ȑ��h����$�Od��{>u���O0�ON�[R�!R4q`w,��D�fe���'_Z����ߑ>X��cK�)��a�!K܇�p<Y��W͟l'�x�c��$f�������w,)�L,D�d!���M`�t�Sd�����i-����t�? ���Ơ�"�� [��P�)@���b�D�}A��n�՟���M��՟x���;=��Xe��S�
�����<�	vY���	L�S��O��AՉJ�'դ%&M=n�L��Ė>q�ʗE���O�
(0��$j]��yve�(T���J�h��l�O�b��?�e&C5W�VAbA�S�6��yQ�>D�@�s玊$��:�O�\���)>O��Fz��ƄKٶ��G��'��� HJ�l7M�O��$�O��">�����O��<AC.]�Xǆ	,�	R�����'k�s
ϓc�Fl2���9-u���i��
�@�=��@[\x�8it)�<k�%����Z�C�Q̓����)�3�$ ]tX]�QOU�p�m�ݶ!`!�F�<�tI�P�^P�Y�&돀vc�ɡ�HO>er��(i4	��-�L�F1�1i](t7n���4�?����?�-O��D�OB�Ӯ/ضp{�*���ܐ1G��C,ั�,����ɾ#�(a��c	: X��DK�f�Z��\H�����\��(�Ӟk���϶�����O��$�O��D�<Y����'m�]����� Y�P�]�{��0��'�0�pf�
Ʋɡ ��; �X�h�y�K{Ӓ��<q7 �^ۛ6�'�Bʅ~�(���ʎd67��]��\���I�ϧi�4a��[�I8[2�J�/3@ƈ�M�=KD����v�O��Y�^=zS��RCd�.�R��p�'��My���Cg�
��Gh^����N%C����2������Izvj!�҂
)��u���M�&]-ll��KZ�L�i3� Ѩ��'�M� q�����O��$JEX|��!kK�Y���x��)
-����O���/�Orc��g~�R�N[����]�DI�`pkD7��I*�Z"<��D���"κ�A
�T�8���F�dL������
H���ߋI�,��nC�L!�C�}*�Y�s��N{�
tO҉v�axB %�V���9��ؒ-U�IzGm�01��p%�i,B�'�F�8����'Q��'p�	�m��P�ц�:�T<�7��&m� ��<��c�x���!�
-R v���ޮV�x��'�,�:P���"'pT@����Z� �w�-D\c�<�w�Oq��'�d�k����]#Ɲ ��	s?���
�'��(�B��L� �c&��	�O��Gz���&j9����K������҃,T�-��ɦ���ϟ���~y��'3r<�0�`E\�B�8���c�y� MI#�D�N9e*�N_[X0ϜJX�t�wm��XF�B���V�T@7��"��X���7DFrh6GÜȰ<�bO,.���CL��|�n	�勨�����៼��Q���O��ܸ�B�1.� 1K���4+�y�
�'�l-z��L�#
����x<̺�y#�>�-O`��C;O��D�OV9�u��#t^"p���S?(�@���Ohʓ�?�����P�1(b�떂�V~"�B4}��t���\ �XpQV �p<�!�_�9��ݩAF)?��c�7lCUZ���Ҡ�І��M8�iTi�O��D�Oz�Ɏq�@M�U+E���2 �1-���?	���	�=B�`�@�S�%��av����!���-�F�R�*�PU���jm�[�	��P�'��	PMe� �d�O2ʧ�
�DHp���I�1��}	�g���T���?��Ԍ�?a�y*��I8"����`�0��(x����r�>1q��[���O� -O�p ��jю?5xia�~�dգ{���¾R��Z�:t3��
�:�!��W7|�A�C���ez�
G'��Y�ax��=���R�%Q%XJb1 6�Ґlr���i���'�������'��'��	�kW2a�4��(#h,{�Nˑ4�Ƶ�<As��Hx�@��Oۍq;hTbb�S�W��O;�	�4��F�L����gr��,�@C(�zb�09���Oq��'�A�F�@�L���Ps��w7�t��'��`�d�Y��f�m鎀H�O"�Fz��I��?J����NL:a�bl��T8c'!�ԖҢ����C;�H�8ĪܳY!�AT.���4@w�N:@!�D�[��s	����A��9�'$�M�'b�,�ڰ�u�\5IA���	�'���1����G����W>B<�S��� �PZ�K��f�Dh�C�ʾ�	K'"O��1&^l��y�D�$o�TAP"O�-�bOR�T��b����vKd$3�"O����(8�H�P7OPW�٠u"O�Ub�NH�:����^rt%3�'�H*tGּˠ����A�,�v%	�'X�;�iM	FPԳ5�U�#��	�'�6��a�VZ��B抑~����'�d]�4C�^���9G���X� 1��'w>��%nցbƜ�F̊�f�Xi8�'�`0�7o��{x5���0�r���'�T�v(�9�H��`�+>4,d��'�b��g�?oDt0�a�Z0����'Np���ESbdPE�bZ�\A�'LUJ��!hh�)�".�.\�'�Ɲ�rO�:�&ta��,n�F���'_��E��1�Z1��l��:�(�z�'��DRp�O� �
x0��Ɋ"�n]��'o�����^]y�"E�-�����'?0�c&g�(R���J��;�t���'��ӄ��q���jZ<� ���]u�<)���+
5c���|؞��Rq�<)�n�t�����ʊHÌ�Uh�k�<����+Lt܌I6�@��L��w��c�<�3gE�R�y0��& Z��rc�_�<I� ��EQ�_�CB�t��FU�<)��^�n0J�Т� :�!S�P�<	���3o��	����v�F�:Sa�P�<)rˎ�8Q�n��-2���!�c�<��ل'��\Lُ�
@ �a�<I	�2���@��"[�M	���b�<� MF�%E,�����B똧f*T���Z�a�Ҫ~�щ`N)�l���N�>�A��"�.,�&�C'yEf�ȓi
^��bm\;ot.���� '5A�,��4����LʥX�}�bY��t�ظ�ON�i� bl�N|$���^#R�S��Wi��1�N;)K����j�رB!`�PD�UI��I����ȓ�<�ye$ُ�A�+ާ) j��ȓT��h�@��
[T <�,
5��(�ȓi\�t�QJ�]~, !a ���Y�ȓM}�`xBWn�������d����ȓi	(q2��!3<��EP�(H�����a�B���H�D�̗k�"|�ȓ`�Z�(�(߁�����B��r��ȓ7�<����\,j�������\���?B�����
�i��s)�*�9��>D�};WFI<s��c��E��I:L�}�`瘐0e�9B����3L�U�<1�)��Hy�����x�7/�Q�'F2xd��6F�������T�͏{�~B�	��FiB��>Ǟ���CI$P�G(�<;���	�`����FUN2XJ�@[9U�!���o$�����*E
�ס���'M�YW�'��YZ�鐧LA�4*�fN��>���O��y5�@�=M2���ڂ��#��y�� C�rwH�[��\jCFݕ��O]8@˼�лЎ�Z�:.aj��$�� ��\�+3�ybF�%�D�S���9݀Y�3"ĭ��d^�w4�dT�c̩Z���Ǣ0�+�cM�R.L�GώVh!�d	E��U� ��F:er!a�(&W֐R��M5ȸ�����O!xV��@뛶5(:�ڵ`�0"G!��Y�ʹ��C�.t���y�󤌋
�$��S�? ���"ΒeW:q[d�m±9u�'���i��I?��	^�l'�xQ��>|�t���Z�<�[>:����A�����Aظ"<!& 7�e�S�֝S@�هqp�7@', rB��;K��ԌP�v�,���m�t�@��0gˋMqO�nߴS�����C[~`�ىM���a#�j0,B�!"j=�w����3I��r��Ƀ?oHA�P��+l�Z➨�C�A��a2��E�7�<�3��>O� ����V�ޭ�Ɣ7;j�Qa]^*�J�oܠ@�B �տ(�Y�O(�BH�?�:,��$�Qxj'L��mOl��N3ń��'[��$Ľn�5�m����Sn��U+�0�R�{p9�gY�D�
ң�"to D�o�3�0?�$�ψ8����!�>x~���
	r���G�=!������a^�Ao�U����'��4��]3t�i�l��c�� w��sWO�\1p@֜R�\�kf6[-��5��q�d�+���`����(�0,6Z	p�c*Oc��-&"dRp���{�I��'��5��4&4�y��A�'�05jf6O$<�vD9;���;g�	�q��,(Z��͓C�~�q�a��[�̀�m?Y�D8E|��i8HQwMI�-�q�p��/&��b���45W����)�M7���D�Sc���$O�Y��x3 ��\�D�;1.�?�p?��VQ�2Q���,e�ް�	� ��|� L�k�F�6�D����D�FM�hȷJ>(���I6 þT�E�_;G�"�įS(,�R��t$�(���Ue?ғj{b��!���y8��&T����'��u��.8��esP)�'&��쓋��O�=�Z$��Mx�6p��B���8{��A��40$�ق��{��7mߙ\��u1���r�0�g�1���(B�� y?�������ʰ����d��������i��JX����7e`����s�i��c�pQ�	&�Oj*�D/�N]�S��g'8k�ր�azr욓S�����w����)�	JH����^Nl�H�P.����ϡt*���'�A5����V�Cz�� �R ��'�$	����4���b��*�L�M<I���ץN4"#��i��p!  �I�w� J������(�F���*;}bI�S���:��Λ>kV�
/l�I2��S;��nňPp�y"�B-2d|Ȉ�O�r4��,Q�yb*� GΗ�}�m#�I��M��ɍ$L�*J�569�ai��		V�"B�e��9Z�$��H�q� l׷<��Sb�I�,",J�a�_V���;/J@����4�c�!�\�lk
�L�ج�lK3e��(*�Fo(]a�\>⬝r��@J~�*�l��X9��T@�b����OФ��ȗkk�|0u��5�Nii5�I��RqPc�ەq�.�xBʛ�'��yP`���#�^��ȁ)VsN���/�H�1�|�:VI
;��� aPc��EZ��W�#5�����8H��3�ND��:L���S��"Bn�W��L�R���MZa�<1C&"=��b3��'@��P��s� �G�>!�;��) v3�} �	O��XϓE�*��S�^�gp4� ���u������O*��A�U0�^4��&!��m�$�
^LL���Uza6�ζ"ay���;,] j@hO&Y�X,�󡈺�0<�!@!�"��jѼO��|���6\���'�;JT�\"!FM��P�O�2tHK�`�����
MN7n�[嘟LI��xn�³��h�Dcӱ�R/-1��q���Q��%�g)��yr�4�ص!���`�>8!��կyG�'>9#��ŏ9Ǟ(B�M;Rɨ`�yrII�-�N!�`D�L�ZlAƆ���hO�|d
�WN��(��Vې�c���eɶ��'  �=���d�0t$�����;� ��'i�>
��|@2�B�qF�S�50�u�3�]��?�1*Ec�.���I'zc��H^+B�sB�C�5��i>���CM�R��Y�EIu\�9`��h�<�ą]4a;�P@��8nMlpa%d����D��ELH��R���4��)`FJ�">��6Hrޕ��!W� Q�y�)�x��)A�.�O��i��O�]b�a����a��dM����|}RO(+�F��$c�el�@���L��(O�d1��Z�pO\�q.�h"8E��I�"Q@�V(�eF���)�(��k���\(�u�Tvp���eC��R�X�ʁ��.'N�cO9�Ok�$
3'@������,�� �'F�3�dO�eb��S��B�M i�,g������<ͻ�N��c%N&_
	!5C[���Ȅ�x����kF��@1@�F�-`Z�D����L<fe{5!P��@�O�.ˋQ�� #�mݢ�8yF8{�!8w�ܩ"��P�m�����Q�i�ӗa��=%�I��X�r����Ҁ�+�v��'evdSA��k�z�r���iz"�c 7�"���LP�V%��ѩ����OpLC`f_�מ(բ��q�:R �@��}sv��V"`D�&o\#-�������'��}b!
V)r���� ��6t#�
N�{f(T�ԧΏ�qO�p�W��!� 5�����b�1G���� �	��j�=l�B1�Gř9%fH�I�"O�����T�i{�C�?x(�q ,�B�	��������=Q��9�^��צ��&�U�� 1=��"��'���姝����isl��Zh5����n	��'5�h��׳o\	��2t��p�r�٢$�܅(�%��� ���'	���O$�&T1m�TDR`4}� ���ia�Ÿ�j�[��-RD ��L�QH�N�+/���c�����dϊ)Fd��$�D� ri��k��'��2E��CWB�[5͘�v$���{b$,hFAdf����T�!�D]�ݘ�x��Q�5� %ٵ�X�j���ԅ�g/�7C���S�iǎ#٪d̻dx�ء�ڻ���"$��,'���ēr�@��R���;b�A�ǉխE��D�Œ�����p�"�R��q�qO<� @!	W�;y�~Yz��E0���I�r���	���p)��d�%D(�Q8�Hߠ{=^���Ź*�����W ��ę?/t!�� �ʔ1��_��I;C�>	*W�X*>� �p��[G՘�s��B̧P��|q6&��C�l���<���ȓ�2e#��ׇ4��$�b� v��i%BF�n|HG�Yk.�S��yG]I��R��ńW7v�kq�6�y2b�QT�;#�CG��孊�yB-��wʮ�st�L�V�Y��ɽ{���Ц��r����q&ą�x�<�7�ƿ��4�ޥ�tg�;d4[��T�9y�H�)o �e�AFXB�I��I�� �T�a��.Kh4a h��5(0�'Ն�*ƸiR֡�d+Qn���BU�RoWy��# �=L�Ɓ��"OJ	�6C� $< �A������&�i�v�����Mӧ���I�Mcw���4�8�h���=h�T�� L�0�� ��4���b0O^ q$��K,h��@Q�P{xA��"On�Z��]�%�$L��˙Wdpy���J�L���i�:2���1��۩]s�m�O���!��ԓ)NlBB��Dd���׎��n!�d	� ���EЬRG���Q�B;=!�C:a#dlX��Y�CX;c!��>"P0͉&Ĥ^��$)�́�
�!��gBT)5l�:�:<KtO+a�!�\M��bf�G��s���]�!�Ĕ�P���z$#�&m�m���b�!��߷w�Xy��0l��@3G��4�!�DK48M��2���~��=�'�ՌK!��I-L���`��?e��È �T!�d[$�t5�f��F��K�ߗk!�^�l���r�̥-U t��>�!��*�iIb$T�P�1�O�^�!��^1:�4�3�Z3� a�5hA�`�!�D��t�Zw)A�`�8 �����+�!�Y�@�Ti���9��4@���4j�!�D�Q�@���LY��� K�5�!��|�h�e�ݐW��Yq	Y�)z!�L/�D��u��O��m���-$!���
D. A�"/����^�
�!��x�t{Pe�#v:�u�C�G�!�$��4�Ƥ�$���z=R�!�!�Ěi��ФdH0~�Z\(4�Ϩ�!�d�<�M!�*�{��)4�-�!�$[a �y'�Z�f���(���!��Z��A�iP�GGd(�4GX�s�!�ă�.�����X�fG�Li�� 5.�!�$K�^�����׊36=a�g�%�!�."M��'A��/�H��0G�Uz!�$�E�nM��X�d�*�Sg�.E!�D΀Dǆh����?z�Z�x��I�j�!�϶ L�bC1��}#�C�"n�!�ą�M	�:bd�$eM΅��/ޤL�!���Y�lq#���hR�(�I(G}!�dޑ��!�-42�|k�ǎ�^!�d.� �32
St�L��bx�!�y���#"6u<q� (�� �!�� ��o�k�Ќ��#R�Wjαi�"O���$��(q��v"^��-zT"Ot��ƱT4 B�NЛX��̓2"O� �D�5:����)(�d蓖"O�5�2�7b�Fi��dN8�ě4"O���Si�q ���m1�`�"O@x3�D8SnN��R#�	��p"Oh�(D�O�wII^��p=��"OhTɴ��W�,�)�׀�6);�"O�M� ��4Ӹ��R-�M��"O���G�@�Z¼ƠΨv��%�$"O!z�nؿR%�����7���g"O�+YukN�����<,P*'�Y�<�F([�4�ᵌI�)l2�IV�<Y���8��MAmʄr��1��S�<���7]��B@
%�Aq���u�<9$��3 zU;�C!�jd	�c	u�<����r,ъT�;s�49��^t�<IVK�:> z,��^�S�|m�sHHm�<�7��;J�"%Z7a��kp��Z��^�<� ��#Z|���	�]����gc�<Q�n�.|���D�wd��i�<A'����s��ʢ{f����B�d�<�S�ʮ4T<+)*~=! _�<�Ve�)�0����m��وRD�t�<I�bӷ_����&GJ�a_����BXt�<16�ғ�b�GG�M��D"AZX�<Q��;44�Qj�+ܾv�6�I�aQU�<1G"�X� �jCf�8/4�!�`�Q�<�ņ�#(�.�u�L6?#Z!� i�V�<����ߘI�SeM�!R� �M�<��h�r�)W�@ ��J�s�<��OZl�:�qV
���1�jr�<���2g�b]hF�< ��	iW͉d�<Y1jG�d��i�5��2mٴ�I�aAa�<����#@���G��\�!�R�d�<��.@#|c��K"*
�r A�tN�d�<!��́y�$I��ރk	� ����]�<��	YV�xq6�[�u� �~�<Yր6I
H������5���PCev�<����PH��^"!.��'��r�<qTDC�x�� ��R�Rl3F�l�<i���ݤ�2��)(���0�g�<YbOD?V3Ҁ����+
	�=;E�i�<�!�:`8�U�g%ѧ<^0mz6�Va�<ysMO�(
YC�� �D�]�<�C,�ʩs6��" 1h#�HW�<q3�	�qRx2č�c����Dd�k�<�ޅ]̀a�@m���2���Mf�<�U �?+��[FHC�\�8숷�`�<���'�80����+x�lYrvK�A�<�V�"
mЙ�7Ǟ%M�\k%�AV�<Q2��-[Հ�û6��	�e��R�<�F�Y�.!�`M�5X����LO�<A�+(8�0쫱��W����<T��q�ļ.�`�F�"=eTԊǂ(D�4��)A��i3/	�| ��Fe+D�H�V	5jr0�+$F�Mj�a�5D�(xb	9)��h�@��yjs/D��0�׈|�����>x�< �+D�$�5j��\f�tI�J>Z��h��E<D���4bߕw�@I���D�#�:D�0��A�{�"�(Ab�T���CQ�-D�@��F�v�3��O�	*���!)D�� ��*��uh��@5Gx�<�y�"Od��!����)Q��-S�8��E"O���ł���Lp��Ġ
�v���"OT�+���>�H�f�T#G�ؼ��"O2b���/X��`�$��3sH]��"Orh��]� ��äh�	$fiH�"O��h�&�'D�� �&ha:��"O������:
(`�R%9X��qU"O���G��b�N���-j>�d!P"O ms���.#���`�H EFJ���"O����7���r�9��1� "O`-z��[:(F�<{�d�!�R�;�"O�,ђ&�#;� �QS!�3l���x�"OL���lQ�R�a#fU�>0{���n�O`���iH�Pwf�K�e�4Z0����' V@�W�ܥ1hL�i�@�fy
�'�v�x`(�x��1��Ȝ�7���A�'��Y�g�8)X`���%������$5<O�ᠧI�,�Q7�o��͒&�i�ў"~n�<�ЂCo`}��̞1<B���j�K�ih ����3�VB�I�k
�R���"7 *YzC�I��z�;�Z���U��B�	�UP� ��"�?YݮM��cO�|	,B䉊Sz�j�B7J�9Q�LL"q��B��)� uh��Ǉp��\�$ V�>�B�	�4պ�N��j��u"�7]jB䉾Fy4=:B⑛.>u9v�ؒh�jB�	;vGB�)W�*a#&M��(��Q�DB��#+ 
�x�ۂ]�x���Դ@6B�ɿC�PQs��R�T �	P��c�tB��"
"h�סZ"]H:r�R9 �.C�I,=ג��e��Og�D[vio�C�)g����bU5]�����M�B�ɻ*Ӝ�d�4	�, !�-J1'W�B�
9L �a��j�.بW��"FXB��/#������Ϩwmލ9a�g�2B�ɓ)0ĵ�	��{]�Y�I	4]�B�ɲ'84��O�z��)�ƕ&�B䉠!�4t�a��!9a<@���@�C䉰���iP���`��
(��;��C�0f�d1��
W�Qp`n_N��C�I�4��C ��"w��E�"7��C�I�$FX���+�.w��w/ۤ&�nC�	�T� �� K�7[��!��&\\�C䉙>@H����;�q����C�<b�L��-� �FD�&HҿǰC��<L"�1�ݘq6Fp���Ny!tC�	0 �[4d?�~�����rC�ɼɺ���_4Y^=�U�)2Z�B�ɰx��܋A�!k�v%#t�J*ŘB䉩n
�hb�I�6|U���(7XB�	�x� P��G��eq.mY��S�zC�	�z���ǣH>Hh���X����6������a� e����᎐;т$�ȓ>2�K	"+��L�33p���S��)����;���Ə7LaL���:I85TbK�����K	V�`Є�� �΂�>E�ghZz0�Ʉȓ\��dX��\=�,�¡DZ�Pٖ���yGR�H�+��~W�Eq�R�\j�Q�ȓ_��1P��7�za�ɜ.�P�ȓ#8n�����qV�� �S�H����<�G��9�n)�"�ۧ'zu��S�? .�Ɂ"'ਙP�H0~�*��w8O�=E�4���"�  8�I&n�Vda���y���)+�iH�#��im:�C������"�O�m�'ʅ,y��|R3jW
c+��ʖ�'��#<��BU)#�-"D�'�H��1��a�<Qc�*M���bg���Ԍ����]�'{Q?�q�$ĚN����Ȕo��c��-D��P�ě"w��G,LI�YI� -D�2Fg��ɞ]bt�E�	���@GL%4�����S\]���3e��y��Om�<S+�k򼹤߈
W��
��]�<97�ĩ��͒���	*���bAS[�<�����^��`!� H�s�Z�	�F[Y�<�gI51�ʌ*B�� _�flyvKNV�<q�%
b�4S��:_>H1��n�<��,��h����(�F��@��g�<�p	_-E48=�c�M�P���GK��!��� .�x5Ȳ���+T���V&�!��,�eqW��Xp0xXČ�9s�!�дTQV-�f��%Z�43��,e���hO���4/έ82I%��)��y��"O�	�G�+^�ذ2bC��a"O�5�fD�v���*��ZĚ��$鉤e��?q�L#[�!��R�l�x�I�` D���vaY7h�vek�"��K�@�@��O�Y�����24a8U��[���)��OG�8?�y����@�G��_������;5����'��}�F�7^��ܣל����N��y�V!f��A�AcB�ېAsE��*�yR��!w�6���M8ŖX��Ǟ1�yb�#d�FI�`薱Z���yB07��d�D.M����L���y���a%6��b�{���eE�.�y�άn��Iʅ 7��|0&�&�y��Bۼ00p�2�.��d,��y҅S"~ִ,�gڽ1�&1r��P��y�m��k�dUٵ	�'���;�V��y^�H��yy�U�$��h� �y����_�_ .�q၇� ͚1[�'� �uE֥bT�E[��A4����'��E�7��0��]�dS�6(��Y�'�e���&(�4�q�65��U�	�'N��{B��*WD%g&A<KC��7�"  ���{�0)�6�نQ��B�I<HQ� 2�	
���"4��B䉉b��K���p$��0Y���B���εS�,d�]���A�;_�B�I
W���
'X�RM�,0���Z��B�I�|�}XA�t��P���A�*B�-	7�p�!!Uz
`����.O�B�	�v���iŬ	� ��qSaJ(nB�I&���QjG��� �4F̦B䉫ך�V��:J	��0�@V-l�,B�	�=o�]��N���m�JO��B�I9/��������T! ��C�;"غ���Ȃ�q����l���C�I>�|`�*K��K��3f~tC�GŐ離̍z���[Q��M�ZC�+$��QU�H�m	`=T�BNJC䉑q�>-�ѫ�/�`؀S��X C䉄����\
�s!�̰b��B�ɹ ����<"���5e�7)L�B�I�:)�AY!H͵R
��ҬɃ[|B�I�,:��%%nI��Fț�bB�)� 2� �#A��P��l)W�m�s"OT�P��+*n0��jT}p��e"O�LaA��<����aI�Hmc"O��{T���u��dhB��[J��Q�"OH9��-Ђ ����`hķn.��aq"O�1W/ߍQ}�)�2xqd"O��s&��$4%�q�� ٨Bu�՛"OP�����X�O3]=�!�b"O�ՊW�Hz������4L�"O^x �Gǘ��S�DA�\��	D"OHȢ��
XM�i��3h�$"Od`
�+̓O:并�R*nWvD��"O���4�
�G��Q'�ҐMA�@Qt"O�����;Q`�(E�&|�%"O^�*R��4|pb�ص-\�s�RQ+�"O�IY%Vg5@��"o�P����"O�T�B.� TÖ��pD��|I�T"O*�J�H]�
0�Y�CH��<��"O�`�fʴl��͹shBa��%@�"Oz���ʄ!U�z�z�&7���ɦ"OR����B��j��٭1�vm�a"O�p2�	�0�<- �E�~�^xW"O��3�#/A�iCJ�%Hȣ�"O�0[��j����h�u�p�Je"O΀��Kz_<t1E��Pv�is"O.�V����A$.V�=�l1!"O<����;Q }��k�d"O,!��D�'x<+E��`��8�"O����9T��5��N֒)x!�"O�5�c�X1�\�w-�"w Fa�4"O� 1 D�-.�� M��6��|��"O�Aa��R 8Z�
6�q��"O\��BGǥ9ʥ�U`�$"�I�A"O�X�1G�bn����h"��"O�m���W�x��k!��kfܩ��'Hda�׈ݷle�L�Q,�91�̱��'�9H�N�-*_�P�ƃ�(�:H��'�T�6�§ �j%2s�O>#��Y�	�'��A��³K�dX[����غ�'NX8��C7\�"���ͅ���mx�'>����#�<AѠ�$�QY�'����O�k�UALDz2x��'�p�#�H�d$�S�O��}2�'������h�>���R.(�a �'  � ��SN�s�Q�yHZ� 	�'��7c�#jenI�RN
�tۦ��'IvD�%�9JZ0�j�#.	�'x�]��%��f��G% �&y��'>r����A�qyh��U�9-�9��',ܻ��'QS�`�"��#��X��'XTQ��GS�5���D�M� tY�'����r6�R�JRL 'K����'�*�(�NB�6q[��E�xK^T�	�'�-�'@@=V�ç��<kϢ���'jB���F�~p�E���đd�F��'���H��|�̠C$�@�o`��h�'[T8�0��;$4|ы����1Z�'AT35��.���I�e����@�
�'P=��3C2șH��5
MV�
�'A|�`��̆i2�)xЬZ��2���'Ċ)iBBP�v�ч���\�}��'.0|q�A�"�6�	�A� zql�'�&M�v�ҥ{�����y�Pr�'��5z�r59F���v������� �Lbb��%X&���<�t��"O�K�n�p����9d.��
�"OT��®ެf�j��E��3fBYH"O�!rN*o�F�2�N�DSzA�"Ox+�,��r�Ґ���
 C4e�c"O�����W0a�
<!E#[�$&�4��"O\`��O�C	��g��JLp0"O�%Q ��Z��ibVa���|�a"O��0҃�VE@����ʶ�j�J�"O���⣀F��1�b��!H��H�"OZ#��Ȳb��b��#a4qj�"Of�b�72vQ1�HGȀq"OV� C�1Ț �w�X� @�Y��'L�|rQ!M���M�c���
�'9��J�k>2p�����ZƠ�'� -��<jG�]���QN���C�'�,��>e�"�	��ӌFp��	�'��	��L� '"����/��>��͠
�'�Z(v+V�N&�a�c�4m��
�'����g�,<F��$��;b0����'`��h��*@.���[�1��(	�'N���	��0����R�G��	�'��t���u�r!��$9.��0	�'�H}"��)�L�`��Ρ4bތ��'h��e�N�H٪T����-dQ��'T*��T ��
�!qG&�"�����',����[�`.�ٓ��E�8lZ
�'F60S�	
�A1�ԡ�ԈDZ.��	�'��]�5f�"�@B�חl��5��'���ba�?*����MN��@  �'��@�r��>nF,S��N7����'�����!@nּbsn��VX�	�'9R���ₗ3��ZS`�>�2���'sf�{5���i8��Is�TuPl�
�'�������\����`�T�	�'�` �!g�*;�
a�jY�R���	�'�
m�$A�l�l�j�ʌ/ք���'��4[t�ҹ`z�9����*0H��'��ұ��9%e^�+qJ���l��'��P�Q��܃�c��V ����'5���Q���=֊x����"S����'���I���B�nB�;�<��'!`�ģ�T�跥W4�܁��'����/Ղ��8H$�Z��(��'�(�v�
�ΉѦB�$|$��i�'�V�yBC���R�16,�y�H�s�'�p)y4F�6ew�3$Q&n��*	�'�0�@F�S+6e8T�S���pG*Lz�'�rU�enն>A����懐u����'�f9�l��
�4,#�-�^μ�	�'Jv��`c��(�`�:�d��3�'��န�4�!b㋫og�d`�'|�1@j��y[�8{q 
�����'^r�`�2wj72�V] !����y���1X�d%����A�L�I���/�y��8)!w��4p*�V�8�y�L-t,��,6�e:H��y"D�02A@��W� XV9b�k�?�y�T*��r��M<|��@�0G��ybL��l.���"y|��c`���y₀3@�m!�ʧl .5���S"�y���.~S`�ˤn	�_�4%R�A��y�[S�D)s)�*U-�$2�H��y�D�*�0M��S��ܡ��Z9�y
� D��kRi9v j�/�[���2c"O>D�v�S	=�:�ʐ��4��"O�����J� m�@���Q�m�d�"O�P��I2-��1%e�$UŪu�"OX���b:�����2-GT��"O�͢U"�=u���+!H0E�p�g"O��`�
Ԕ "�����"O�9"���E���:��(�V᠁"O[�U�F�v�B�h劓9`8��@"O�8	ڎ���	U�#4�M�f"O�pЯ�y7�]��(W�F�sB"Of��%Iٗ:�ش�SŃ�shI8�"Oѡ��-h(A�$��S%^93"O�kU�I/6�98�mXvD�
V"O ���m�=��H�C�&�t���"O�	vH��y� ��G �u�D�G"Onx ���7�t[-I�jp�ۇ"O��$�_Y���I�F[�( �"O8�d�������7�v�@ ��"Or0��B:~�PqU)��c�J�r'"O���4�O�����ˆ?l-S�"O�M��cԴ~}��
���# �ʸ�"O� 3AÖn�N��� �P�
 p�"O��Vk������Q'�9�t��"O�K��̿9z�)�k!NX�l�Q"O�b�� g=vJ���U�1�"O2��QB�J,cTD
..��	�q"O�|����-ur�l�P��X�ux2"O樂a�ޥb�h�ӣ�5dH���`"O�1a/C�$i�y �BE�C�P��4"O��S�"�
+��3��ДO�|X�"O���A�إa���is�
�G�j9��"Ob���1O=���.^�[t����"O�+�
�[9*�a��6��-�"O�&N�M�VM+�,J7F^�ś�"O ���
��U! ����P�=���"O�����;%��;�c��.��u6"OLԍ�>l=v���#���~�YT"OJr҃B�{Bn���O�[�\� "OJ��U(��?s�����ld�"O���@NKĂ<�u��	hM�#"O��p���e2�EV�_����"O��s���9�B����#@t�"OhU"�lA����7ꁡo�*��E"O�PP�ʕ�.�!E�Ew�9#f"O��PG���V���Dآ�r�Z%"O칐`��\;eˀdl�̫#"O(@�� �*A�mR�bǧSb��iD"O`�B�5��	��_8`O���"O�ॆ@	n�5K��f�N��"O��x�L!#Ǫ	&��"�6@"OZa��.ͽ �iC�gU�E�*��6"OL�:�B�0ay�s,������"OT%8%�	�u���Q�WD�z&"O~����<f��k�䌭P:�"O�A��D�<�Paz�O�e(���"OZx`$���l�@�K��H�T�3"O�i��8� )��b�*c�b8C�"O��Ѓ(O�2�X���[�x�r�)a"Ov��7&U!6@�3"�FV�~��a"O�|HjQ.����G8W�xܳ�"O�����X~"�q��٘w�X��"O��s a�J��tjc^k�N98a"O0���c�)x?`;1ኰ%��<��"O� T��T�C�7$�"�/RG�*ܫ�"OV��g��@��zP�3��i�"O���x��X�P�tu0��"O�Q�!ON.9Q�BG86ь�{�'[�H,s��L��@�4���'`ș��aK�Y��ʒ$A��j(*	�'4�`*��_o�l�Qw&���z�)	�'��X����j8�a�1+@8a>~���',ୀM58���k�nI�\�& �'"�����D5�����	�~���'���ѦL
}!�P��
L���	�'D��\w� ٘b���m~`A8�'��A	�Ǜ7p�F�1��{�l��'O:4�����8j��ޤx!^Xh�')�ۤ#]�SK���5ɾ�P�'Y�aa�	=n�×	kJX���)��`X�M�\l��.^�DS��y"������	��C�,��W��y����]:���SZ0����5K��yb��]P���FBˆ=��0ֈ%�y�.�6@�D�Y���9*(�425�Q��yF�;|ud��Pщ'a��B\��y�Q	\|�:� ���P�船�!�d��L���eK߬�8t�wb[>����%F�s��NH�4�uD���ya�G0(���&�5JG�y��?$h�H���4 ������й�y"/�9j�SE�	�K6���ՋR0�y��7J�@;6#G09݂i�Do��y��A#y�		�d\�4G|,�����y��-0��AS5₇5O.5����yR$�2����$E�A��!b�nT��y�va��i�͐�16�lkG�M�y�C�(���bM�0����FIѲ�yb���]�;p���&:Fi�V!���yb�޵��S�B���pp�4�y	�4�(-To���v���]	��D�<����'r�I<3�<�2!ޏR�<ig�?^��C��1@޼��1��/@��8���3b��C�	�1��8"F3$�N܃
G�Y��B�	�W_�D��E�xj24)�i��4�vB�	�@�<�ɶ�G�^�0�(&K%��C�	�wl�u����Of-�f�JF��C䉭V�����4Zj�* 		\�C�I�'��%{�j�oPA���ƲcthB�	�\%q��֑2�W�R�I
�B�	�V?���dԬF:X2v�N���B�	�H�,�
�	��x2E�>'D�B䉓$�&-�� �t�Jy��"
m��C�i%�2��-g�^ 2G R���
�'d �Q�	W�*ξ$#W�И<�#�'�@e�0�U�(Ҍ�����(����ȓMV qaǄSE����_\J8q�ȓ��9qծ�<���q��I:R��ȓ/C�ݚQ��lr�k��̇�R=�ȓ>��
�C����=;���>�� ����-ҥ�£_��e��D���e�l�r�:O�iw�׎V���&�\��	<z`l��J-}(@�4��_v6C�	/?�~��cýq9D��B�Z�"pB�I<�Y�Ǆ�#�<�8q#U�-�xB�I)Y}�\z�j�*���C��`B�Ɇ���(�0:C�l!�͊2.B�	 ��ʓ�g�r�	 Oς-�C�)� f}�ף�U�|L"(�f����"O�؋��"F�ŉ�$L:|�Q��"OD�sC��X���yC�5C��1��"O���w�E(k���6�� b�N@��"O��ЖΘ�}�Ƙ���d�aU"Ov��*F)��[��.+f� �"O,�3͆2RH�p���2ֈI�"O�=�� &"�I��-�p#��[��|�'x�Oq�F�Wǝ�%ox�Y��ܬ�"O����JK�z���P@�%*��z�"O,���$�^Ԙ�:�o�4֡�R"O*��A��.���{�N`I�"O����m�$,���
���:(��+c"O:���	ԗ2�z@��,ϻS���`"O��;����l~�D��nN�r�����p��B6�Q�y�ڍZ�֊��P%x�!�$%S����p �3V���kV�*�!���tC��#G(���hp�K7H�!�DA#"_̰&�R�i0���<3!�$L,V�z�k ���)Bi�����u{Qk�)���g��aw�ȓ"O2,��%���*�����M�I{���������
h2R�٢�H,G����-D� RU��^Ă�C�dE.27�����-D�$�e�R	󀍂e�>f�3� D�䣖�.
(L�� ��~�@|j�h?D���0�R�dGr���)Ih���<D�|�&kÑ'�h�r��$#�|���:D��&���QߘU��ҿBS`)�'�8D���u��:c��sOքY�8�2v+D�0��T2"��D�wDӆ"���Q�!)D�����؂$��,8�3r�����;D�L��(�z>�� �X$rF��X&@-D��zf��K�����Y'~(rMbR+)D��`���%uRp�!�<+�6���	&D��S�==�M+d�W�Q3��."D�"`�K�C�� #F3S������>D�`Agʈ�z�ƣ�*r��pS9D�(��>o�8Pb)&Q�	0%1D�DP��(^Ʈ�"ro�P�����C9D�`x�ń�J�Js ]�wbn�a�$7D�h{����1�a���^�6d�S��:D�H��� }Ͷ�q�gZ�'�,�y�o�O�C�ɾ]��ak6��9<ۼ�����9+�XC䉁4��yt�z�ٸ���)$`B�'rn�H$
݃G�:����WBB��-9� @�%��>uN����Ik'
B�ɬy}`��Ĉ^��Ri	�h�C�ɈR��0f
�$�T��"C�&cRC�ɥ+/�ڀ��Z���)A�^@rB�I?{l����U���- "n�B�	蒑��+.�&Y�#�4W�F̐"Ob��)�"7�&<RdA@�6��-	"OĨ3)
�vh<����#-o
(s"O�	T+'�9��K@ND[�"O (�dؽe�(�9�('el�&"O�;�`��:�ּ�'�'z��l�P"OL���L�~��y�&�$l�j�:�"OD[��Ag��Dң��+n
��W"O,���i�o�Q�d @�%����&"O��;ԣK����=e�F�8T"O: ��T�y���œ?p�`"O�(;�M(a��j� @��"��"��`�Oh�����"�#��Z�!�mc��� 8a8W ��_�����'�-"O�C�d��c�Y�#�в_&�q�""OPA��2bEP�,�;fp>��"O���E�K0.�Șa�ch�A �"O8�"���� �j��f�\��"O�)�˅ k" )�b@�^�HI��'�ў"~��-т�9P����|,��B��yR@G�I+��Vj�)j�.>פІȓ(T�qE���mJ����J3*����`�d,~=�h�MA�7Ū܇�g�j��t]{\\駬G�n�T��>�ȲЬ�"Tf�0��� ����ȓU���&���;���|!�d�Iy2�)ʧ'��axŦK(X8�JD�Ó=V����l�h1kC���x&��� �|8��ȓbH<�rN @'� i�J�L8栄ȓ/
~�+�cU�|)����Rqh�ȓn׺���eT�bc�Q�I5X���~g�1�.�ș��L�?I:t4�ȓ6�&m��2FN܊�*��N�콰���.�	d~�튡rQ~��/P��
ǥթ�yB₴r��#�P��a#���y2j�bd��D�3��9�$E:�y� �	\�� ��.B���+��>��O��w$�p
��ƪ�0Pͫ�"Ox�t$|��#Hx�����kr!�D=vbSk;��9�b�%:���zybT�4E{bg	�C��㴣Ύ}KD�����!��R�6�"E����%Aư��K�a!�'�Ub�Q�:͘���
Ac!�Fq��e�2e��`���|]!�d�3������
4\�q�pk͟5;!��'�tP@���R���"�LY<!��#@�0@Ӯ�@/����+�2R!�Ę7w������EIȬ���'�!�ۃ���ɲ��_Xd��$�39�!�dM�f�y,P;FK��HD�{c!�նD���:�HK
3��q�knL!��B] >���e��5�4��;p5!��G&tZ�8�W$/4�F$���3t!�D� 	�@Hw	�����g�[�J�!�� l�-�#��s�A��B��j�!���vDD�*��Y������q�!���Қy�'F��B�M0�H�=�!�D�3-�&#����W���_�!��b����w�L�^5�(�:!�	�#��xXA��!U����*�A�!�$^2|}Dؘ��H�ctp�5��^�!�Iq�$�%J�����K�ae"Ov�P�����4�G�ro`䪦"O���A�X�a^�js�Ƣ��qy0"ORQ��а����,/�� ��"OjhB# �( Bl,�CN��A�H�"O*p�ϡLU��80n"+�VŠ"O�<�P&B�#`��j�͖���y�	��

^��'JF�e!F�� N��y�%ܯ3 �8J�GF(d���*`NX4�yrj�6�������>Y��T!�@K��yr�&.�=���YU�0�gN�&�yr������P7�T�4�D�y��`<�� C��zB%�cfT��yңA`&δ��,P
s�XQ�0CQ�y�n�RϠ�"vo]$Ơ�X�d���y-D�C����e{a�]��dJ�y
� `�B�\�0�:!r�n�M�y#e"O*��6���d��(B?��R�"O���!�0;nL���g5x�ȓf�T)�"H�Yw���Q m �y��g|��C%)��)䜪a��xP�����ܟ���� ��i�ĥ֚4ޘ�!`��N�<!5c-/\�9#c�7�84	��H�<�g��F��8��.6O�A�%�|�<I��ϝ����c�+pf֘�
x�<�s
h�dnn�D�a!u�<j+�8@��.� j�d%� ��Z�<1���X�7�S�b��\�$�_�<�b`J�h8"��wK�� ��53�f�B�<�f�!G�U�k��1�� Á�{�<�"�tlT�%�׌-£�{�<A�n��D��1�Hu�4��1)�O�<i��-�X��R��)��fdM�<QuaM��j�l�R"�S1�BF�<i`�,~��VኗoĞYibb�'�ax!��`a�ĦD�"����aO��?��'�����%|��a�fɂc\<=c�'�
��� �ʁR�^ǂ��
�'֡y���R�&%+&O
�l�@�	�'4>p`��Ґ)y��V��2|��0�'����IJ�z�d �5ƨx�$*�'�`��>%��$���A�mW��(M>�	�'w
�����n�����Lهȓ6��L�M�&j� Hs$!��%�ȓk��,9�o��^Wh�ā\a�8���Q����C)�:X��		%+Z�$��@r�I�!�^�PQ��ӱ���rA$���~�"��'S>�J�#�!J$Tf���z���둚NeJe�S�O����IQ�'�L��7-�)�!!T튰#�F���'��� a�+�ҹY������L8�'C<)c��_2p02�B\�����
�'y`�Kv�p�B��b!�'D�4��MŪFrr 2�j�+��
�'Iz�R��N�K�l�k2�X�
�Bt;
�'��e(���9=ل8�$ҁ���ߓ�'�HȨf�1	�Xa���cM���'�aA�Õ?��0u�ғ.��`b�'>F�8��/ �l �D\(9͋
�'�J�	�3=�^d��e&�
��	�'��H#$�ݏ7޺��'�#���	�'k�9XV��9:��s$�W�F���b	�'�4(�fk�1uwf9pM�8����'�jQZ7��;(�B�(B9` |�j�'��`�Wk;�غqFǂQ��
�'������(�l� A�ǳv��8��'AT��0���l*0AB�}^e��'�����D�2��
��)<�!��'���w�	-g�|p�g������i�'Ypm1�$�= >�\�"@��:���'L�	��K��m�:���R�v>l`�'�dt�d�_��2kA�@;kfά[�'�6bF#+6� �E �=����~>�0�lS�o��b�ȃdb�ȓ6ȼ���h�l��4�����D�@���^E����`��Y�1�+޾bX�h�ȓq��C�R0`�~�c�͔�T��H�'�"�)�ӚY���ap�ުXb�ٛ�fQ5���0��z5`�%� 	���
�UH<D��a7�S1��,0ӥ-!�@�R!�'D�� �q��׶5s
��F�D�A~� �D"O�(B7��٘9{�%�]m���"O
u�E��+s ����=A����"OA���i�d���̌�U�0���'�� �a�O�mN�٣��BM�qc�,D��֭]5wrș�e�L���e$&D�0P!&��	
b5�WDہi�lB4M#D�����23{0��I�1��x�T�?��Ԉ���c��9F�*qK��_%N\����"O�dA4OA�_��� �i�FEnш�"O�A0V�3�Uz���,45��zWX�4��`�S�O(p��|�p	�:"����'ɂ�SdE�{�y���k{ �+�'��"U���Z��r�^�H�x�',ܩI#H
"4l��p�ͻ�+
ϓ�O��i��4d>�p�V+=(�� ��"O�S��<T���k�)L�:��tP�"O���������jVnԚ�bXY�"O��R���9���q��;(W�Lٴ"O8���O�Y�ZY�c��"C�F�J�"O�p��h��>!⫀Z����"Ol1���6[˶�����<C����q"O�mЫX��]ү�7P�Yd"O���
	��5N�D��u�!"O�`WE�ϒ���y���b�.�y��P$>
�+w�P7#�Ipb)!�yB���XX�`�����b���IE �yd��H���ɣA�3��53a�W��hO���dT"26(��`AB1̀C�^�!�ȖA+�L�-� _vMJP��%/�!�DO]��8�b
P;H�^P W	�+>�!�$'F���g�+G7z���ˢT�џ�D���m"�as�&�9�ެ�v�X��y,^��fΉ�H!bD��y�M�/;�ش��l�h������y"��$UG�(�7�ltF� ���2�yҡ��]lA�VgǨ`ZL����3�yR�ҙ5$��&FC8f]z��2ş�y�j�/nl0;ŦسbX ��½�hOD˓������jT��D�G2ٸ�"O Q	AEO�,�K@,�;�8��2"Oz�cB�*uv��	�Q��1Z�"O^�	��c��yS���Q��!q"O��@��!�x' �O�<��"Opu!ǒ��t`{r��([/>uKD"O�d��O�8_5ҝ��A�H��@ht�	�X�	V�O`(�4�N�%��W�9o����'��(�!/ XЁ��I��\�$���'L%��.Vx����B�� Sz*$s��hO�6�
�4���޳a	�]hT��?#❇�8(BU��Cȕ>���h3j>3�(�ȓV���Qe��~�vL+��	�x$�ȇȓ<��M�>ƒP3c��W�($�ȓ,e^���1 =q�@Z�8�1��@H~XɌ�c��0�&�^�jtR4��7b����X�<P�HU�D�p�G��S�{K����A�m���`��C䉪!�t�D��-i��n�7��C䉓3����� ��k�@�:=��C�	QG����-�jn���OY�ҦC�sp�@��-5�]��X?�C�		+����"@��I�0��O "C�I�hj�B�-�,�����5&a��=iÓ���fЉD��<!uL�  ���S�? b���&^����b�N�p{��v"O �Qf��jG�A#�↣`lN���"O�)�&ާ�<������Y���"O�|" AE;a������;U���@"O���d�.V�Mj&-�K>�px�"O&�����]d� ��1|;�)z�"Or5�ՊVl�P�FJ��
L��"O�E�T��^��0�+_v�ź�"O��$*!��h�A�=0��{�"O��C
�]n�)�Em^	m!�� �"O@H���<Kw-�J��Ey��c"O�,ᐦU�[�4ti$��3B��H��"O|�G�V�GļDB�!��3�"�c�"O$�	B-�"C��
!��2t��$"OZ8S��)s~�<r�!�s�f2�"Ou@W%� f�^�B���*2}�e"OL���I�CFլ8x
�W(��B䉡��ە�I�t0��80B<��B�	�;���1��Dt�����X�T��ds��YK��t���MșO����M3D�̑��ҟp��K�ǀ	c<%H�=D� !d���I'^�;Tņ2>q�Cc/D� ��`W:)^��:&��i���)��:D�칇�lk�ǫ̻`�����:D���v��Izڭa]�N��;�8D�<
��Y<{��Q�����P#�f4D��³�ӗ_�,�"�M؅euTHG %�?�Sܧ�D%��P��C���	o�d͇�.��]����,D2�2#c�U�ȓFt�3�K��ڟL1��ȓ��[���6�,:T�D�� ���I{�'�윫�X��0�
U�p�~Ի
�'S���М&�P%�D�^8c����	�'	HH���k@�@�d��j�~M#�'l�8�d�Q�0|���+j��R�"O\(��aF-��I�蔵.��pz�"O��Qˆ"h�4��3�\�`��y"O8ՠvdϓ,݀��1N�/}c
��g�'k�OR�?]�OG�Zamͺ"��*����}Dz1x�"O45��(c�z��@�4��aZ�"O��f��/����t*\d��dE�'�ў"~2Ï�G�"����.S���&-�:�y�h�a�����Ըi4H)��L�yr�H
��{�9 �Q�J��y��_0GG���bI5t�NY�p `���Pov|Q��<\��R�δ��ȓR�$�c�-{��qг̀4{�\���ff�<�֢��pB&$�T�.Fj���Il~Bm�1K`�B�	�zbXt���y2
ʍ(tpR���l��@��EX%�y���B����G�,g���S��Ҡ�y҅R/���r&�^ڑ�
�yOO�AǪ��p��� ��a ��O��y2��
�b��N�e{�����y��QE�m�61J=�p����>y�O�y��C`Q�po�8d�.T�6"Od���LYVJ%p7� �^6�0 "OȤ%H�FmZ��ݙw#&�t"O&q�D�)t�y3.̔T���"O�����A���B_����g"O��'aބin4 ��Y�D�8�"OL$a ��X�r��$gu>ts��A�������� ��zy��#�O^˓��S��{b·,ԅ[�r��t�3�R�:-�i���� ��9�˚j��%K�J�6^L�!�"Ol�� ]7T�L�yU%�J6E�B"O�u���ؐa(9�#"i���"O( �Ù�K"$��ļs���y�j�U�1R*U��%�aa���y тbج$��U�\ő��?y	�'��� �I9=񸨰T�O�}xx
�'nА�,�V-���cA�*� eC�'�Pm���\K�mX�
͛$��L�J>���IL�~kh�ZG&�/^��89uJ �B�!��(&�MASm�q��mi�C)��r8O���F*R�@�ζ)�Ԡ�"Ob��]�"��b�G��
P�5"OJ����U�t�����cC4o�P	�q"O�h�mXl_��Ka�UW�0�"O��r�$΍nS�pɴ���W<ֈq4"O�(���_����j]/ۨeS"Ov�2Ǆďf��q�cȇ!r I�$"Oɲq��t>:M1G��#U�d ��|��)�ӟ���r%���vQ@Pǖ�s����(x-Z�r�e�_����&�?/��Ą�t�ۡ�Zk���K�9{e�0������rGڜqQ�]��� �ȓyR�)��@��)Y���D�˔���Nd��I�
/	J��4��{�6L����<�'�&jP2	2�"�[D���n�<��c��;h�Trrn��xhZx�A�r�<yp�Vu�x�Pa�Bh3
�i�O�v�<I��,<Ǭ�h��	D��	L_s�<q�,ԧy�(�BFh�c���Q�q�<��TX'J�k�Cކn��[��D�<�6%�`�&�Y��Q
M]�4�R��D�<Y��ˠ:�TŊbP�����g�<A �3�P��ed�+b���8T������9�0ف�e@-1�(��a.D�d�'$\(c�Y �gK�A�b�2�o.D�8�cȓ=!�ReK09�g� D��QQH����K&��5W-����O=D� �̔�>l��N��*2q��5��0|b�JX�8�{ca�?Q�6��Ah��hO`�G3��4B�r���FgED1 �B�'5���C
�R�4�񵪓�1薰��'j�k��^.��e%�0��1�'���q�
I�1,hcԂ�.U� 	�'6��ՅO>W
t��nՃ.�Uh�'�8@0��@���A���g�&�	���hO?� ÕO��߉jRLP'�Gh<�AmεG��Q�=�Na�ק�	�y��CCl��4-de�&�I�y҅V3b^��V�������bEU��yb@[�����	)�K'���hO���I�mI�,pt���(a%�\Y�!��E72�<�����n�s��ƎWHўt�'c�����K"a�(���%�A\̠���O>B���c�c���,~H !���]~ B�ɾN����o�3��j��@���C�I�/�>�8a$L�@�ĸz����(��C䉢z����!X�&l��X`.Y	4�C�I�C� ���C�@��x���C�,a�D���O�)����t�mrX��d;�	:8V���M1on��B��0e�C�I�?<.̓��|�l��OV�}B�I(T܌y��V�\Xh�D�C�ɞU��1R&B�-L���+�͘B�)� ���i��,fHI�d�z;N�J�"O�܀��<u�@���$:�l@f"O�����	O��˷�щC&9����F�Os��8q%)MI0@���(���'\�CMP�H���ʃ-(>�lܱ)O�=E�tcT&8�X۶�X�5����^��yҥP�y�&��p���+��p�#'���y"㊐`T���kK�!K�!�r��yb��F&�ݚ�bĩ}�!�r-ޯ�yb$_FPР�`#]�H��eyg����y�@*N�R�匮?Y�)7$ɔ�y�Eݔ�S� ��0����
��y��0Sl(6H#<4�i��ɉ�yrDB�J�D]�(ލmXʴ�uE�ybDF0X�~HEќL��I���y�	X. ֘Y��	}D��DM�.�ybK��p*��G#0�� D��*�y�藵U��(saCVjK
`0c��;�y�DN�İ�2�EA�_$0ezwM���y"�ݏH>4Y�%�.]�T`	�&��y.��:����A�R�Iys�@8�yb�߁Uf��i�!��6��3�Ө�y�h^.&̀�q��z�T(D���y�DͷxLZ�r^�L�,�Ƀ�Y��ybM��Y~� e޷o2|18�/˩�y"�ް]�d%8�o�[p�0c�[��yr��	}h���AkGԿkH���v�I�AnВ"}�`i0�9KCp��ȓFI �)�KNfH��a۵A��t�ȓ
���g��N�z����A�]��j���3 !V�$Ȅ��C�u.��ȓ�d1ҕD�Z��0�"��H�Ԇȓ0�@����^�$��F�Vӈ�ȓx�@A�dϟ�\L��`f E<K.��m4$t*��>Ϯ0!��F����C�t�����e�����gϦ�ȓH�ȩH��%n6j4�p�YN�Ȇ�� +�=]�*�2@�w9r�ȓ>
�x.U��B�ܢU��X*R�;D�8��	���lx�N��Y.hY[ �8D�$z�/.^��L�įF�;-,!QD9D��b��UY*"���X��E�Ё7D���h[�^��IAȄ�8=~U)�*6D����9��x�.E�(Sh݋Q�3D��ӵ��$p��X"v.�3{X�07D�,b&'T0N��Zs�	�g�H���5D��G
����v�[2\��)3D���2o�����^�.���"Uj6D��K��X�co�P2&�;J5z��!�.D�(��F�4��	���|�z1㑎8D�X�a��O �б%�	e���ۆ�+D�\9���:<S���@ ^����)D�P�) ^���'��6t�Eғ�"D��b׉
��`m���=kF���d�2D�9RDQ�A� ���W?]�d���.D� S��5r稡���%�Ri�-D�䛁g	Ju�5`��s6N���H+D��w��>2�Q�b�Q�xa�F�&D�l!󨛴V2@����R�b1��)D���&ԩi�Bl�[$C6u���#D�tض��#S��ѻqɛ�I�X�xSb-D�@�b�z�\@�_7G%Z�-D���D�\�SR�<"��
Z��@5!D�lqaF"̠aȷ� �L��7j=D�� �!��D�D��Nr���"O�qaF.�:9�u�U��#q��"O}�a$&e��h9s ,��'"O����!D�&ٚɚe�W8o��""O`����}wN��P���#�|� "Op��s�Y��2PB N�G�hh�"ON=;�@�N�� k�A�8�`���"O.aQ���2��w�b�	c"O�Rŀ�>N�N��u�Z
O�V�"O � ���,����0n2��%�"OFyqr�V�j"Ǆ�"5��J "O6\�v(Ͷlbj� �_v����"O¥c������u��`b�1�d"O�3&�#�f�R�+A.{u^��0"O�h˔eܿY���0���e��x�3"O@���G���
�7g�:E�ȴc"OR��4�֕w�h4z���lup��"OT}��'�s$4�X�AR�`f��c�"OF(pB�=9��\:�!��(l0��"O,y`b�+S��U3�+�%{\�)�"O��:�,��
?i񏍪XAn��"O6}��n�j��d�%D��^�<�b"O��GiΧ`����i��f��	�A"O�+��r��(�3s԰�"O*Q	�"ٽ%J`y0g�)�Qqg"O@�(@'�uU�@� � �h9�"O���#�ȥc/ �
3Ɋ�7�q��"O��1���M��r�ؚ����"OX� �f�\�
P�AݍP�d�8�"O�i"W��7)��a3A�~'4}��"O�{'`�U@F4� Òe:p���"O�i˳�@,v~Ա�pΎl:R��$"On�8��[����T�='�0�t"Oܴ@��K<\͎���{��t�G"O�	0�I�y��p�J	g�>l�e"O�l��h�F��ѧh�1[���B�"OD�0&�MbZ��k凃'M��!I@"O�ಠL�"I\���"7��I�"O<����	4VĖh�$�	��F�Y�"O"dy��̞0�L0�f'Q����"OJ�:ED�>l���2W��g��8aG"O�] 3�
BS����)X*UB��U"Oz(����ތP	L	\F"��v"OR�*�V$
���	{�|y؃"O>aq��J�E�	 g��h���K"O�uZd�_�Q���5��C��ݲ�"O�� �OA�X#ʰ�R�"���p"O��a7-�7!�dB�"Q�`!!"O0����&V� �ʐ��F1�"OZ P��O�T��J�T�;�"O��2���o6�s .&��p"O0��C�?�B����ό&���"OZ���l�. ����C�H�Du#�"O��B���%vd�@��6u�&Yh�"O�)�w��<������/y����"O��)l�(hD4�����.���R"O�3��/J��R �
��Т"O��Д��� q�dQ4a۠(�La�"O4p����m����3uJq��"O|mi���?R�a��ߏM�q�v"O
�@ɐ+c�̄�V㙺e-
5�u"O�]�/O5j����#U��xB"O�4�v+L�#g���G�H�%�S"O.�u&&�c�mQ�c<�y�""O� :��c�a,�-�6���"Oļ�$���CBl9�0���F� D R"Of!ZA��L�R����3~^���"O�Q�?e����IO&G�|�#q"O�����ֹ"|@`{6B ^V�� "O"Q�pN݇6d%�U�fr��`"O�L�t,�d^�U�6͏	xq5`"O��Af�	�e���5-���zq:�"OT��VA�NI���j�H��@"OV����&�(�B�kE�[��q�"O
h��)H���(��5]r<1E*Ov���;XC����"($��'J��B�R�n׺�����0��ؒ�'Լh�`�S�gg�$!�΁_BQ��'�Rջ��
P���A��@�&�\P �'?��J��Ͷ�ԙ���:�<��')��J�����2�Z�	ڼ��'�6)8�'�HD|�`*Y�����'m�hiei�ĭ�IΞSO�	#�'�X,��*U/ �6 �G�(X���'[��!��]�+!�1�G��{��d!
�'���Jr��|����r(H���' dy��Z�dA(�C͟W�J$h	�'���5��."r�Xa� �y�� ��'}x|r.�88=�%� ��-yn��'�h)�oԌT�j� �/�
n��a��'��t��ȃ�ՙ��(U^�
�')�sJ� c ��2F��8�
�'���CU0g���Yrǋ�Wnn���'�:  a��<���	��W����'堸S`��c�J�p�M�e�P���'}ޡ;W�א'	( �B]�_k�i(	�'�A�r�ǩ0�='�ٝQ5�H��'5��n�H)�@+F�D>ȤY�'
�`��.p�y�5B�;�Z�!�'?���j;��$⍧�%�T�<������Iޒb�z��6CXv�<�1�[�.WBxJ�!@�yH:|�FXp�<	f��(���C(]b~8hУ
j�<iA�W����3T�F���\��g�<ᤥ\!EFh��Μ���h�傚e�<q`,�
A�(���ė�&��|'mA_�<a��ԣ3�^�@�.�n�0��@\�<���ӪC!�9p�% �LZ$�[�<�%�G=y��|��
9厸1��!�ƣI��Q�!� dz��8�`,hX!�̔�b�s�gT2���j�ʂ�QX!�DI��MX�L�G�*�Jv�]j!�d�\������ P�⩢ՍI�s.!���BE���E(���F��6mΕ^!!�F|�h4ж�D*}�l�:�I�!�$�7�<C-Ɔ9����ǐ�=�!�D-@KZ�F� ��C�J� ��j�'8���e##s.���F퇔�x��'��j�AF���HA*� }&����'�.%)B������.6hӄX��'�Li��
�U$�!�h]_rTċ�'-�%� )���q���Q���J
�'�8�Y�C��V^m�Ԏ�1�d<�
�'bt�+�@�P�)7d�$�v�+
�'7, ���m#�mJ��S�:М�
�'��a�#�@ @��;(� Z�[
�'�i�"E��&��c��g<��	�'����c+J�[l�(�f�M��
��� ��[ԋ����˖��2��Kf"OR��S*  �n���Cͩi�Di`"OV��L�3+�4l�'�8*��퉃"O��S��_�L p5�Q��-̲�k�"O|<4��8�maUX$̀MX�"O<]WIոe�0 *�f��A��Y8�Щ�OI�	�����@]+j�4`.D��i����2>xX#*%�V(�Ch�O� ��0&B,�=�<��o� wԄ�xa�d�OF����f���)U*��dx�@"O����:'#�TZ���	 `a[T"O��0e.ˏty�-�ĉ��?�T1�"O���u]�n�L�:%
�9�܅3�S����:�S�OZ�5��#��%��	�� �j�.�P	�'����D��$�J  /��2vX���'Z���Q ћH��!㦍�{du��Rn7�>3������ -Ī��Ո��r;!���)8l!��咉�����&�5j�Q��D����35����< n��e?�y�"�!}��GL79������yrhT�=���PukK��|�y�#��y�ï�i���y��p�g�X��y�O׆IQ��4g��}���!��O�#z�$��F|���q�8򑍈z�<�E%q�%9C]qUlْ�mE1�Q�E{*���V�	�14���J�:\wԘQ#"OZ�i��.4� ����2���@����"d�,{��u���Y� �thrB���>��O �0���3 ��P�Q,����Ǵi���$�1}��xAԦ�\��Y �Y�\O!�$[.���!�Н�l�a�<!򄑴>�ya6bˣ��ڀ��)2�)�'F���8�6xj7��e�L|;	�'F�X��#Kny�����XjF�`�'��$�N1]�J�y��a��ɱ�'��p���;�:3�b�p����'ў"~dfB<w��d��M�\
\{�d�[�<��+L�f����O�'.�F\�Ȱ=9E�
�ڔ�+K�q~H!A`��8�<��4G�~�����$�M*�dڦt�"]��]s�ѷ�".���۟L�6a�ȓ\��8��@*s�0� �Ť\�lH�ȓ�l%P����b\��Ś���<l�q����0l����k���LmH�N�F�C�ɵ/���ϓk4a�)�-U��C�ɵi��q!W��PP��?]�nC�	��Np�`+Ù%㞈�+6�:C��>ag��c&�U7F+>8A ��Qz�ʓ�0?�2Ε!Y�ҝys	_�<��Tjx��3*O@X	�حBHR Q�^�����"O�Lr�/L�h���A�>�Zex��ɒ2Q��)��^<a���7W��HG8Y�Vфȓ=f�lq�A`��}� �W��F���HO(�}Bp���
�kg�[# ��yc��K�<1c�W83d	Cc�6]~�	1�N�<B�-xӚE�0o�D8 �J0@N�<q ��o��A_4L% !2���A��F{��t`@�ȐMϬn�R��FHN*�y��-g�N�� ��B�FgP��yIÜ
J��@c� #Ԙ![�H���'Mў��(��k� �8��R�k���۶��6lO��)���,En�éB*���W�Ib8�+���x�\< n1/�e�&h���S���	��H	U�S:2�09�-z�z��DC1򘧀 F�; ���Yеe(�ye&��d"Op �d���Moz=��1wI�9���'8ў`���p�$p��F��B���it*.D�ti�ϝH����3�H I��R�.1D�t�B� c0��bG�\N@���.D�x�2 L�Y�X �����WX��rO"�O�扁 �j�Ђ�:(ȑ�]�d1B�IjN�y�i
���9��@�� �"?q��ɑ�#x���ƛ3hK�a�Rkݑ �!�䒇K���:R�W�lI�5�����������]y��I� <�q�,E���*c�ޱUJ!��ҧ?U6:�� �ڄ�N�@D�'�|�t�m�C���Dъ\IC�˫�yR�P5`Bg��5^E�U��O>��Z1,��0ceFI"O���sO�ߑ���?�O�
��EF�nz�k���:w��\a1O�|	F=Q���IŘ�����<G�Ԍ�~�d���
:P8Y��F5�yB�[/N�;�O0\$����yR�ֿ6�F�d��^�QE�٠�y�
�%;��!�4A^��@��J��OV���
9�p��kѳ&JL]���Û3!�d_�e��HS�@�7��ꕎQ2&$C�ɴe�d3�J-k�.5Hd�ϞB��B�I"@մl��I���m���4O�b� ��	5?�����U�(��P��Jh�O��=�~�'�ӻ�vL
槞&xR���o؞��=ir/�u�A�a��2�L��Vj���=�f��$q���+"O|�fg�<��
�#�t��i��|	�r	�c�<��K߂M*� �r#_^:PB�-Z�~���~ښ'e�p|Ƭ��m��P�j�0L�Q�\���۰?�����|����$bך ��m�O|��w�$�	�?O��D�&/ƴ#��Ҁ�H)�:O0���K�h���Q�(K����`�L�I�!���p���Y�]�z&C+�!��ƽmʂE�!N�c!��kR ِ|֝	��d,�S��/�1z���Cō2g�֑q!a���O"�Ɛg�)yq�3L6.Xȓ����G{���'��`0C�,��xAF��O�n�m�������)��M��О^�
��4�	$C ��`Q(�O��0�^��mD�Y7ZY �%X+h���6f^(�,�8X��I`7��Af�d��#t ��`�[-�;���$�����v9�v��0�P�C#ڜ� �ȓE���Ūz��c�͛I��D��'p�a[�H�Tz@1��Ѡ=p4��,,0�
�`�\��w ��66�H{�'�T�0�U7�< ѳe08@<I
�'W�P�בd9^I�'�B.0�%�	�'	���f�T ]I��j��3/�x�9�'m,�,��4�b�K� ͻ+İ��
�'�$92�[V�~�q���)"�$ �'�rsvbkW��Z𨊦�$��'��@�w��_��ᇌǋ�>]��'[�%��^UE& ���I]H��'�B����=)ن�1�7J��l��'Ʈ�u!�B<��WJ�V��Y�
�'��`�3���)�M����'~��C�6�2����\0=ε��'��@4��i^��J�FߡJ_8q�'O�Xk��)z��sf�2>�����'��X ��:T�kФ:0ļ��	�'���H�Lٍ�∢'�>�0*��� \�Y�D�]�z��� �_{��X�"Od`:G��/ZX4Q���:|�A�*O�(:�ˋ�~x�G�	l�q�'=�3�i�G�
�2a�;ňA��'�&��#j�x?
�8��M=}���'~
���)�:��A�WE�y���)�'V�j���S}�����O�kB�
�'GHqt�ٺJ�va`���[���	�'�*=Cs�ߣt���ǈ�2\>���'�R]D镩C�>-�&�	5�͒�'LN��D 3,j�GP�,�V�"�'%�;��ɺd�F}�eM��5(��'@� RO�M�>��E-!+hzl�
�'骡�ՍųW�����͑)8VhP�'[��2���QRh\�t�&9#=c�'0��
���>#���)���g�� �'J.���c� "Q���v�/S�����'���N��<8F%Z��f��'�j�#RÛu��٦�ıcK�I��'^`̩"��*?�*�A��݆YWr0�
�'��O�P}�z��ˁSv��x�'dp5��͏#mtJ�Y�N�!P�^�B�'l��2��J��)��RS-
�	�'�ȔP��W55�n]J4��'D��p��$���֪��Jc@�z�'v��;��"R~|!��A�.i"�'̚<�"e�Ui��B��I�'����_�gy~�bÅ��^Q�',�����Ƞ��"��"�8Y�	�'ȊHj�D�v�1`��]�
���
�'8]����8TFJ% vc�<$�	�'���*�!�Ey�Q� �lU�	�'���I"Vz+��B��5��#�'��	h�ϣ'/XZu�]'�D��'�"0L��/Z�"T c���'VHAJ�F��"�4�{���.0�
!��'E�������J��X�m�+/W�H
�'�d-AA##&�\���N�"1
�'��1!�%[8I�(�(��^;E�ȉ�	�'���ip≚��*�`ܸy��'��9x"H˚��}�c�	�Y]�ur�'��M�@�%����Ȼ\�%��'��!�"X�7<&A��ӜW�-1�'������~K ���VE�.e��'���s�Y¤<�!�D8S����':h�t!��">b�Ҁ �3=%>���'��K5ŝaN(1�,a��i0�'�ּ���V�n�n5
m�,
0N<
�'������Z�4X:F�ґHO���'��(��nX�DNb�yA��L����'�\�0sA��P���e !Bo�pX�'��|�g���]0d���A��o�ʁ8�'��pQ�K���>�d�*Ƨ�)�y�`\������0�J���!N��y��z �Q��A�"��\Q�A��y��>	���	ǌ�+J�"�Q���y���)�VQ�Á�>Y�LUR3�y�dۋSa
`�W1�x�����yR*7qJ (�0�4v��$�%�y�oR0b<%z��3�J�Z& ��y�/؁(E`��&-�(4G���J��yB�Z�t��á��4���2N��y��B�8��q�@�8�60[r�7�y"�J8�ؐȳ.D-0�|�{�߃�y
� ��{7a�h)v�?8}��r"OL�i��_$T����eY�zo�p"�"O�ej↛�_<|e�����Wo����"O��玱j������0zk>|�C"O�j1*	<u���fJRG}�1"Od`�EE�^�t�5�'6����"O��2w��]�T�ڦ�� T����&"O�ī`�3-�I ��o�H���"O�\���J
^�X�樜#Q�t�a"O��C K�vӨH*%��G"Ox3��.����� �a�����"O�,�� � J����³!�8��"O �`��)w��yaCq�z`�"O�1tK�<|�ex�"��z!�$L ���roJ���*AJ�S!�O�;�qPd�	�%3���Ys�!�D�����O&�e��`éI!��*~`�� "��G��`�'��Q�!��	�J��A(�3���WcL�^�!�d�) )��Ӱ��p�0��� �)+!�U]2�}�FdQ>��x����H!�$�ir���,�;`0�pk�'_�N�!�/w��l���+E"�83Q�×C�!�ǻEd�9� ��������$!�d+0��o�.D �Id�9>'!��	�eB�!A�U�q�64�'ʵw6!�d�:mpb��_�<�>�+u@�P'!��T!z����M�8������)m)!�Wq&*�`c-	o�	
� P#3�!�G-?����폅E>��Ů�	
�!�Nw���b�_'�J��S��Q�����v�?��(��B�f���c�MZ�&D���'J"~"jQ�6��*?�yQ.|V�0�g�Vu�)��<QA��s�^Գ�'�9u�&����](<)!�B7[����a�"`�mQ�O�-E��\`�Zy80:6aY��=	 ��.6'4��4�6R5��C�(�G��)�I�&C����ф� @�0�޴x7 ���̆z!��Z�D�4��)�ȓ�~�ac�R�b�#�-��v��8�'EN9�%o�k�!r" ��Zl�F��&I`ܙ��oVt�	SĊ�<���pA�]؟P�!Q,�Z�B�n	?�N���Z}
	�"ME)e������#]���l/H5SǄ���c�R
#k��$dN�IV*�/���S*��*���/)�����7G�`�B
�1|���򂀎O�"\sA�'(��K�@��B�_��8o2��d�;Z�fQZCB��D��?٤�ȑO�p���)��Jp�{�iZ'-�Iw��@��Ԛy��Fh��v�F�'� 8���Qb�g�I-)��bJ1m���ڤ�]�X˓(��Y����{ul���JD�~�?A1���	@�u�u/�(\a�-�5�V�n�����[�a~��ƤW�4��%��4i��RSF��@�vp��ÚZC���MV`���a؟0����X�3g���O(j`�F)��d��h]L<���',	Z?��ӆ�7t�<�cѱER$�#��:kt^dC�Π84s��>���"�SMń<�BҚF�88[�!9�J������ ¦�X�C2ёu:O���p��-O����Z�E,,��r	��
U�9�Tx8#�3�3��BN�D�� I�5����ǥ5V�ɶj2Zac5F�Hl�@��	64T(��D�H8 ��	aWL�}�,�ʁ@�5��;��w�a~H��cx������%<����ӱ���g��X�( >s�2k�0a}��Ҡm�$>���ӼKQ�ťE��]����Lk7��N���s�CE����gMN�l3XH�l�T}�p*�����@�v#Ձg��9Y�GLg?�v���  �Ӵ@��}��j�"�J����,6J@D}b��;�*4�K�I��	�rS?]��l���}#W�G�TZ�Pe�<��M\��vpY�",O�)P���8v�BT�d��J�ƴ*`1O�{W��J>8 ���* �!X��TΌ�� ���8L�5 "/�3rbt�����Z|�ē����ǀ�v?T���,S��^r�x�Åc*Ԛ��@-��ѩчA	u>��yG�ʔ$�z݂DJ� �r��nP���>����hR�A����Vk^�lo������q�X��뜽d������?}2�8~�`�ۃ��4a�� ՚������~�J�`� ;sў�Ab�ȴ"�6��&&^�0� 脮��|� �!�惒�e?F�������J�\��8�/�;��F�'�l:�D�:{����V-�#t'�ɀ�N���G�Xmؾ"�b��[�d2I~JW��[�b �4o�0��)^4��-[V�ӪZ�B�I68�*8�rG�

���גjH�O.t4������d�A 69� ,�2'J�i��;$�A���p$�������*�O���U��Fi�L�/��6TM� �J�
�AÔ��W�j$0��	�O�pyd%��')B;싻Bێ	1��@�d,��ú�;��8}2EE	a!�Y!���2'� 8��l�$bS�Δ�4x� ʿ*&R�G���7�!� �
H9sp#[��0٣j�&	���T33d���K�8��M�@.����A�if��D/���G��.���Ѐ�uSR�\����ܵJ�Dl�-��*@(Oʸfn ��N�G��\˖O�0���k�f��N檁2$IM7���	�v�0��Ā'�B��3��ׂ�<q1��s�$����/?���Z�~�AR�L�A�Y�bLZ�zqz(�q�dl([(����K�d܊��p�@�)��I�.]�#C��c����Xb��>�[�V����E�9mީ����-sH*2f��8�̍|�p�1$$D���	��۸��S͗�N��죟���T�n�|�7,�aJ��Io�D��&�&{��S�*6h�S�	�3*.dm؆�ٽJ����$[d�2AJsJ��|(�u�	�X�:y��	�
ـ����X��䓶H����H���3�	�Bی V�DQB1�$�@�Z@Ң<�E��Gј9G=�'��)�傳:�t=
��Z���D$$^$4��m7�ON�qC��.+ ��'��8�!"�T6�����@�}�1kF�ᄂ� �槿ta�J��h[B�
����F�<�r.G~�Y�e�9��([�}?�#GM�+�f�i�9}��N�w[����H+��j4-�����=�
��d����>�4$�r�46MZ�C�(�0�S�EL<��5�
0J���X�3+�c6���Ջ�ޜa��T+O ���GKfG�~BÙ�U(,T�F^�q�R�R�����b��6d�Q
�iU.d�a}2n�n_\`�gU�q��i���O\x۲��=1���{��*bBZ��&H���ʑ��!��u���W�]H�C䉕y��*B�%�E	��|���x�X�P��-HE�4��t�?=�c�9xG�!85�K,V�8��"%D��c���bs^H��(H8�VP��?3@�v��4N��l�3�Ŕc�����'Bց���T�h
� 1ynP����4)	��Ξ2w(�##��]�f�;���*���y�gB<4.0A�(6�ONI��2D��E�,�5~�d�+����u���p�b�R}�t�٤m��p�q>�0$Ș���E�Tx�� �#D���E�մd���3�`�	\�be1D�	YaRYcFlX:%��U�֔N8���5���yWo'����+A=m.)��j�9�yR!��%�tm�<���E���S���2Iиi�cڌ*\L�bQ�9 �9�����Nf�$+���*"q��A&jݧ�z�
�"o��
W)nq,���X�ƽhլD"mm|����I�А�����U�N ��I�]}���)K��8��E8R�P�La�b�Z��ܺ���w@E�6G-ʙ��Oin��EV��Fi�#h��,[�'%����UsP�p#�nϓadJ����^�Dm	W�L�0��,	f���H'��?��39�$[b
ϥ"�
��l�P�n੷"OT���ME1�1�
�&J��Z�GE?s��$1�#�t�
e����tyax�H�mE��@��5I�&�cW�ݩ�p=�0���̽*�j	#�M� $��n^�S�ʤTn DK3,@@�<i��Ă'f��{�`9���Xܓo��A�p���V 49�􉊖:�,`iT�؇xoR(ڱ+ŖHP!�$\�䮽��A�^��ͲqL�J�ʁqN�:[|�'��#}�'BH�'O�f
&���]"Re�
�'���`èȧR٤P)⊉�W��Y��6��t:���0>y5aC�'^�[�JX�}.l� �`
@�<1�F>\�>�yB�I	2�Z��gK
x�<�K}i:�k@"�p>�� �x�<q�3�f�G˛<-9F`bMy�<a4��!v��.ټ�y����z�<фb��]�.|҉?�&�h��Y�<�B�Dk�AB
�fd0��%DQ�<9�h��-[3�Rq
Dc��L�<�e�ا
� ��b[�H(Cm�O�<���$6��Sf>$�0�J	G�<!�+\$ܰ�Y�&�'(�^�CgM}�<� �	 �C�$<��<r���R���!�"O�pA䠛�g�}���ڜD��بv"O�dbI��8�V�@7���v���y�"O �X7 ]�~��F�B�M��t�"O����6zr:�J%'�l��`�"O����B3_P8iCF�.tH�"O��e6Uҩ�Dd_�o$n��W"O�):�.B�o�-@�B0�4{�"OD�'dT�+@�I�&���"O�p@4$ӗ"�z��e�^5g�>�"O����fH V�q��@�^�6\�"O�i�!�ԓ=>)��'�I��8"O2�����bp�l3�i�3�J�"O�TC��A/z� ����
���"O���WbV6�&Ȓ@��O��!s�"O����-�'_��97 ++�i �"OFU i	
�^ɸ�j�rg�|0"O`ͫծ��K��銓��T�#"O�hp��G�^��J�.J����"O
	����xԄ|;%�E{i��{�"Oz��԰F��h���4^|�s�"Oڱ	�,I�t�c��=D�x��"O���-?�J��O�0~d��rw"O��;t�U�Oɰ��H.Ch�"O��ҥÏ1eH��"--J$��K"O�̫���h4иv�H�N)<e�"O�PDʕd@5LƢ0+25pr"OTp#�B��b24�b�NR'��G"O&I�f��
;����
;+Aj�"O� [cB��{���%��P!<��"O
��MǸ'�^�*�`��s�"O��A$hL%�<h��>%2��9"OFMxv�O+��u�c]&�Hy�"O&ɺ�m�4zǨ�sp��u�:i��"O�Ո�K�%�t`ۆa�4R@��:r"O��ȳF��֮�) AVAh"O�DP���	!��I����K�V�("O�:�f�)I���� �
5 $P"O,�����ū�צ3
D�hB"O,��T���;W� �瓤}�0L�R"O��b�EI)�p����j�>���"O�HA���D�� ĨU#X µ"O�1A��B �*�Ͻ7-��4"O|�0U���8�M+Q�K6>��9B�"O�4*�A ,%���A�1�h���"OJ�B�cN!?�I8�L�{�<kw"O���nȪ4#�q�G%Ѻzer0�F"Oh���B+6�ƌ�҄��,k~t"O�mq�&5O�T(2�B�'vID@"�"OX��a��?Hkʐ�wH>&Ya"O*5��l�I�TA��9^�D"O&��s�ǾKV�ҧ��'6�\��T"O2Q��^&h-� �*(׼u�"O̜�qDR)c��X��Vm��qD"O"��U%�8aDblzGj��0�rP��"O������'_/\(�1�����q"O hä��w���GaՓ{�|	:"OR��WIE(E��a��E�&ƈ��"O��b�`%\ڌ�1�X�-貅�A"O4�D��\)��q!�7μ��F*O�+$�KR_$�P c+]:�T�	�'��Pj�Az�L��Q:����'�⍢�'�e�J�&oT�x�h��'����bM�:b� ��[�z������� <ܨ��R�7�y`堞0�h�5"O�It�=qJ@ԎڇF��,h`"O�� ���z���- ���A"O��!�ـ�,h��O�8t�'"O��+)w�T���Z�^4<�@�"Oj���C�z�=��I�(.�r"O\  Ҍ�7��`����/��"O�-�s���~�{"�@�r�4�P�"O~�z����N�2�W�q�$�;�"O��lq汈�/���� �3"O���H�lڤ3���f��!*A"OL)�t �(h�)�A�X�Н��"O���#�ˆ/�Z� ��5$9y2"O�i���i�%��C����y��"O�!r%�k2�u��cL�{@��"O.)�@���p)+gE,D��"O�hsr��o�xkq�_2@ rQ"Opx�J�H�VyJ�-��bpPl#�"O�e�7	�0�!E��]HH#�"O0��c@��8�J�#v^�3"O�]���8	�Y���M�jK���a"O��"��$�:snۇ)R޸j�"Ov��n��|��g�F�H*24��"O2�Y�c�%V��1HR�(1�4� v"ON�*�b^8#\h�Θ�I��t"O,�ѲKC]�Yz �L6<�lc "O(i�f��	t�����.�']6���D"O���@��>(�#lX�+p�	3"O����QWȜs�+йQڸ�"OL�ڒ(ڪ;�c�L�#_����&"OKV�DF�E�g!�+LQ�S�I+�y�ˇevID�Fl$��^��y���'� ���n�
?I�����F6�y����~Wtc���5�ޙҁ�C�y2�دw�T�Ab���*��a��^�(O���X/���*@�c� 8S�U1�ĝ�B�ܬC�"OP8��㘜 ��9ҒޤZ����,i9��)�J=��s�x0e��qф��2"
i L� :�8���CC~\���^�Cnr)���Џb�\9*$���l����f�B؞���1l ,�VOK�h�R 
D7O��@S���xX�]�4B�"���oZ�2���;D/W�8�.A�#�/XhC�	*p�r$�Q��<����@+R�FKT��d#�H�`QD�]�9��|��"�v�|`���9+(� ���?(fd�A�*�O`�1G�9"����D��[۸e[3��8OnT�S��K� ��ڴ1e��I��p"G�o�Ā4N� ���=�E�M�z]��e@5K�œH�s� �ؒ�N�~�h��Q?l��`ag��)+���GL�:�Q\��O|BEy��H8wE�&W�@#	�J�'�i����t��B&x-��;�:1K� $4�s��,��ݓ0(�s��ZV=��L>�f͙Y���B�N4Vv�����vy��ʰ>�@�i��-TװEC6�x�'j�"��Gꙿ�$�t��lDcdA�e��Fφ4�0?�$�%��q���8y����=M,�q �
��MgϒFH� ��O'��!sEC;~��8�'{0	1��ٶ]I� p��&I�E���ky:	V�#t���P dR%2e� ��%֬X�p z���J,U
��_WlٚM�P�d�ܑ
�@ ҒF�fV�]HwA
�D�axB�6�. �B�øZ�4�'Z�Ay�%��'�8T��̿|�X�%����	�}'�l����|%;J��DxG�Z3
�H��	����I�g,H�KӯZ��0sW�)�yS���4'��PĒ�	�
*�Ӣ�u��ѫŬ�0?�d)�7w�����9N��ȥ���J�xiS��9�� =H�zi[�Y�/������9%�q�!˧)�v����9D�܈6
�T�1L����VF���=�R�1*�U���t"V�- �>�K���r	
�P���'�҈abX�<	��V�'NHQs3M�1�H5�)cybMM56Ҍc���dX�x��k�>F�%�������"�O���B��4{�����WQ�l;�H�9a�<�&\���x
� h�3���l>ɚ��M�WC�Zr�I��X��g��M����@Z���%��$1��C�ɉw"O`|u�	Wr`h�ѷ3�vP��'�� �' �S&u�O?]��o�B
q�cK��IT����y�<����*B!�!E�̼��ȕwy���8<tDp�"�cX��YE�E�;-�h�� ;�: c�-$�O8K���V2P��F�aB�G�,eA�"f�ސxR̖oBpE�ӡI�M�;4�\��Oh����H�
p8�?Y���gc����$��Pm���*D���ǡ �[Z�y�I�Z=Hf+��@���M36MqO�>=�qi�x��a�FѲD�9���OIx����������x��[�Pe���6(H�,�pa)D��%e�4G�2T�F�e���4��>��!�7g�%��ep���G��TQ�m9��D��Ą��.X^�b�Y�l1��tK�=���C
R�^JN��F"Or�/�b��j�) ) f+��ɱ �b,R/��`�O�v��ŏQ�d0Õ��;Qs8bF��Z���z�l�򃞄D���g#�2L6���'�.3�ytkY@�DO�,StĻ�H�s����ICN�g�N�@���3&�Pe�"O�1I*@�����H��]�'�Opz�H�5:<�XL�� ��Q�hstܡ��\0�ͩsVD,�����P����n&�OFuk�Z��P�l�%u�Z�9��s�	Y�G��I�%��%B�Ԏ�axbL�>ӊhI%��-C�JL��.�(O$���E͊;ۆxYM<�u��qL}a�P�
5K��.tF�����T�!�$Ǯmڵ����
?&5`d�۝}Or�ʖ`��:������>��m��p}���'}��8���S��|޼\PG��,d pM�ȓUOvD�T�U�)W�9@���3f!��{��u��<��'�\ͻ"��&.�O��LHq�R?㈜j��;@��	�D�ˁ*n����ƣ����`��T�U�>	���%Sˬ��v�6O(��S4P���QR.��D�Kg�'�֍� ���݀���DŶf�ڱ�F�ٳJ5|(��MțiKPd{��'��y�#S�iP�a��!S5�:��$N#���h�*��O;���/�?A3%/��j��;6�C��<��;D�@���E�<���_�y[�؉a��>�ǡ�M�������h�,lHb���H<B��ݿA��*/K���$�W����(	xǤ�Qd^��)���M���'�JB��q�~�?���O�E�����@��P`x�a��4��;Ӗ�:l�=Y^�	0�Kԭ|\A3�nK�ϗ�o����ɢo�D� %��~��s��	~��⟸)�P�D�ȕ����t��ۘ�ͧ(�̈ ��P=��a�������ȓ9�;�J1ݴt��oA#�J@��`�<d��@�J��a���<	��~"!1�&�ÒB�R�b���aѻUY�i��"O.L�dBCh-q� ްu��e��&M�<p)�a�=;��_5t�.H�4΂�@�(S��
ox3��_<3Y�����0\O`ۗ�͔4tf
$T/�4�@��աoa��kT�Ӛ#�zԓ�
G+P�vf<�0>�G��1LPt4��Q�7��h@��\ܓQpH@�Ə>��y��CI����!�Dse�)�4�ĸ�%��"T=d��&���`!��<ʖ59 �B��yH�� >8@�c�X�U" Q�A݆�z 갃BG�'Ar�݇�T�	B2U����ڪJ��C�	?)�����#n��:��4t��r��5��6N˭R:Z�Pc�9OP9������v,	e$4*�ʒ�'IJ�!������bŸi�P��^�)���!J5&.�U��'��!��=9:|-+V%��  n!��{���a'�N�͑>e��M��T�����}�X�0P&D�L(�jJ�K�4�K�GS��:"��p��0��Sz���M������[,d>2�jP�Ln�!�U�5;�l�s��>n�����CH�;����'���sUB�<� �68՞��'�2�ę+h�����>�f���'�b��C/\^|��, *1�jk�'k�8XÍ_<)Lȅ�Rg�*+���
�'ð��!�S�b����bn !m����'���c���:%�n�A5Ou��'1Ԩ���@�Ȍ@%I�|t΁���� �e��.�[h�R�#҄V�usE"O"H�n��7��K��2{Č��"O4��;;�ZUb��N) ]�D"Oܤ�r�O�t�p�Z��P#""O��1�LV�J�������q��)��"O4��`
{$���6r�I��"O�4چ��gu�غ�У7`tE�Q"O�%�� �
f�8l^�{^I1C"O����^SҤ`r!kW'w�y�"O����n�;R��3F������"O�<+6�hT�0)ǰ<����"Or�k�J�8 �����ٝ0  	�"O�,@c`أ":� ����q�H��"O^�C�闇cȑXW��1m(@�"O>�ٳ� 06y�q���K6\!�"O�Ejզ��|�h�#��	 3����"O�1���<S���j����qz)C�"O,@�pC��S�"Y���JJ�AH�"O�� �((���93��%S����"O�0�s� r*>}�7��S3q�t"O�x`N�<W���eDtE����"O���0>nA[�N�ob� D"O����D8#ߐ�a��Г^X^"O��rP�'��ڂnԜ8S`�R"O� c$��j�5�0� �9D���"OB��� �$1�u�î�f/��#�"O �Q�íw�b��5`͋�"O��i�f�P��$�FئRА�"O(���j��+/�PV�,6��"O�t���Ĕ,vT(�n�9?JM8"O��oM8��R��-g��#!"O�QK�	�Aa`��AZ��a"O.��$�4I1:I%�n I�"O��J�-�(i�|Q�&��0�0��u"O
,���&�� B�E�3k�A�"O2p���T�0X�K6�ڮg�^r��'�uꀱi�f(ʓ�˚Q4 ��-�>Z��K�{R[/��O1�<Qrr,��FAS�K��1��	�L����@�Q�S�'M��h`斥&a�����ZH�r�مMe��̒��Lv�6I�A�S/4��� ���(�RIɟNS%�Aʖ�`��-�%%�����t�Q�d�+���s?%>��}:�@�<܄���I/M��C�l�aLؓ�@M���ٳc a�t��,1a𜩂��bE"���2�2SV��rP�R��xb>��W�{j�Q&��X=�f��y�'�g6@@@��2e��������v����Ӂ؛O�U�w�\��X�H7	��>��٤NQ�z���9a5�'A2x�&fր<�t��2D��}��� Q���hfn��?�M��R3���<��^��FMпt ��B1�Ɔs:%rVf�k��{2>�������)�/��O�T r�'	0*���#:B\d��'}���B�,m�p!�cD�>E�����_1ȡ��W�iI��B"E�-T��U;�re�քYp?��ӊ1<�$�� ~�ȡA�f�/޾�8��AJ���7;O��آm+�h�9����wӠ��݋MVfQ�r�a�0�[�4@�j�[�I�-(_���i����!j�@��JпA� q#���y�	5n��;�
5f��Q����(�l�V@+V�(@�.�����Nơj,�B-O?7��
.mĐ�Pg�%*|`�
L�J �����q�L�J>�Ϙ�j�O���faD-�$S���C�<��鉄Bc����!F��ږ�@�<���\3 @  �