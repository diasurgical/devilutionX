MPQ    �    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h�F����|I�,N���
��8J߬�Q��᧕� ?R�vl�+�ꗍKJ8J�����.m��j����v�fմ�o.� Q�zMd��g�F���L�7¬��C~#p/�p}��N���*��gVW*i||l��_�t�;N(���:�HB2 �ܴ"���>��q6�)�˜L���i�v�X�h˸�Z'����4�N���z*zFAS��]��:쪹~ꡚ��HD�07n�Rv�b[I� a ��)�6�"���i�tI��X5 �0��n�!�0�������v#����q�>d7RN��D���5�<����˶�^����_�I�]Cs:����_a�Ʊ��Z�7��j�!J��0UE��)qFϵ�ra{��Y�	���2��V3y<��پ����z���!�<�E�iς�A�1�s�Wٹ�q'�qV�,���k�P����]׬���j��Ϗ� p�ɻ�3��S�;Y���w~;W�D���M�]g�� ��t��5rY>o�,c��wt7�X����S����a<����}�5C��}�����^t�����޸�U7+���>�V����:,��1|n)_w�>M8�/9L�&AJQ��b ��C��a��s��)¦3A�T�X�0VZ2��e�)�#�Y�_Bq6�9#Λ�Đϰ����_�k5.y��l8�O�ꬃF��ry����Y�u$S'"Q��:��|��or��K�M5�M�X��0�T2����˶��e���(Yt����?h�T�۽�7�m�$) D>����z��{QQ��Um�����X��}Ty�G�)J#~�r�H;0$.O�*
����4Y���h9M�����~��j@��C���N����LKStt����R)C�xE���4��h��'o�,�����L�tJ�o������Q�3�u�z1Ev�@�G����PV�u�u�0��� ��1��Q�aZ�LE Ψ���R�˪��4骀v��:�MS���ůӐ��"ry�O�&���3��%-m��	�z3���/b�.���f�|c,���d��TO���$�+���"��J�P:��6� ��ߛ�U-R�������8��?Ԑ͗��9=�ES��غ��nӡ>�5M�`�m;as����f`!�����]�~��ر��͢ڞ\�7_Z���rx��@)5�>Z��0ő�t����'h�Vj�o��o�����L+0F@����b����xo}C�>�|������&V���?Q��Cp4X�]2��J�������]][�0 ��J�hMR�@���BAU��P����R��m�3��;��xli����G]��ͳ�T	���S�.�z�a�؃}^���
0��"��ZdT32WȦM3����	@�����х,��H�ir��x�~�����r�P~��/EVE�߼,G���m�)�9$jAU��e��o21�ڑ<��F/��\��Z�H!���{��h���n��A`��P/�βF�f�v�(��曄��4��ƚ�r�vW\ҡ��ׇ���-:&=�F�ƺ�j/�SW�1�rk����2��X�=�ȕI��({}	2�V�R(�i��~Qa>��� ���s�,�,����3���P�4����,��Y�O��A��"[�.I��H��-L����K�
��C�d#B�������WU�&�SA� �t�~R��Gw4��=KF���,�v����0���(�'��� ���5�l�1�j_R�������'�;h��ϒ����>R�x���z`z-W��Yy��Y�zV.Z��԰�#�n 4h%N�w���0� mf[����@1��yPD}�DB��eZL�V��\�����k[ຏ$�x b5P��R�
r��gք�"�.�#���وOc��'֫WD�&���d�-��%F�>���qf�čQNJU�'��2�HtO
zg%]�C�$�����P
��(��7*����4=y}�ڈ���h�c��`���Ӥ_�/\w���k�<b��Nr��g8I%le�_��&򖉃
/L��?�0��h�j���(��: &~���ˡQ�_�`�[���v��B8۾�)�h|+t�ã���<l�&X�!�e=�F��� ���,��$�d/
��.s�B�� ��*�Z ��o���R�K)���8�<9��}�NI�t-ꀃ�8sߣrѮ����UxD��Q�z���72����墎i��F��A�￁\������D��K^��$b�Gc e%��3�C���a�&����޽[K�N��������5��JZ��Uё���n7|�T
z�ޒ�6�Ԗ���X/X��=U�)������":�'*�= x��$��f�Ļ�N�n��3�3蹛�
^Dd2�i��A�Uv:���pWŢ�.T�1�R�6j$3�|R���{J-�`ߧ�w-`)�b�f�N�bN��#$>?2��z��R����BgK��6�t�7x̒��N�oe�Wm�d;�,��y*>t9B�U��j�fw��SD[��Ψ`-NL8~m:�ȗ���e��N��,j-h9�tǠp�a3�9�t?�- ���L��Ѥ�A&��YF�u.��i�MDCc\`w�OSl2+�wz�]?8Oƴ���������a�3dp����P�P�<�H>j��;����$C��|L����e�1=!�M l_���1څ:����{4^-r'��F R5%yw\�?�%��sW���9L�qH�h��|'@^�p �3瓫���:m�_���t�T�l���	<��%�%��鿲5�Fʐr[dpC�̅�ۉbN*������������I�u��#�� �����6i�.�IV�kp(hǚYd����Ԧ��,&gJ����B�������׊�]�C�M�q�{ו�˳mA�F��䧘!�ޚ�3M�U��2H��|3v��, z���ihC=�J���n�o�d���7b�9�"�Q�RեԢd'r�b�b�z�A���ܯf�Q�Y��Q�]�&ўp�O�r&�%��I�}�|���N0?!��~��um��wr�5F�:ӄ*7��v�^�孑h�?���+<T5�:u� R�Sl��wp�?uTcM@ڲ�RppV{H#~ JF��������K�-)�&|�۾��������OO�p2��e\�!���� 6y��i�3����{���E��*�Nl�އ_ �X;Ih�7NH�� ��6"n����uqq��fT��ό��t�XX�:��ӛ�'j9��uo�4�	�9��%�uA��]���ű���_��D�ʼ7	3+M��b��� ���DiO��=��D�RI�e�X�-��+��nK�60s���Y��}��[���dҵ����ݟ�5����
�����g�9�/���b��X��:=�E�}l���U
�ս΅w�{!���0�L"����F*��-��{�! ׁ{���o�0�<s�8������U��WK��7��c�l�M�����l*i̀s��Em��\P���]��]�~AJ���=uWW���S���%�~�_���鑖X�H�R�4��y�t��Yr���Ѱ̲�D��\���P�b�8�Y��3R�]g5�[�Ѹ������^oy��׸�/1+�/,��I�V����uk2��3�n$Yz������|�L	#J�/�b��e� ����VVs�Y����C�X��Z��@�q�^ꤸ�>'6�ɘ��`쐊+�ĥ_a��.T��ls,�ą�F�P
y�x)��O$n�+"�2:�0�|V�/ooK�s�����XU��0���2=�������cf}o޳��jhdp$�؅�7do��@Dyz�F#2�7�Q?;�mF�J�ڗ���>%�rT�}oG&=4#�rW��0�E�j[�
et���	�Y�jh�ˎ����~��j@F�5��g�ɉaޱ�w���t�����k)�e�E�<Y�O�e��*���),��GY��G��JWfq��6�Q����P�y1�.�@M8����V�P05ۋ�爊�l� ���L�*�Σ2�_³H��4D��yT��!Z�o[sӋ��"͆x�
�箺<tm��	F��ΰ��*v�."���!�cG�D�P�͎/�r̺�V$�Se��v��sR���.�QN����0�2��r Ϡ���rV���	��Tΐ�CӒ�l�E.8��0�V`,n�BAJ��>";|
?� }f�)�����
�~�	��DI�]i\޹nZC��rS#��{9<��q��+Н�b�<�VVbh�z�j4�P��5����筘Fz8�g?u�ؖ��Fo��>͆S|NԂ�IV�� �i�奷�4s$2s�/J~1_���u[��#�96|h��@�#\B�FZ�+'x��/t��1�.O��kx'KF����G��r��TD 1�s��.�|�a��}{��
�t�"�c|d���Wc@�3�o��vz@��R���LX�Ͷj>i��x!�D��^��IkP9/N�J��+n,��̈́ls����9,tU�������ꚶ��Q�<%;�/���W�0Z�52���+���L0�I�A�^�P�:Uέ?�f��(S���l�����u����\mR���K�r-��üa|#�2��.�����'�ʋ2���Mw1Ȱ��ʃ�k}�U��5�({��y�->St u�Es��ϧdǞh���B4v�ܶ�Q�鴙lo���j���X��y���h�H�ms5�F�
� �������+?�U�-Q�n 4<~Mn���؞q�Ka�����(vc[!�ks��:ߎ"7@�[$��җl�9wj���t&��n�����r��e�����x��^z�l�-28ɔZ1���AV) ��~���	
#�L �	!NfH'�� ��sfV��
��z�D��bB:�<Z'C��S�G�lkV�����x�~�P�R�������}���.Yf�W�k�
`�Bu6W�@�&qaid/;���@>���q���5�e���w�2��{t�"ng�|C�7��=�PŨk(*S)�ݟ\�y����������)	`L�ӿ�~/��M��>�<��?��gq�I�4�e����9�N�8�
���LP��?A����jv�(�� A�(踵b��Q֣ `g'����v-8����D���o�֞wlS��!b�!G�_=H�L�-�ʉ{x�gF�$��ʫ��)HB/V� ����u4��0�-�)� �8HI����N�4��t�����
���B�� DSTx�u����b�G���Nd�	�w��t�����Zdb���VvMز셰��}���e  �*#c1����b�&#�A
l[f[·N���]�����О�!J��dc�%�|��z��6�e�N��O���R^����n����v��������=ۣ)�_BU�!��f�&���_��� $3y���^;���J����-v5�f����]�T݀R!H�j�䬷�*{E%cʻ֬��Y�`D�6b�A��{+�����>��8����	��g�r�6Z�t:k�-�N��Y���n�4=,���*��jB������*w=2RS	����Fh`���8�h�:z'�����7��=�(�H��j�pp��T��?צ��fLؠȤ�&rsY���u锅�:YBN�P\�v�O�R�+��zAW�8
����r�ś'>a1>�p$'�K]��n`H���	b6^����$~��|�lc���J1�pvM��;�놕� ���i4�M'�	R�a�R���4=��Z=�q����+d9���H5���w'^C {�������:�_�+��TPj8�`�	�k�%��� =
�����k������g�ۄ��*���e`������yKZu��x�Y� N�x��46�#�Huk�Q���T��q���O&,��*��	��F��v=ό���hD��+g�:��0�b�h�F8.���~�<ږ����M��:�J���n��v�j�{!�Ж�<CX���}��n��9��)�:��4Jg���%�`��dBG�b(ۥzٙ�����m�Tڬ���yp��r��D%����)�Зi�N+H��9�-�0:\-��w���Fc��e�Lܺ6!^й����ͭR��<o� :��R��Z��0�ڠcH���tp+��H>��J��@���'�.��ȿ�&wd־ M݀Ҙ �	��Oe`��u�\3�`�C��6t�i�ۅL'3�}���*g�#l�_�-�;D���;H}�' �@a"����8q�mI�,\��Wk�ϪX|�����j'�	��PO4	崌�ߋ ��A	S�]N�h���hꗱ:>�D4��7��HH\b*� ���_lp����0�I2W�XBF��&��n�X20.���G��lf���<a�dm9����8vU5X`��%tL�w�d��3j��Q��S��:����8������P҅R��!���0��w��#�F����j{��n��@�^�&��M�<a/��.��n	jZ�r���_j�������[���gM�'�Т{�������]���U�q�䌆�+�lS�=-S�������~�ؼ��x��ΖSq&ɭ���]�t��rO�Ҋ�^`���忎�w���h��a�+�N[ɂ�pn5Д��Q;�4��^jkg�Z2��s)�+�`��4��V�mE���|�gzPns١��ܽ�pL$?UJGφb���;�v��+s�>��\Ѐ�S]XBZ(��ʩ�_��[u6�y��Q4�E�/ߗ�_ܶ�./��l���� ��F��]yCS���m$��"G�p:���|��o�a�Kӹ����XI0��B2��m!��Gr��Ùj�[�P6h���87�z]���D�������Q���m�,��5��N���BT�)�G�pV#�r�5v0������
� ʽ�E�Y�!Choj���c�~W<J@s��ND�!ތ�6¯�t����� )�A�E;�1�j4K�^m;��r�,Uz����B� Ji^�,���QF�G���+�1��@��)��o�Vf�8�ɋ5��co�G�@�� �L{u�Ξ��`�}�J��T��v�����X�
/ӆU"(��ş��&�1����m�B�	��Ziі�%��.}H���Mcb�¿˷
�
�F����$T�֦�u,��0���m��l/ ��ȯ�5��8���;���<���F�g���x�/��E	K@�N�@���?nɫ��~1����;�����f�Ǥ:3�4��~�i�E���PW\�[&Z��{r.�&��iw�t�9�&�eҽh
�,�h�Aj�����&�$��ȂP�Fu����h��8�\�os�>�q�|IR ��dV�D}�����r�M4�r�2�o�JY�R�<^%�.�[�(c��A�h��@�q�B7X%�h���I�`)d��B�x�L���GSX��k�T�P�ћ.���aK{X}�_+%
&P"���d���W��z3�\тs�@}����e�J�͑��i�aGx����J��(�P�Ѵ�e$;i��e�P,�q���9��U>��Ͻ��e#���F<`Ν/O�,R0�ZZC�?Z����z�^ T�$5�A��JPe��ΨXfg��(`ś�jF�*�
�P�L�h\#���/6q2�-���|"���6�	-4�y3��w��:g2I�3��0��K���p�}������(���t%V>�-U 0�ts~��"dB�C�s�P�{4�.���~�*c��1ѡ���e�T\T죒Y��`�Av
@����[��m���<Ubr����1 �#S~HIA�ˤ�Y��K|닧"~ v>K���^("�n�ݹ����ݫ�l�aTjUKj����Q�)�q�4��T��>�3��i<x��zV��-Wn��[0؏� V$\��S:̰�0�#�JH*�HNA9G���:�fQ��e햵5�kD�l�B��_Zߏ�k��ԇkQ�y�E'�x��?P
�qR5��w���j�X_�.�$Ʋ����9�]4IW:�f&LS(djh��[σ>�fwqA9�ǇX��Ne�2ebt�Z�g[�6C�j�TЗP��(/��*�a�z��y�V��)>�����`v���?/R^��^1�<���}*���I�Dea۾�TP��
�1�L��?�f�pjk��(rb� \
����==dQ�`)���v�U�8Q���_crԺ�yk�N��l��<��K!��=P��1Y;�+0�B�o$Y9�em��$=�B�� l�ؐ.2�e��B�)7�{8�uն��N������Uߙ�ﮜ����xmD��V�p��p�E�}��<���j���d�.X`��f@��hD����m��ʹ��=�1e�JFe���Ď��&~Z���U�[�>�����S �Qx�/�]����G���^��|�?z]��@Xa�ǎ�����&��ݰwL�5+��=��Pٚ	f�Ef��!.�^�k3���	�^�1���@�w~v0��&���d�T��R��Xj�G�����/��{@=E��ш�\�`_G�b�a��r�������>�֓߄��}��?�gA[�65�Ntu����&,N��*�(U��L�,���*4��B^{����bw���S��Uߧ`�u-8��:��`�mJ�A���m\#�s�*.(p:���o�p?��yx��L�s�!�$&�4Y���u�N��+u�V���i\֕O�Y|+Э�z�p�8�/q���o{�vv�alh�p�~��FP�ɤ�H��X�$)K�p��z$��V|�Il��%o1��(Mv<�9��{R��4ԍ�'BQ����R�9��"Z�u�����m�q{�9��HЭ
�r�^p�f 6�����0d���L�fuT�O�1�	�[�%P�w��\�+_|�F�B��w��z�*B�a� �%��$��l;ut~ �7 ����Q6j���Y&k���ǐ��pm���/,\c��;=�����1��8)Ȋ��V���p����bq�cߔ���ZZ�W�֚�/M���,��	��v�2�����Q�5Cs�����nӛ3���0�V��/�g��8�0Ad]<Lb�s]z�AF��#����a�Oc���?��B�p��r��%�b����I�2�iN&q/��W���HT�wh XF>=���i�U�^˭�p����<���:k^SRw���ࣇu��cC���vo�p�	zHY��J<W#��Gc�i`ècv&r�,�[���!�$H(O�o(�t\n�����6oE�i=��������;TD*B5	lA��_V��;?(���8HH8� �3"d�!�� ,q�]���#x��B�*�X7F��	�'`�x�+O}4DఌoB<iAd�e]	�������;Do�27?�^C�+blʃ �Æ�z����*E����Imh�X�~y�!3n$�0�O��Uk��7�ή=Y"�
dݘ��).�l�5"��@mV������8��!0`�N��:�����p�����lA�-D!��0& E���rF�:�Bh{�E�w��9����2<�E���� �ɀ�%�1��jN��g��Ҽ�����(h3�b����n�]ͨ����
]hT(��*w�O��9��Ѯ�d�S�.�,�~̶���;�R�NJ ����>a�t⑺r�y�����(P�)^Z�~F��+�ϭ�i�h�S��5��"�.�w�ϔU^eڑ����.Cq+�n��<Vgq���I���>n���OY��`��L?{�J�b����v�R�2�ws�Cj·���I�XF�Z����r2���w�0�[6�IXάߛ� �����_Wc.
��l�LgĻC�F�fmy�M$�$���"�>{:�p|�1EoCt�K�ƚ^"oX��0۬�2���H|���(D��A�e  ���>h���7�W��2D���|�M��Q��m�s������!.��,T*�<G\İ#s�rܳ0U	���
[�����Y8�=h
)�����~�
@�oų+pH��M�g����&tE+3��?)T>/E�+ԅ�����X�$�,�g�}b�=հJą���J�l����9��{1��@��Ӿ�b�V�a�P��Pn[�~[��"԰�UL�/Ι���j,8尬��������X�������Ӂ�6"�����Sx�A��2q�mq��	�Ѩ�� �3.���B+c}�h�F�s�����0ˬ$����)/S��7���0�����c�s�Z��腫�&:�I	d�"�n�����+�E�8�	E��C�n�`��ңȑݗ;��h��rf���V��é~��[��#��Ӻi\�Z9��r	m�����!F����!�h�bj*3_/h�_>e��Fp"��ʼ�������o�>�|-|��fԸ"xV�%�����-�4���2iVqJ4}֌w�P��[}Ծ��l~h~��@���B����Ȃ�=Ӡ�$�ŶL��x�n��3K�G���^wKT�D��? .���a���}���FO
��8"g��d��W���3�iw�ήI@84	�jB]&�l�i#��xW���"����jP��?À3����@�b,�A�������95�U�Z����#���%���<���/꽌M�Z�pt�2����L��d����A�%P &�Σ��f��(�����E(��#(�+�>r�\����3t̵�-k�����T�(�{���*9NC ��	�2�JA��J������yE1}��.�(�]��o��>	m 듇s2Oϝ�)� ?܋��4��������j����m�LX�xƪ/��އ~ߣ�$�<D�
��:ȕ���;�!�1U=�7��) j+K~CD:X&����K�H$��~�v[��i���Վ����f�l	�jЖ؂��%Č�X��F���♦3�o%2x-�z�yP-�4�
}��*'V�����Fw4#i����NJ�?9��պfL�����i����D�uvB0��Zݚ�B��}��kL�P��XFxQ�P%|8R����F̡=L���.�_�m�����x�W��]&'e�d��m���^>��qwȣ����Sx�r2@�t ��g�C�ؒ���P;�(Je:*I� �U�y.����"���t��`��R��߇/�{�9D�<wR������I6%e�4�o۷��<
��LƐM?w��|$bjƼ�(-� w�g;ѵ��QL�y`����v�8���zfL�X��T��ZlP ���4!���=�0�L���S��$��; O��R�B�[ ''Yثe����>���)rKy8~�޽	NZ�{^�o�?B�C��w���)�D����k����hh�z�1I�������j�i?���޾��(���m����e����g�Վ��&ٺc��T[�·DX���i	ČI������Ѣ[����|_z��k�$�G� �)��bi�:�z�2�[�-���_�=�[H���J�W�f�J��_^���39Fl�|0�^�HW���LFv+z���ȍ���=T�R�j�	x�-���8%{;u��q%�D�`z�ob���t5�(�P�>�U��AM��+oޤ)g�cU6��t�M�c�)N�yׁh�����	,A*��B9>��wsݹS��좰�g`^9�8Ͼ�:pD��^۔�Yj'�Q��4���\p��W㊵*?�xS�nLN�Ҥ�lj&�1YW�<u_(�=O�F�NR\�O$��+˧Lz���8��%,~h���Q�.a��pZ>�Aǉ�$	�Ho��?�T;�杮�$�--|F���/1No�M1|`�!U����vӽ4��'ݸ���RF���(?萗^�g5��L��9�w�Hk��m9�^��� 񅼓�L"�c�����wuT��^�
"�	Ml�%�6C���U)�!d�����<�z6�*���ۍn���z�o�HuO�3[R� ��ꞡ"�6z�'�z��k�����K�2�W^,��󮖍��SId���S}\�^�u�Ԙj�"_7�fL��^������\9�r8����MZK����3���v��1����RC��w�s�hn��]�z�p��*�$�b���֍�dxQ�b,�z�	A�8�ۯ7�-�J���b��W+mp��Lr��d%m���.�^��tN!����W���c?|w�N�F4J��b���^��=�y˭ȕ"<�WZ:��.RRNH�V�ˇXc>};��-�p��HtaLJ�;R���n��O=��L�&m�߾���H�&�?��O[����^\����yK6j�(i���F��'\��j*��l|�X_�f?;:h#�HxuH�,� %�"�p�ժ�Oq"n9�7;L��M]��_AX����$��'�
�oI4� �
�Z-A�]�]�8'�Z��H��+D��7ڛl>:�bǊ� M�������ў���MI��Xx�|�r�n\
0��ţ�O�b)7Ή^]۶d�����`���5�c�[���m�B����I�ˎ��I�^:N���R>�2C�F����!6j�0������kF;�^:�{����-����B��<DJ待>�$��?��DL�U�^���i�k���v�]�H�gL�c��K���rb]C̅��w6z��g�"�j�O<S<�����~���0���Y1�IC��c�s����t�,�rExf���o�c���U�y
��sb���\���G0���5�f��iZh�j�X^`i���?��|�+#|�*��VB�є&��g�n�����k7LZ�	J=n�b��֤�,"���<s�h���_���X9�NZ���쪩������6�9���#��[��_ҁ�.���l$��V�F�!9y�g2�E�v$��,"=�Q:�@�|��oަbKɥ���ghX�
�0��2v���#�����4ߺ`q����h����)��7�^� D*�����+uQP��mwz��+�P�D�����Te�1G�7C#�Y�rh��0�o�V�
����~�Ys�h����~��@w�c�F$�:���B��8��t�t7����)�ZlE���ԠR��TR���,�t���8�Jͅ����
'�=�����11�@6�u�V�as�k���sݶ��p�M'L�j�Δl@#�-{��ŪlD¦+9L��@܎�|�a"�w�;'�\hP���mL�	�
��rіr�.3��R��c��6��������kf$�Vb���&لM��<!���Q`��1�����ܮ ��q[��0���Ra��R�9��%��E�(!��c=�'��n�55RG�L�X;͏I���rf�G������j�~��j��͎E�\/ �Z���r�A�,*���x���*�s�e��7�h�Lj�qV:�����&ȸ��FkX��x�p�NZ
�"oiqo>^�B|�>!�Sp�V�&k�z ���2<4Ę�2�\$JSꌲ`��O[x�6�J��h9mp@n�B-�?��I�x��Q<
r۶��xX��N�JGIq�9��T���Dμ.�B�a��}J�Xa�M
ˍ"B��d@<,W4͈3ܖ��){�@�j d���<�G��i^�x�P���=���Pjw�Ûm�1D��Ӥ,3�Ȅ=��u�9�3�U��*��h�[��|y<<�TE/���H,[Z���+�����T'`��:AL�tP���Ξ�f�G(�G���@� �Q��fy[�\>$P��W�'Yn-&�0���)��P�ҿ��tB�ޙ����2��~�{��2��9}u��B��(LD	�jy�>d e ��~sM�*��|��.��ƹ�4GL;���Ŧ���/�g��󗲪
�?����>I��7��
�#x�PN�r
��_�U\��?V S�~>_�����bCK�ń��v􊍴��X���A�l�G�!e5l$�jK3�]���������P���[��v��*�x#�fzL0�-�B��E���ŏ'V4��	D��?#� �N�z��z��p�[fGG������D�lB�'�Z�v	�}���2�kG������x��P@�gRD�v��S�!���:.���h�"�;����W0��&��d�"3����>���q�o.�=���=J�2��t;+�g���C�0h�
USP��G(e:v*�2��0�ryi=��_�(�
ў��,`}�>���/H���wQ<N
����˟I�Mne�"/����
��-L*a?s[w��j!�(�� �C����.�Q�0�`8J/��<�v>2$8�%$���}h�1�/�V�Ķl���@z!XK�=y�w�gX��������$ύ��P���B@s# ��Ƽ��[��5�)��8/Ҷٽ�N����"��ߏȾ�R�|�A��D${<�f�E�&�#IC�Lv��z�I�s�����q�+̄��tg���U��A�3�e�@K�u�:ގ�%/&4;N�rM�[�N����}����:�e����Ey��w��	O|9Mz�H����Ԃ����}��zY��ذ�ot�H�<�\O=l�����hf����n��&�3T
���w�^��U!H����v&թ��JŎ��T..�R���j��Y�h�e�{6����||����`�[�b�yO�N/���!�>�
��I�U�>���)\g7��6��t�D<��;�N�g`��bB�Pޅ,+�&**��B!��V�.w��S�g�p�`8�=:�Z�9io���S��.����0p�\���?��.�L�=�WH�&�jY��u"�0n���4�2\L4�O��&+���zR�8;�G��㎨�,t�a�up����<�?��oH*�ڻZ�%��x�p$/�|�bF��e�1��M���<���qPZ�Q��4Jn/'x@��r1R��DeNh�t��⵴�'{ 98'Hs��h^&�� �6!��&۶��Hw���T!#f�3�	���%�T�Q��!l���IjP5-�8��u�*�iD�T[�A ���u*���� �����|6�VP�5��k܌EǆK�&ŜԒ�,�!ܮ��������sŌn�X��� ��T�]!^�V��Y9�Wm���������4\M5ݷ�����?��v�" ��>��t�C�ן��n����PR@���%c����Ց�d���b�1zj�sʃ��!ҋEڽp��4zp
�r��%Hh��i���h*�N#.�J�,�a�B~Jjw^��F�q�\_܋8�^����Զ9���g<�MC:a�6R-7G��ȧ���uc9|)�,>p\=�H�B�J2@��bOJ��^���C�&hb�	����Z��O���gґ\��U��I6eO�i�D2�}r�ޗ1i*��l��_�3g;5�D����H�w� ��"ZVcՅ*�q]����r���xp���X��p�?`'V;Y��e4�6���g��AC]���1���8˞�D�#y7u�r9��b"k� {z��5������lI���XP���+n��0_#�,�[��:��d�Y�7d>�8�ķ�I��5���v�B��Y$ڥ����fݬ�D�?:�^�i���M&&���d���!q�g0\sH�{��F�3,R,{!���m����;��}e�<�n������������>���ò�vv�X��^gr�Xv�8Jj��<=��0��~]d3���t]�絕}̆���S���~��kX���V�D\�ɾ��ȝt�;r��B�s��̞�B�_�g�t�Z��ŝ�E+�����IM�5a�UѤ��^[��k}8����+#�ч�[�V�ϔa�T�8$n�����OqLuS�J�mbf~ܤ���h�ys����mi'��B�XT��Z�*9��3�J��fq�6�I��b�ːvV�0.�_M�.�	�l_�����(F���yT��� a$�h"���:a0�|B�oy��K�Ks���XA�0�b2�*8������[�Ϝ�[�<�a�hP��D�7�}pkFeDe������g�Q�h�m2���F������dvT���G��#�`�rÈo0�L��?n
Q毽Y��Y��h@���y�~h*@2��a�s�'��'s�"t{޳��Y�)
��El��Ի,���7�n�p,�����3��Jz4{]okࢴ�����W1lOA@�EP�z��Vwr�-��x��t�ƶ�C��j3LL�Ώj�q�y����8u����y�t�
���2�wP�"9hw���w��(��m'��	2d:���.�"�� �c�*-�<�Ɏ�4�̦s�$%B|��2~�ߋ��*B���l���������o�v���Z����>��矐T4ג�j7E������)�¦Jn�*)�ۈ��;覲���ff����iT��~I�V���I��\J>Z/��r�6��g�a�En�<'����Bm�h9o�j FO۹�T<�S��Ff����Ԅ�	�%��o�L�>9��|��O��݆V�G܉�@:��~y4�[�2_��J�H�����X�[s�ʪ�#h�C�@&�B�L����M��`��3)-��x�i]RG�-��T0}���|�.��za\_�}n�|7�
��N"cd{MW���3��7��g@���
8���"2�i���x��%��2j�9��P%z�ö����u��,nʄ��qX�X�9�u�UoV�� -v��|��Wq�<H/ S�C�vZk+7pD��,���ZH���(A��7P6�Ιc�fx02(?��\�� ���L�dY\�T�޾�D��-��G���&��Қ�(�V�y5���2Z��9������oN'}P%�}�(�JŦeS�>�= a�Ysh�nϓ"<��}����4����%'� ��[r���ƈ�nB+�����T���%t�2�
Q�����)$��UU� ��zB� ��c~9�`;�؊H�K�b����Pv��Q�W��D-��O��y����l?�\jƍy�8���S�B�R��g��Og�����x>�#z�-��qɀ��`OVл�d,p��d�#:����N��ǌ��J���fBo͙v`P�f�SD�B&��Z�r���pF����kB��VQx�1�P[��R�PQtE��!�)\4.��I�Å�������1�W���&���d��,�>~^�q-7ٍ�?��G����2���tv�Gg,;C�ó�eGP���(�/z*?�9�<Hy��F����h��*��`8p��+�1/èX���R<��5�U~&��oI�Ce�v���QA��1�
a��L<�?�S�r�;j|��(��� ��F���װQ���`ӕ���bv���8����������
����l�m��!�j=4Σ̂��u���Ӂ$
h�6r�ܪB�g� ����3]��[}����)���8�������N����Ã=��
n��-8��|�D�rC�av+��Ko��O�g�0���ҺN�h������.���*H2؞������L7el��|��ߎئI&�۸�-�M[�'�:E�X���L� &�����Xҽ�@o|T[<z}qQ����Խ s�_!��up�������1Q�c����xc=G���K���f��e�%^��s�3o���r��^��u��S��H?v!���7A�I�TI��RR'j\�K��DC� �{1E��'���$�`�Ibvw�*oi��w���qB>�M֤f������Vg��'6�st&�̙��N�uŁ0I�Wf,FA*�hB�#���M�w�S�@:�fhg`� �8��:f���ډ����|\��;8�pk���a?���	e7Lı���C�&n�Y7�u�;!K�-ETo�6�\���OZ- +���z�|�8��:b��^N��#�a��p��5�7�q��1�H���u>�J0��SB$j8|S��|5�1� M���W�����,�/4��'���R��� ����q��]V��+�9s��H����c�[^�� g�2������������T��e� d�	��%��i�lɄ������O������-�p�*S��Q;��3���e��uǮ��~ �-=���l60�8��N�k�5���!����D,-����2�	�Y�bp������T�����.�yלn�T�5�i���K��Țu�DM���6�5��#�v�J����Ђ��CĀޟi��ndRB��J��� Vҹ#��L�-d���b�LzE�&����m�N�@=����\�p%P�r� 5%#������ ^N��楈רIB�u`w�KfF���Qu8�&y�^�I*�/�H�>�P<�cT:܊jR@����7�F�
c4�S��
�p�H�C�J�d��=�����4ZD&cLY�l2���+��u�WOQ^DB1�\崯�6`:iN�O�8�9�[�#\*��l���_' ';0H��V0Hi�� 7��"�[��`�&q����m����?�;�rXh�>�Z��'ы{���4����@*�IAu�A]:v�Lj�_u��[D �J7�p4܂b}k� Æ��˸E�~v��GI\{X������nFb0�$�G@��Xl��? bӳ+dه��.���5D'�đ%�c�Qڀ��V8 L��?�|:���$���hjq�<c����!�n+0�L~�v��F��>ԉ�{<����K�ʝ���<z���{���ڦ:V����X@�K ղc��������&�S��L�Ў�[�6�|�g]�1�A�KH����#D������S9�,����~]��W#Et�?�v�F�o,�t3Èr;�*�Nֿ��K4��ϒ�o���)IG� ����7��֧5<�w���e�G^V�y��+�_P�+>eo� 0SV�<��������n�`����T�L��^J3��bA�Ҥ'᝗/s���m�z�fXo{{Z�d�@̩�tK��6�y
ν��1q�K�R_�̝.�n<l��SČ�F��y��x����$�uk"3�c:<@|}��ol/K��oR{X�Ko0,%�2lvq��Lu�3�jz�Vsզ�7�h���_E�7x�F�VD�൜MN��ïQD}m���a��:f?�T�8G-#�r��0�)�H�
��4uY�>'h�$���k~�A�@�%L�|�0�Z�������th���/)e��E'�����1�J���I�j,A�CN���.jJջ��1�~��32��QG1��(@T�"�u� V��Z��,��-���|������͠L���Ί�
̢0i<�S��bk��\19���v'��r9�"�p��.o��^�����mze	m�Փl���.�U��Ⱦ�cΠK��ݶ�v�w����$�MΦ~��:���T�������i�w���$�ϧ������ZE��S��o��:&Eu���:x
�]�>n�?�����<�;ޣ���fA�Ӥ���I�~z)\��a���y\e$�Z�\�r�K���jm�������)����hT|xj�������MFa$z�.
�����@}�o_H�>]�|5��ԉk�V~�I�0�O�^�:4�>}2�ɮJ�^(�!QY[n�z� ��h�:�@A�B#�
�r�;��<���� ��]\UxΓz��G?
��ZBTkd�zK>.�f�a�@�}�z���
�{"��5d� bWj w3�PR��s�@i�96b��T���iԖ"x(zZ��j3���P�����A�'���ь�,��t�s�I�[�9F�3U*��;�K�Q�G�2�r<L[=/�ͽ>�nZƸ(+}��2|3�J�����AµnP�v*Δ�f��(����&�����Ƽ���|\t�H޹�����-����K��U�u�/ꊣ���62����w��7� �ꂔ}+���1.(�q٦`M�>S� bs����g���@�<.�4}O(����{O�b�������0��l�'f�t" �-��
�"S��#A�D����jU����J ;�~4��i���EN�K���@Yv�Jf��K���	�9�"_Eݗf�lZB�jA9���m�=ɞ���L��X��w3��,xY��zB��-y��ɻ������V���g<�wC#U�y�N�<���}9䦕�f=�����c�!��DQ1B� �Zn�Ü���Nek=�����x��Pv�R��:,;j��è��E�.����BH��1���p�W&��&�Z�dV]���a�>yFq�����q�	[>2�Dt�{@g��$C�v���YPl=�(�DF*�����nyߣ%��(���-��%`�XB�F�b/>����<�<āՔ���=<IG��eM���<��x�c
<�Lw�D?HT�m �j�(^�� Ȣr��@���*Q��u`n���_v�8=���I�^����z�:��l!D��t!�=��̝I��(H⮠�$Eb�ѳv�QDB�{� X�����{�Q�n�t�)#��8Oh/���Nk1��
��Xe�߅3>������DZ��\���ܵR�����0��p�'�)�_���a�)˼ W!�Y�)�9U��)�feG�Q�8�׎�G`&ꛣ��Đ[�j~���B�3k��=}��~�����ѳ���J�3|o��z�b������<����ƣp���K�԰c�~�n�	��="_نf��(@$f��5�pf.�J�t3����f�^fM�˥ ��ov�੒����rTd�R�$/j7N�ޡ����{,��ʂ���u�"`��b�i<q��ߏ�!�p>���('���/�g-=C6��ta�4�2N���y����,a��* �5B�F)����wDNS�9[����`�D!8 0�:�߃���ԉ
�h�"pb :��{�p&�A���I?u~��#L�E)��_�&���Yh��u�urf0����eZ�\�RO��1+�U_z/8���}2F�-���� aXQ6p+���2��5�TH�hm�����Z��.��$��(|����w%1_�3Mb���rAa�g��4��F'����ȢRW������Ꭰ��,����9�y�H<�.�^k�^�0� "��M���"��b�R�/TW>]���~	^]*%<,m������xʲu��ך�n���k**����B!�N݃��2yu��t�� U����w�6�������k���||�ܜ���,Ⱦ���C��d����3��9���[�e������7�]�O���F��õ(���M�`��q���u�MvΒ�BF�=��C�
���Fn?����b Ag�iùs��g�d�P�b�5z !���ϯ��;��s������p@�rd%��@���UО��NU� Q�����^wT�-F�M҄�����ٕ^��ʑ�}���Q�<���:W��R�hU�1|��Z�c/ڹ��(�p��H�dJ(����q�Uݣ�ϐ&^V ��{e�y���7O��%��\Z_h�J��6[��i�m���+��'�&*�Al-^�_�,;+�[�Y��H$m Rk"P�U�;��q�^(�B��.˖�^kX#�P�u�A'L�i����40��fT�A�ݠ]����g"����ԛD[�7�$g/�Bb؋� ~�~��[�����fZIY�XI��v�nm�~0�jʣb���ӽ}��P�dt����G��5�h�Ĭ�O��r��[(t��r�ڣ�:Q:_����X�Ѓ�$ҷJ8���!� �0�F,�q�>FL�Q�� {W��c�,�����<�v���5���@���6�Ɲ��>� ��c����N���nf�I���([���k]��~�|�T��ˆݱ�3G��P�ASTR����~8Ǽ��0�ꉖ:�@�t�3�*��tN��r�3�)@�5����՛j��쐨�(8�ՙw�?��5�I��r�;ò^Q֔�!�i��"+Y6U��$�V��<�׆^�n�in���~J�Ly�L���J���b���b�I��`\s����#���5�3X�"�Z�bu�������6��(�]|�쫁f2�_C�	.v�"l��'"�F�y
w|�v{$�6"� �:p�|�ao��YK�������X���0G��2���'H�nAD�x�Q$j��hƶ��z��7�ʹ!2�D�!h�趦�?�Qa?�m�N3�|,���gQ��TgIG�RK#�άry�+0A,r�
G_p�QQY$�rhvc���}�~��@����� @�67���Z�t����0)�o$E⊩����řG�$,u,|\�����)��J0c��t��h��/�r.g1�D@�$��pn�V-���p��F�j}���3���PbL���΅�9'�G$�2�n�p��.�7d���}c�mB�"���lbt��	;��m�W�	�v�pTޖ�2.D����}c�6��27ЎQ&����$[yX�yP�ٕh��m���t]�����R���_� �B�뫹S��qa���ɒ�)�EPe{�u2�����n�t�cdn�}��;5���f���B�y�;��~u)?�a�Ϳ�\�f�Z%��ru�ô�:��{�)��T҄�ϐ�8Yho��j���K�cȉ]�F\�މ_͠��[�'o�c>��"|p�	�$vVy鲉�!�v�4Bt2U0�J����c���i[i�F�[ZhjQ@\�}B����M�ّ)9�"g.����2^x�5���9G�o��4T�k[�:.�(�aB>}{�����
�A"���d�kWz�3���:��@$S�Q�.����ՙi��x�>'����u�P������$�|���,�������~�9�Z�U����V��̭����<���/Vh~9�BZ!fz��P�M���!ݥkcVA��Pl|=Ώ�vf.��(����A� ��]Ɨ�*�3\�޴��8-W�b�A��K�P	�%�A��R㬅�2D��q��RT�e�M}���(�E�[g�>u�� ��s��.ωA���{��w��4Ӷ�Ϭ����q���� �d����=�ʜ��?$�(D�
��ȁ���_�f���U��F��" ։\~/pw�ϟ� tK�V���-v��ʴ�֯)
����}d��RXlu
@j�˂��e�x_��xW?��i!��3�[T2xt9�z�-T����A�ؖ��VhA�è�2�:#p!j�r�N��8�+*��Aɛf8���,M7��D:��B̈́ZI�X�.���8k8�E�^�x=��P��eRuʐ"��Z�_O�.��#�yۈl����ϠW��&���d�*��bֻ>tN�q�%��nk����Q2�R�t�Smgb��C�I��MP'��(�y�*5\�����y�X�0sNۄ���y�`�aZ�a�{/�����ϥ<�o锋�Q��I��ne~6��G�����
'�L��?�t�h4�j2�1(�� ���`���TQ8��`	�]��٘vOm�8��5��*�٪���u��l�:��>s!i�=��̸��kx���$�|l`��YBQ�{ f{��"��p�O�O)^ 98�4B��}NƐ�JU��s�� ���Ah��)�D��y�W�+�7@vTj5���Ǣ�I���U@��S@˷�Ax�e�Q��T�.��#�e"�����Ɏ�s&E|裰W[�"�0�s���x�86��������+��|��zst璇\�3��Ǖ��k����r�W��t��p=�JG���'�Îf�b�����m13�4�h�^A�T�{�~rvn���9�ſ��T��R�jQ`��6={'����Bm�0J�`���blҙ�(���g���pW>�3��Z�o"kJy�g��*6|�ht����ːN��#��*w���S,|��*���B���jHw߳*S�Rx��g`J��8;�3:\�*���_�EOQ��@`
���lp�h�����?�o-�v�L:�X�(��&��Y�3JuKχ��f;��@�\�dO�Z�+��zcϼ8lg���'T-�Ž�Qa��pƖ�-J����H[�<���@�A�	V[$��O|�x��r5K1��M�[܍�������&b4�� 'I���uR��|���F�S�����9�dbH�
��Y�^7�� ���h-~��:�\���� T��L��%f	���%������r��oVʍ�^ٯ�	��ffw*	<I��h��iہ�[�6u���G�2 �4p��~ 6�J�f�k-� ��5��8��C��,c����������������Jq*�@���(���2ųJ�bh��ߘ�t�k��M�R��·��fv��������/C���_w�nl��^�Tl��p��'Y��Dud��b
N�z�hM�$4t���ϋ6���H��C�p[0vr��%��G�;�9�N��[9�����+ew��F������\Z�^�Q���F���<��:ҝVR��d�B�t�|F�c*9\�=g�p��^H�xJ���ʽ��Ln�j�&Y�C�"��45$��OG�s�N�\��ߴ�e6V�;i�����F�{��}*�fwlh��_]Yo;&�Q���kH�l mm)"������q��������H�X��ːw^'ǌ$�r.�4k���v��A+�_]�{U����y��\LD��I7F�U*��b3�� 9�������~�A)I��BX�y{�btn��:0�A�}|q�N/���!�Iqd���|�ZI5��c��*��Y/��6t�̦�7���5�:�Bk��E]ОR@�2Rąt�#!"�0-`R�l(F��dJYq{r�q��������.��<��r�q�?�̊��ԚA;�����	L��/ֵ�I�gI�D��d�C�/�rT�]������~$ǆ�_5����So<_�v�=~���~Y���5g��V���S�ti�:r1��RP�O>Կ01�eZJ�߯z�vWZ��߂�IM5���U�3��^�^L���|袸գy+t'��9�V�d�����	�n����ͽ�wLƇTJ),ob�
����9�s�<3�~���QX���Z
�_=.����7��6�9��s̄�����m_��!.Q�9lN���i�F�M�ye��1a�$+��")A�:�|�i:oJ�\K���%�Xrp0b�2bm��"����搠��L���r��h���ە�7n�����D����?���ZQ�Z�mc�������0���TQ�GcF�#�5~r��)0�!�'��
��B��LqY_�h¸�ׯZ~y�@c?ų�4B&�ޮ�b$�CtL�����)bE������@�!��}�,����)��$}GJ�*�'+��r��)}��M+�1��@���krV���ME�������K�iے�9�wLհ΀$E���ߐ����$�XE��!%E������hk�"J�w�'�����Cm�U{	�/�5h���.�C�>\ c� ����,ϰ�W`T$���t���d�(܄B�x��-Lܚ}���9!���?����e���xߒ9HE+d$��𓫎n����X��8�;9��}V�f�.;�}�*��B�~pI��g�\�z��\��>Z���rP��+!�������F�s�ph���j�s���`���u�$�FWp�����:�v�NoU�>ʒ�|���Կ�aVtj������!J40es2жiJ{�ڌ��W��[d/��%�h%�D@w�Ba��(�'�dU��
 ��)'xD����G5#N���T�s��H .�
�amc�}6��̓�
�"�#�d,EhW��E3Ȋ����Q@�*l�x��ͳ׶iJ�x^#���:��J�PVB��PzZ�Ǝ,C� T��M9���U��1�q�N�G�����<��/�"4��Z|3,�N<�h| �@���Ff�A8R9P�HΊ��f���(p�Û\m�<p�r�\e@\���ޯ'P�&*-f����6m�+bN`S�J����c2k���j�C�mR���KS}�Б.�(�
�V��>�% ��Ds����e*Hܲ"�4������)�1x9��_���8��ުv���2eߪ{�#�
b���<y�z�բ��U����+� q1�~*��ػ��K�קa�v`��������`��؉���+l��j7�Ղ�P�ĳ��)���[�`�����x��z8J�-/���1Q�1rVVd��u>����#�߂��Nc~y�f�2���f3də��ʵ�� DU�B��pZ$&��i����ldk3 �g/�x���P� 5R��R�(��?h ��x�.�C���n�'!���N�WRe&n��d���j�>ov�q>M��)�"&#��2��~t'L�g��lC�<��v��P�X�(��6*�T�ݜ�yU�߈�ݵ�B��;��`i���|�|/4����<:~q�&���/�I�.�e�1A��rL�n}d
�.L��x?~�gc�Uj���(��� ��Bx:�_�.Qs�`�8����v�k8��n�,Tϱ֛����rlWQ��')!�0#=el���s���\�d>4$��5�����B�D �EN�2YQ�G+��*��)�e�8�!���N!��Ѓ�ɽ�{n����-zD���R�E����`��j��fm6��s>�����/˲	ӫ��ю�oe����e����Ncn0����&�|��^��[#QϷ����鶨ĳ?Iя���5��i�R����|�E�z�t�b�C�n5�0̬�fu=�+Ѱ�6���k����h=�VO��T1�^�@f�T��&Io���3�Z���,^���A���L9v{ܩH�@�z�TT�*�R~)�j��T�R��O{"m`�8S��@`|b�/v�5�:/�W �>��Cֵ��*p�e~�g#n�6W;�t�QB�j��N~_�/X��<�`,��U*��B�쁄B(9wz93S拑�w�`�38V��:�<���z��ΘX1vƮLb�p�Wg�T'?k��/Lu�<���&�z�Y�uIa�ro�q�\8�O+!�+�i8z��*8'l	�Jq�LŘ�ra��paȭ�(�����:Hh��s��8��$��|$�me1�M��4ܨ��]f|�C46�.'����Rx}Q%��)����ӝ��'9$pHr}��T׊^�  �9���u�I?�7t�ȦET��4��I	�U%�� ����@�h!{<�X��JM�a��*d�肯w������� u���� ��]����6A�s�!dckH��r=:���f�~2�,���}e� ���&2��\���e�[]�Ij��m���Em3�����Ә�S���~FM�d���O���vĂ��4�г C�ڄ�n�(�<��w�)��ٹ)���}Bd��Lb��iz��ؼ_�l�>�ԋ17]�)&����pv��r���%���U����@N��AبM$Z�swJ��F`����<���^�`�@�5�oo�<,fx:M�R�$�}!�Rc%�:���vpH$�H�8J�����ٙ���^�&T�¾}nV�����00O�l-��\�sK��G�6Q��i_V��iE�a��a*dнl���_���;!���9H��� ���"F,����qI�!�>�:��d�LSX�hA˫�C'B=��M��4�c�2���A�(]k\[�����7�lD�|w7�<%?�b�,� �i��;�u��)�I�o�Xr��non#��0K8��J���������d�R�S���<5uL����|�����>���W��0u]:$��UR�й��ҭy��O� !]�.0ș�g~�F�w��{�y�Y���[���i��<KA��lT����� �/g�����i��DTr����D���cп3O�^p��\�]���b����-x�A���*:S��T��@�~�gj�WA����0 ��*���t��r�P,�߿�̊g���a��`�'�:��1� ��o�53�5͢�ѐ��q�^G������}�+�8���mV�(�M���n����q�0��"BL�kJ��eb�yU��_~��cs���:H��A�X��;Z��/.��6Ըң;6��9��[��b�����_9��.,]�lK��]�FШ9y��C��f�$FM&"��y:�/�|.�go�7K�#����X-��0}��2���j=>����;ӃG懦��h<�۰�(7�3ם�DQ�������Q�m|L������k�yT�_�G�Yi#伋r/b�0�S~B$�
=Xa��haY���h�@���~ԕ�@�׳͈���4މ��_�t��V���)vȟEX���'Ntһ�����,�q~y�e�J��I�]��W��ĕ(H71Xp@%��f��V㚕����`�d�D���t��L��R�{�,����yL������a��)�`��G�t�c��"�Ix��)�㿪�h|m�s�		��5
���.��g��Z�c×�(J���U̒D�$�0�o�4�Kŧ�㑗�)�n��gӚ�z��lL�x���B��k�u��z���$]��h{E����e�.��n�>�mT��[;TC���Чf��������q�!~k�ٱ¿��5��\�J�ZMr+J��S;ɧ��Ń�r�:���.��h�c�j�������ȿBAFRF��?j���]��%^o��>�]>|潓�Z�EVoz�A�����4K�z2K]YJV`���%���[_|3��h��@��B�R���%���ҠX�	EͶn?�x��1��BG�_y�^�T�_�Kw�.{�aȤT}�`���
�0�"��Ldg�YW;�a3�W���X�@�"��ϭ$l�͎��i�NZx�'����7���lP�v�"p$����b��,Z�}�Dpm�$�9W�U[��䌁|��^��Ð�<�T�/���/�~Z� >\���,C�h"�!�DAs��P��K΅�Rf���(+��w��:��M����^\EWrު�6�i�-���9-��
����e�����㢃`2� V�%şȈ���[�}��i��(S�&�Q��>+�^ MP�s�b���r�@����̼4NĐ���"�<WG�5��"ْZ,��Q��@��E�4��
�����S���,�kU_�n�f�@ �5~%�~z��vHK9!�!;v;Z��CM�_O���� �3����cl���j��̂�˦������r����h���+�x��jz��D-
���l�\��z�V�7���a���#�����2N>Oj���=�w�4f.K@���R�DpLuB��Z��󜤍�K�k.��� �x��uP��lRk��Oy�zj�����.����/7��ȡ��W�Ԥ&Ip$d%<���>j��q��ō�Jo=�=zc}2b,dtbdcg���C�O;��P�P�^(�C[*+m=�w�y����fh�� ,����`$Ӷӗ@f/�v%�[U�<u�m���]�؉IX��e~������+�
�L(q?g^�@j�E(�Y� ���3=�:��Q�E�`?���7�v��8nvk�M����v�w��l���1;!zv= �<����aw	�?�r$�D�8��p�By �E%�MP������)��8 .0����N|���J������C�����h�8D+���Mb��}�u+��7���ﺺ�%��^�2��˭B�.�؊rװ� ��z}e���3	~����&��d��q[>�&���Č����lH➩���?�{[Y|��izi�-�=>'ԩ�����s�a��\�ﰔxm���V�z*�=��'�7�����fж������{�V3۾�^�^�q��|\��E�v�������5*�T�y6R�[�j�4���y՟l�Y{e�ʓY���`>�bb���b��u�����L>�t�0B�����g�6^62
t%��!�Ny�򁊥%��y�,���*��'B[oV�}�w�3S�䦢҉h`�o8q��:R���&��ߘ�A� ,����pWf��,:�?�u
L��Ԥ^r�&�iYy��u����C�1fR���\s��O��+�#�z�x8��#J���s�a	�p���#�F�H����6�����$V��|��M�h��1pk�M��1�×V��;��U4q�p'�_��ORh�+�3�2���Iڝn*�9_�.H��O�R^��� S����ݜ/�O���T(���g)	on+%m_���U����5�C�'w;��?�2�\>�*�m�=���7��Q�6uq���;� &�����6��\��Uqkcq�퉋�m��Թ��,���x.�uQ��N����a�@�������m�f��@J��n�w�˘S{�aa_M|� �"�*�F�`v�*S�`�n�C0i��U�1n�M�wkw4��b������8`�dp^b �z�X������v��,u�ڄ#���?�p���ryN�%�&���b�o��Ng�j��Xjb�w���F;�k�=fܒ�c^��T��ŭ*._<G�):�0�Rt��������}�c WU��C�pnH�?J�6���ƙ����U&O4����������HO=\S��\.��IK6L.i�*ƅ$��|R��M�*?Zl�M_�;��j�'HUͣ ��W"������q�o��h_��/֖�}�XT��Ʊ�'���(Τ4�>Ȍ�t
���A�}�]&]��
V�o��Dc7|� �kb�� ����7���W���^wI
aZX������n~3�0O���8��DrQΫ�d��dE֝�J���50������O��k\B�cmF��+7:p%W���Ժ��(� �*�!���0c��boF]ъ��^{����!�6e"䤷�<�J�gn�FDgB�F�J
�7�Ӳ����|!�e&�?������z~�y�x�h�]e;I�-�g�9F���D�����S��1�l�h~�Jd��Ow����+��Ʌ�t�[�t�or'E��M!�ŰĿf�/�[B!ꕖ.����&(��<�5�����s���^BcN�2%U�Kws+�i��Vd���D��?/gn��ơ�*t�}��L���JK�b����o�s�N�4��fQ�X��6Z ��gЩq�Ըm�J6�y,�)��1��)_��U.B�l�.i��X�F�#ny�����$a*J"":��w|i`�o�v�K�i0�ۧ"X�N0��e2X��Exa�����0aB��(9jh�	+��Qa7d�����D������&�svQr�m�BO�ͦ�&,;�
�T��G��L#�c�r��f0r��]��
�̽��!Y�[MhG����s#~/G�@��γ��~�U�di��A�t��+��J)Ѥ�Eb��B���6z굁�,-d����m�JA(��)��x����1�H�@�c��a��V>�~� ҋB��ۦJ�������LSJ��v@�8X�U�o���D�N9i�ȼ�����=��^" ���������n����mn��	Y�AVĖ���.Uc,�y2c:�V��%�‪��H�$,�G�j�٦����;�D��nl��S��|�����-�ƪ��?�����B��E��F�&!��N�n��2t��Ȯ{5;o���sk�f��������~f鐱���%�\��Z�2r�/��k��L�'���ҕ;{��Ylh��1j���\N���<��Z�BFM<)ޚ����h��UoKv >�H�|!���!Vj�׉�b��J�i4f�2�#UJ1�3�h,�s�[ZT�l�h�U�@�b�Bd����ӑ��H��K�K��u�x�ڡ��:�G+��[J�TWA ���b.v.5a#�}����
��i"d1�d�	?W�F�3�D��K�"@U:	��j�^@�i;!i��?x�L���q� <�P�g��=j�դ�=�$,�3>���>���9���U���fr�=�H��(�<8�/'��* �Z2.��?��m�6<����cA�n�P=MG΀��f?
I(��㛒�8�YH�(�8�r�\�'[ޥ�9I�H-��Y�T�q���5��s-֛U���2�2!�����ȣT��֔B}�8j�n�(�K��Lu�>�x� 5 s������N���(��4�գ��>��� ua�	���v��,���{����T!�C
��ȲNh��~��~ �U:K�c� ��6~ ���k�1�HKTT2��tvJٴ~8���M���{��4�݃��l�"�j-'��f��)�U�I0瓝\���4���]x�Qz.�-�eɧ���g�~V����+���c��#��,W�N@�����$�f)R�=�2��}D�5B��,Z�=��ߤ���I�k)�D�2�xn!P�R�p��^���(�0,.�]�Ɗs������5�Wwp&$bddBRz�3��>e&Wq�����'XZ �P�2=�yt��,g39�C��3�,�PX�.(�G*����Rc&y����9��Q�`�;�Ӳ�7/*�&�6H�<���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸�x�rhK9�1�#l����_�)��ToڬrN�'|W�Ds��&�M3�i��P�E�d�F��FB*�@�J�O~6�I覑�	ߓc?F�KE�ַ1�v#p*�8s,Z�9lTA�'8�qEx��ϦIq4hF�w��Ձ��Ýo�,�b��<YAΓ0u��YH�T~�M�&a�l�"����|ج��)(_�f�O�jE�x�`�07M�8-��I� dh�
`�irr�����A'璩
�q��ƲLZX���h[j"�@����� f����X�'ߢ9{�h�2(k�J
>�
]�t"�*m�}j���B�I�"��+�E;�%	�B�	�LR6����4k�4T�$i��oj�C�I�n�F���F- �ѱ��:^��C�Ɉ���R��!+1Xc�6Q/�C�I�Vs��k��'M*���f��a��C䉃D~L��R�4}^�Q�D]�r��B�	��p�Q��ǘV����)zC�E�V$=y=L��dȫ^BC�	%X0�p�E�
2b����	u{�����!Ih����bEy�B���kT6pՆ]h6@��?y��&%A�X,G*�\�r�i�u�`)p!� JfJ�)Y#�M3�̘Ix(с��<!��Q�S`<4$����_�xO^3�LƷ2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  �.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   y  /  D  U  '   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=��J�E�TM�P������PŌP_`��7ju�r�d�O���<�'�?!�Ov�%ʢ���)�-#�E��-�����L9B8��	�}xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�z (PЩH��ɢ(�Zc���a&,O�$
�-ڼ1V�pU猤IV�u����B�ayR�BNj$����n ����ϻ%���OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O�����KO���O�<Fz�O�r]�pc�A�,�̨B��;W��)�1��jm4���?y���?)N>��T���GN��fg�h]$S�E�'*!���><`D��E|B|�f]�p�&��OnTh@�Ƀ ���S��;��L�Q����bi,�Oڤ��E?:���Aץ>k\�s�"O�����E�"��ƀ5h��×����'���e���M����M�@$S���ī�턙ZPyç	hBY�|�Iܟ �'����bĜ�$!DѦ@{u�@��G�Z��1DG�=�2��,�=��E|ҍ��NƤI��ןa�N��A��>(Ҹ���1(n�Q'�X� �	�i2��O�����'�@7�O�6��<��3�! �kUPub$�R�?k  ���,��䟨��\�b��&Z���T+h#�8���;n��B��@���P�h\�>ϐ	��$��>�RE�OD�G=���i'>��'Q��C�I�*�P��N�9��te�'����}����;��)��G#�e�R��-��`�)���HOJ��3g]�DF�YS��)
xѮ�3�ޏ;M�Y�'O^��'v�P����?����?ɉ��DT�p>�M��m���4	߂��'A��'�������(fZ�`�ʊ�u����ǓY\Q��rQ�:������/:j4�����	˟(�ɶW�t��ޟh��ϟ,ק� X����z5�|� , E(5۱矖n"��XSZ���d���g� ��)bH�/MªL��ЫFⴳO��2�X|R�
F�,��*##*�S�v��	$D�Bm���(w����t�@����&�'� Y[������dp�Ȕ��X�������aQ�LH<I�+�E��,����O�p����K?	�K웖fg���|��'�B�O��A�)��mIR��1�T��Ek�0�&p�ڴ�?!��?A*O�)�O��$�U\��
�F�t�q�1�W�Q\��5#װPm����'��Q�p�L�N�<M�&�J0��uv��'	��(Q׍�-~b����ҫR�4�3퉼"��h��X���Gwȕ��H�O����ɦ���xy��'�O�1`�5xq��h��Ձ����"OB��1�P�	cl����M ^V�<B+TI�	��MS����?�p������TG%R���
4.��B�$��?�M>I�S��򤙻G�4Z�'�� �ؔD�8!��ik�=�P��R�qЉ'e�!�d��U$pS'b۱'�If�w�!�X�x�-˗�V�_V$S�GE�Rѡ�D9<	ra��8=��,*�g� 5�H}`���Ȯi��>m���H� ^�4��c�0#6�d	���6�?	�°>����Z?VУ�MrcM���y"N��@5%�! �8�<��IR�yr$�@匰hGN2�~X���Q��yr� }_0:P�H�.�.0X��p<�7�	��R���q1� �F�*pd6�IK��#<ͧ�?�����kP���!�4Ӳ%s$��15!�d� ��أ9�:���`A!�D]�A��e"�-�+���C��G5d`!�	-q]��G�(�#� ��l)!��N�k�^IK#���$Y�f��(�����?U2�	�2�Н�3`e!���$}b��]�B�'Rɧ�'U�0a���@�r�I %c�Qv����d�E`Y���@��$�@L���.���H�*v�=�B�O1���M2V]�2�Uej�a�fIX��5��s���u��bt���1�]�i�=��ɽ%2���'W��eP��W�a�Z�pI�f6���IB��"|�'C�\t씙�eٖH���'�����ٚ���.�?�
�'.�TK���9���J�(L/��LY	�'p���̩A��nB�<��z�'G*�b��)��e���D�	B���q�~�'��Tc��i�#@�H��$�#��5Sd��9D�<���x��I-� s0�Ǘ(xX�2c�#�C䉗'�Nu�1��>�(����I#i�C�	���a�s@`�@�	�y�2B䉏=l��S�H,M�X5��� Q����ĐB�'J&qHt�X���b
*�ƨ��'O^9���4��d�O���h�[�D?PL$Xz2.¸2��Bڀň��K��幒�����ȓA�XSX7`d�1&�Q9p�@цȓ�8��g��*�� �Ƽ	A��ȓ,:TE�����ּ��LBR��p�OXPFz��D��$�Dq�E�A')1�@�È��	<1����ɟ�&���Z(qCD�gg͹ F0+�"Ox�[�&��Xb�uc��'5��0"O��Ѯ�4�t�hO�Np�0"O����G�N&��&*@!Y�T�"O�l!�OTe���N�i�d)w�DK�'�4���o#���v�D#)�D�86�� m��6�'�'l��Y��Ɂ�U8v� ���pf���Ш:D�p@'��(,S��s�#�z����4D�x�B�ң9M�mI'��=w_l� �1D�(xrN�T򔄁1`�*g����a1�� F�/�F�����k\r$�M4=�Q��F�;ڧ�(��"!�
m�z}������)��'r�֧� ���D�һ`JN8a'BA@"z�h0"O1
b���.3��K7@2C0|��"Ob}S���#V;�xQuOþz(�ŉ�"O84�M�!�Ti�##
V�1��'x�<�d��r\2e�1���n�Cw�O|?e�Tp���$�'�rX��:��*��˟,7��Z'�;D�di�lN�9���݉|�T!�
<D����
�Bgn.�Nb4D'D�h�ю�q9�܀0�x���g&D�,����W2�<�" Z��`"�*7}"�?�S��-$�H�Q�ݟ@��x�� �13����O*$
���OL��&�����H�F��'A�R0Y����y���1a�8���O�ay@�yReS�6��1�D.�E� �胅ܽ�y�J�%��pv��=>�R���@W:�y�^�Rĩ�b��/�r|s4�W���'�@"?"@�ß�1�)o>D�`FgK\��4�W�?qN>��S����U�3(H�ID��-p��eƚ7�!�_�yfh���6t'���d�k�!��^�2�� bSd@�x����i��	�!�ЀIЀ��!"�����$�!����h��`h�`�# $:�`TnH �d����9y��>a��㇧Y���BK#
6��u���?�����>�!��E��ى�V�2��� K�<����J�`�b�� �_�<���Ɔ!U}�X�$X&.�MG��r���YB<m��S�u:�p�㉧�(O�h�w��/�<��T�=k@-�"�O���Q�i>9�Il�'Gx���SU���#a�4R��j�'+lx��MA4.�RԐ�@H����'x.ЊvΈ��t��G�K8���'�R��I�
E�H`��Õ?C%��
�'����#�� -M8|�3�!SU�5�N�������3��� ���v�����( )���X���?aN>%?�!�C�}�� �h�3}�*��c�,D�aP��+r ���LǪh$�@�I,D��І�]�_4� B�)�v��|F�)D��0�B�z��/�aX�A�-*D�p��۴�<�Ui\�O`H���'�<��OV\6�' Ƚ��`����4#�)��a��O��O���<�`ac`Tyag��P������h�<��+�B9� �:@ht(�d�<Aң��� 〮L�v�֫D_�<1��H�t�Ќ���ސ:�<����Z(<���߂IA�|z���,u�*��K�'{��>a�X�O�I���a��a��� ~�L��@�O(��?�OH)4H�31�E
ìL�Y�m2"Or`����0^O�Q��Z�G����"O�]tcA	+ :=q�B�z4aG"O���,�h��E����.�>X�`�'�\�<��H�pO �hD�%?��Չ�A?��G�\���T�'_�X��0�׽p���j�DD9TZ92�+D�8�1�� ��A d��1�N��0G/D�@a׬A�@�eQ@|��Dg8D�lp��^_��`�u_�sT�H�k6D����٧s:(�%�O�ya���d�4}��-�S�'dX��h�^vRT" ӑD���OYS��O ��"�����1[�B����z�jL�1N��y�*PW�ƁV�"x�l��j� �y����#��q6k>:j��ֳ�y��;xI��`�#A��&�Z���'�y�+H"	�-p4�˳s�8�����'��"?���П p��^e��P��'//D)ȑ��?iM>��S���D�8�ƙ�1�!����W!�� ��)�Da㨼i�)�:���%"O�@��M&\��a�H,c�Bm;"OR�P	�<!Ш-��F�
!�p
O:�4	Q˞L��� H��mL���O�+G�Ӄ$YH��F��I���t|�=@���?��xt�	��'r <
����Q�������U9�n�qTeF�BXm�ȓ�Ρ	H�~;� ��[�PtdE�ȓu��E�F�	8 q$��s4z���	��(O��8�+�/.rP��E��y�h(�O��jt�i>��	ߟ(�'�ݰ��Z����Sc��'|\xpQ�'����׏�?.���U��3lk�i�
�'��=��O�/2&iCa�+jRT��'v�d�Iڸ
���6��f�" 	�'��а2*�T@.��L�32��PHH�����	H<��X[.ƣI* R��v��8l��K��?IK>%?��2���b�@"�Zq�����!�Q?V�*��Di5�=���5<R!���8�q���Al!�h�+�
.8!���G�@�SÐ�#X4�7�!�Dݐ9=�Yw
ܡCZl�ْZ��qO<�F~b�Y��?I��ς`�#�
��b]5�_�d��|"����	�7jެ�1*��`����m� e��C�W8��䅞3���؃+[/��C�I0����č�'`���G�;m�bC�I9���S�U"hohY�Ձ�W�B�I�5q
�����f�\R��(T6a@����a�@�}��[�c�"��D;4��B�i�~�2�'a}�AR�*_�D�R��D���B4���y�G���)�O}��w�O��yB)�97%L�2
��E�%r����yr�N�>�t�s�F7;x��Uϒ�p<)��	=܌�A��M�F�z8�s %@2��Z��#<�'�?����$^4V	�eJ��DU#�H����F�!�dȻd�TM0���8V�:�0T!�D�G2l�`#��'F��1G�iO!��.P�0(��0@����s@!�	����	Nx�Ɛ���R*�E���?���$¶"�& Xׂ��6d�`*"}BA�L'r�'$ɧ�'^-��j&*
�|�h� LWEy��ȓODP(��ݢ%���l�,���7��yIg�H�"��S ��4Wu,�ȓC���8��[�(�# .\�ȓ<*��%���;T ��r�֓.:���=A��I1W��DK$S�hq����7Fx�{��0ZӴ��	S���"|�'ɸ�`��:a4�X���C
�A��'0dl �!ZB;>���*�`y�
�'� PåG����
oE<�	�'6�5{Qo�!#T%	�L�/1�,��'d���"�`��5�Ć䳢�~�'�����i��y^$������K�P�GA[E�L�	៸��I�\�2���I�$�u�%�T�#*VC�;?*��{C�[u��cj�L�C�	�o7�=af׾c�H��b �/ �C�I"�r$d�#^� � ��ś<����$No�'t&L����O� А�`Ќ{���+�'{B�ي�4�"�d�O��#�����5!e�|$)��bЂ9��Gd�����El�� F'�)^	�@��-l�e�1�8ErL�e�-����
�� ģ͔a�(�=_��ȓe"%(À��uI���A�&Ѐ̤Ol�Dz�����9����1��~�D�v����R����şp'���
HR���l�tl����r4�tB�"O���%�V<"\Y� ��B����"O� 0��&F����a/�5|$t�"O�Uqcg	/S��qU�[�hnD��"O\0+S/�&(�q�o�M^H����PY�'��ɋ�7m.ly�l��j��]��$Qc�ds��'��'��Y�t�W���q����!�zԩWb<D�Ԙ�mB�nҔ�.�EnJ��7%:D��� 
��C&��S�U�F�R�3D����Ҿeꄡ����2�4�iS� 7����<WԨe�?X�Q����'�'G�Rٶ��3�������yub�qT�'�"�'oƔ��ط/ �0�s��*� ��'�n��pG�4�"���0u�(���'B�,ȵO�sG���$C��s�<E��'�αK"�JY�Ҩ��K)r���(ǓT�Q�,�ӬW;M\k� ӯi��f��@�'gE���d�O��2�2W�@��� LN�g h �O&W�Ȥ���OD����Z�g≥U�N�)���72z5e�N�yGF�"��P
P���	P�'4�ф�)�3��^��+E擹f�n,["5*�p��I|~�$(�?�'�HO �� ٨V.H�7DE=\�h�U"Oޱ�C�G�ZU£��f�� ���>Qs�i>U�	d}���2n��+�k���K7	^4j��ᢟ�8�	�P&��O%f�!v�6��Ҏ��l���+��V� �rk
�p���'��T{�
��?f�%R��[1A}��y�
[(c���  Y�G{f�b��'����D�l*�	Jce�#�b��aD��?Q��hO�b�x�C��Z����G�)��c�"D��Цo�$# �ɗ$B�e��!`�"�	��M+���d16�lx�O웦��h�����_
	�H�C�铧 �����<����?1�O�~��d�ϣm��US��� 4x4Q��O
v�ؤ���jW̉c�=,O�� C<�b��A� ���9���4��r&�hWo蒥a),O��� �'��\�(�e�X��Yh��H�R�%��H؞��-]���)sCG^t��� $��;���A�����������䌛nnu��Xy�T�X��i�'�?�J~b�4S��<�5͐6
��aJ�X.�0�'���+ �J���w�p���-�O��K�Te�[�Q�d�ѷX�B��U�3�ēGނ!`�Tt:X�!Dƨ�(�:�(�R!7O�8�TꐺD|l�;$�xB��!�?)���h�X6m�-G$��.�g��8���QC!�d�vNr�� �ʏF"Ĺ�7Ŗ'�xR�<ʓSi^��R��5|���QV�R.!��}���u����Ob��S���D�'�R�'��I���%Q�L�Ę������B(��&�H�!��L�g�I�O�R1ۄc�W��X�v㖲y��$��.Q }Vt�3�|i���xr��o�t��O�#.�(hEn��N�\�$/?i����SS�'y\m� `:}���dށU�ؤ��'v��R��/KP�T���;a��XQM�,R��4�L��>��%S ~��:��Պ&S���gh
'{� ��n�:���Od�ĵ<a��?��OP�x�Gl
Wv"�S�lM�!(Ta҂뛚M�
 !�w�`k��'�԰q!�
?7���5CӊoJQId��#�vp��mR�	���'�pؘ�A�f�� V��<r�2
���?����hO�c�8"L�W�đ���[�>�*�p�?D�XY`��&��X��{�V��qO
@nşL�'�l�C �~��4-Xᑀ��=�z��N�/)V@�"�'��	��(���|rq�A0)� Ib��Ú"��$��B�ʃ�T4�^�q@���way��4\[�=Ѐ�V�GE,��3c}Q����+�,���ܑ	���$]�5q��'!�	�m@�d��l�*e� ��¤Zs�t�p��I�]���#h�3V2ൂF3�HC�	��Zܺ�I<G�ԅ���3���V���ܖ'����[ir�����M��@-.�舘�D���)@G\�z�b�'���)�j�/u}*���4�r�-�@����C_�Z�$����˥O�r�!��
戟��z�k޷i��ӱ����TŞx����?9��h�x7-Qd����Ÿ]��%�1�с3G!�dC(��XC��
1�b8	Ta�+D�x��6ʓp�Nl�_*bn�C	I6:�!��?A	�&�$�  @�?3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  8  �  )  )  4  ?  �I  U  W`  �j  �q  ~z  ��  ��  P�  ��  �  &�  ��  �  ��  �  j�  ��  �  I�  ��  ��  �  ��  ��  ��  � � � � '# �) n+  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�
��.B*�Z1�f��+%��O���$+$�T�J6)M3i�j�+�R!�dI(�$-��G�!P�Ȁ��ѻ*�!����UaƏ�R�2@1�O܅M�!򄕑[>J�!2��+��Dk�N��t�!���-<��A��@�uy�q�A�4�!��wI���E�9��%�k��!�,���A�k�^��Q��$#�S�OT�A���Af�Q���3�ր�
�'ؘ	Xa� �2]t��O�*�Qi
�'�\�9����,����6�D>y9
�'��a KI�}?�!��K��{%�ł	�'�P���]�fDD$P&K tsX��������>�࢓!&\0 J��]�:F��A"O���D�%5��xZGKC�& �lP�"O��c�p�bd�SK8sI���"O�a��HabV�+�'O�}]�a�a"OT��fj*6���l�EB�LK�"O�в�,1	��0�&L1y>�y "O6p�bE�jE��C'�b&��B"O�6� 6m�>�*�Ř�&vP�3"O��p�C*R�TJP@�P�LM�1"O��C1�T y�4��-��X��"O
�jQ�	�1����#��0g*���4|O� ��v��C��af����`�R�"O�Xk���f�Q���X��< �"O��a�Y`&���!O+v���"O��``J8.D����� š"OҐkqOL�y��O3yҬ�8�R�L�o�n1��C�<4½ÖdWv�yD}��M	�i��h�����a�*(�DB�I�<���G�7Zʣ��@�"=ɉ�T?Q�-Z��|�)���!F́P�=D�@�'J� rl�Zg�RUZ��4�p<����v���� O�[1c!��fn�0$��&>-���	Qx��/C�Pnp�R�BP��y��Jo�$���E< bQY�R��~���ӟ��>���۱ ��V�_�nhK�Ig�<Qm��	j�X���ߺM���R3��xy"�i?�⟢|z�!p��烑S� Ӳ�X�<���{�&��'F�f�J���J��=q`�DHJ[tOǵt����LI���hO�'y��Mh�F�X��|�`�G=q�	��|�&���5^�,�
d�I!�������s����`�)�z�PTG���
�R�d�}h<)Ħ�d<�ؘ��Ss���o�o�,G{�k�:���f�S���(��ˍ�yRH�Z;�1���O�x	�����y"A͇Y�(�1׮��t�>e��8�y¬J�;�[4��~�*��֟�yr�ϲb��#�\'o��A�b8�Py�M�^<�a'V�H�����-b�<9SI�6���ش�[(���X`��b�<�v�R�A6PP�7�$^�4͐�`�I�<�7�7'3|\� j�j�ج�ѯN�<A�*�f�42B��Z�� E�I�<��d�#L��@�É5�t��B�{�<y�l����C��T�0���"@�v�<��!ٽx������;a�$��tfJ�<ya��������6N�&��e�E�<��
|L��)�샴���
fA�<�GDޠU�>52��X2{��тvk�R�<p��.[��@U�,C�ɢ��XO�<�
�)��m{O�V�`J��Ee�<)5��$��` 4f��&���r��G`�<I�DŴ^%Z�㧖�i�d�Ä�]�<AQ��O[�qre`W<n=D%R�(�p�<a4D�x���V��A��Q��FC�<�@J<(�Rł.�𢴣�c�<�1�Ð�ZDa���:!	 �zgjYU�<����`/��%l¹!�0ZrC�X�<9�EH�K.����`D�"sz�Q��Y�<9
ԃ,�4���%��3k�(H7��S�<�⩉�4F-��T�`���+!�E�<�'�.v~�I���K�)X����ƈz�<I�e�l�����g�
��P��w�<G���f7�t13��t�rXZ�`z�<!�	02���HU�<
��!���x�<���H��a'H�F���9w.�n�<���RC�M�E�a��!�Ke�<i�/V�R@��@�ßP��A5f�W�<qg!]�On�qɅ˗ca|h�n�<)Q�H
�@q�v��͐7*g�<Q`�)iub�;.-��!�m�<q�&qP�!pC��*є��j�<��	R�|�������8�fEx �^�<�n	T}�+��n��R��W�<�2kT�fZ@�V���6eR�T\�<� �A�f�#y�E��K���p��"O�pA ��T��Eӣ*DG�ԉ*2"O�h��4X�a"+�38�li"O�2��Z�b��4���5"���"OVMK%cޭM�t��b�ͬ�����'n��'O"�'���'���'�"�'`�|A"ʓ0H`��c1j�x���6�'���'���'���' R�'���'�D<��GٛY
F%H�HVW�4�2"�'@2�'�R�'�R�'<��'���'Nx�� �����Y��ӛ$[rظU�'��'���'�'�B�'Q��'��ԫ�i��
6�Ɩ4D��Q��?���?����?1���?���?9���?a�F�k�����
��(oܕ�M_��?����?���?���?9���?I���?���l/p	xa��;I�C��.�?��?����?����?����?i���?�)�+C��!GX
+��lj���)�?i���?���?���?���?����?� F
.K�t�9Q
65�T��M�?I��?����?I��?���?���?9C�D'P5U��'�*Ϡ���E��?����?y��?��?a��?����?��*��@��}�ǧX�*g�Țí���?����?q��?����?1���?����?���B�X�ka[6�
�;�D�?q��?���?����?���?i��?�LL�p8)XF��9��@���?���?����?i���?��\8���'"i�� v��`S.��2����h����?�,O1���>�MB��_S��Ô�W$]��y�H@�<�-O�qn�x�U�����x�3�A;;���A5�C.p�ah� �����3��nZl~B?�V���m���!	֦�� ��(]�g�J�{'1O*��<�����2w�E��� _���"��#<�<��'��I㟈��6��y���l�ܭS��E9T���Q� /Mz��'��D�>�|�e����M3�'T����t=����D;�򽹟'���_ꟴc��i>U�ɘOX�|�N�%�>Б�'�:.�r�GyR�|��1��ܟt�s��3����́�UT0�T� ���џ����<I�O
��"�
9ZRr��e�t��֙���	#:"9�,4��:,���[1G�K�ĥKE#��hcٱ��~y�^���)��<!��G ���×F��~L<��6�yt�"�>�/OD\���w��iK��6Ѷ̨��	�o�L*�'��'��L� ��V��ϧ���-ɾ4�zq9�E3��q��F�u�t�'�x�����'���'O��'��H��@SԈ��)�*V��tr4\��ѪOv��?�J~��I��a�,aCh�HS���j���؟$�?�|z@gK��,:�c��&NR�h�/�*T�fIP�έ���K�L)���:�L�OD��ƅ�R�V56�Z���W'�N���	��d�O<���H#��D�u�_k~�a)��O n�[�$��	ߟ\��ǟ�9H[�L2�X�ւ$F��������v-oZT~"J��p�'�䧲�/�NݙrT�sX�1���&/`q���?�Uh9$#����fZ��X�Q���?Q��?�Y����p$����+֚	��9��U3]ZH��4�IK�Iß��i>��D�]ǦI�u'.*Tsя?{rVI�IB23�4�R��'�x�&��'��O�H��ɱx�ne㕌8C��ٺ"�	:��D�Oh��O�˧voD9�GP�VY��""5�t��'���?i���S�T���"����۷Nc���B�Z�5���*b��6$�j�<�'�@��X�I�Q�]�叒a2Q�1�	@��B�	��M�V��# h=Q�@$*��9���_�<���?� �i��O�<�'��NƆ���RU�l$�L���*���' �K�i��	�ip��HUҟ��u������5�F��L:Z��1���$,|O ��%2Hn��s�j���9U%�l}2�'p��'��l�mzީ)�A�aJ�K*�
#s�q�������Iq�)�S�N�"Em��<�Q��{��� v��Ds*��+�<���h�&��u�	uyb]�@H��̇`9>� �*Ka��Ͱ��<O\��'�'��d��4�	�td ��c\1��O��'M��'f�'�� 	R��@�u���Q�f���.?	b�V�u#�݊�4&��O�D���?1fHZ�hӼ<���6k�zL�4bʆ�?���?����?����O ۧ�Ԑ]�D%�U�C��a�O$��'R�'֖7�2�i��%�فz��D�1 ۀ��S��d��I��,����`s����p�b�?��A'
����&��Yo�th���z�IKy�O��'��'�2
x����2��	a�T� A�-������O����O����YQ�n����Ӱ^�,���!P�1�'b�'�ɧ�O��������\�& kQ�	�9�|��Ћ��v!�V�����,B�n��d7�D�<1��B�S��t����grȬ"����?i��?����?�'��P}R�'��!Z2�1&�6=��ڥ�ESC�'��7-6�	���D�O���O
L�&C��Z�`���$W�d3�����L10}v7�3?����.R��|:�{�? ���jӽu��y�"(�$��15O4���O���OR��O��?a���D��saٶL2�$�ǟ������K�O0ʓY#���|2�U�h޲�Bp�P/]-P�����+��'��T�e�ߦ�'X}�F�	X�h��I�;h�����Z#h����j��'��i��'IR�'g��)sf͓7��)�gE�(>���'L�Z�<�O����O��d�|*����"��T�S�l(��I��f�{�I��?�O[�Qsl��Z"4p��I��2����0'$���CC@�i>����'|$$���F:6��� Qi:D�� �ٟD�I�l���b>��'G�6-N7 O������H��T��Jĺx,��O��D ֦��?!RU���I�O���:&
*O�R�ʕ��9-2��	쟴9�o���'�����Sbr-O��h�nE�v��
؀|�����'��I�L��ǟ����l�IB�EѮ��� uF��M�(B���0Z`t등?���?�J~���l���w�晊�lF�5� ƹp;���'O�O1���ؖ)i�J�	�v1䔳�f�@����B��xC�:O�������?T*&�$�<����?�©E�&��!fb['\��������?���?y���d�L}��'���'@��sfa��5t��%�����DT^}b�'l��|b��p��H��_�|���q������ݿJ�F�k� |Ә�&?�P��O��$ѣR�ʐb��4Ա��#,����O��$�O��D2ڧ�?��	�"�,l�"��7<<J���B��?��[���	ş���4���yG�0P%�T�T(J�O�paBGE<�yR�'R�'*��KV�i��i�	��?)uf�>T���0�Jy���a�� N.�'{��˟����(���x�I�n/�M��Ǉ�72��k�aF�Q��'������O^�?���9 ���$g�M�@�����O��b>��mB�q+!3���6f�>$ e����`y��Ud$��
\��'b�	5)�\I�qI�)LS�0��>w�A�	؟D�	�8�i>M�'����?i���o�*��g�Ƙzf�}�eL���?�ĺi��O���'���'���<Q��\��2�(���D�'Rp8ǸiK�I�I�Dqb�Oq����X�*-�3-��Z8@�Z��"���O2��On��O��$=��%OL��2����Z,�v��8��Q���(�����Ĳ<"�i:�'����@�;o`���#J�J�Asך|��'��O�}ôi#�ɪk��(zP� +S��(���Lm�x��LV'��L�gy�O(��'�"`ŒQ�l�R/�y���r�Y"r�'������O��D�O\ʧR�A�.ǽ>��v�/��'if��?����S�T�̂;��U8�"E�����Q�*e�ʔ��*� o_������~�|��0q0�2E�¡;&1����-��'S��'����Q�jش��C(��
�`#c�S9�<��?��?��čL}��'=��n?�2�y�o�<&�����'�B�� ���������?g���<I�	�Lt����sN� y0@�<�,O���O����Ob��OTʧ]�����t��ܸ�B�K���Q�[���I��t��l�s�@k����q�	�%
r�1��l� ̣֠�0�?Y�����ʹy��?O���H*`�x)K�G��8Ͷu4O���W�2�?��L2�Ķ<����?��E�=�\������imnQ�SGF�?��?Y����D�y}�X��	9�APm�PMpT( 	$��?R� ��ߟ\$��#��G�T��Fr�8���-?� ��z��ɔ���'r �����?y`�ݺi<�铰��H'h���K�'�?q���?i��?���)�Ol���cC�=�ijw��'?2���F�O^t�'5�	<�MS��w�2h��KQ=S�N���דz(ٚ'���':��).�期���!��JE�M�F7n0P�B�2z��+�F2p-xX$�����D�'_b�'���')Z�$�>���X��w ��1Q� �O���?����I�����$f���������?1����Ş= �i�Ȝ��  ���^
q`���Ab����'�*�Q�.���a�|�^�$�\�-�ܐ������Jj���?���?Y��|�-O8��'
�βa�
M�t&�E�\`�"��q���,*�O����O��d�)4F������T�<ݨ���'n:r@��o�(�g���cj-ʧ���,�d��A3�G���fI�<����?����?���?���$��4q��YB�I�a!�49R*� a���'����>ͧ�?15�i�'��t#G�/cj���.U60�����|��'��O."�i��	�6��]�iD	)41�Ǩ�=���� q���8�d�<!���?)��?1�%ˣU�c�E�Y5j(9�+���?�����Ēc}��'P��'��3�^��IM*���9,H�"���3Y�I��0��Z�)����-6���	ceöS�����T:������M;�O�	�/�~��|�m�'zj�0ipm�b���]�e�r�'�r�'����Q��[޴:� �H"o�:Zv��K�%k<A�����E�?��[���I�D��u��Չ'q�ҥ�C���I��D)㦉�'�0�@��I�?���� �!9C��$G���r�]|xFM�S?O�ʓ�?���?	��?I�����g�h7� � ��@���}�'��'�����'�6=�rl�N�jcL���-b��y�#�Od��%��)�bm�6-`�H�Qh�3;��ǉ�~� q;%�j��1�@=p�BPw�I}y�O���	`B���F_�Nb������'�"�'B�'C�ɀ����O��D�O~��E���IBoY&^�Z����7��:��D�O��$9��Z�a�`u *�&� �t, ��^R5+�! Fx&?�BE�'F\�I,V�����f�k��qaK[�s�X���ߟT��ԟ�	i�O��]�OP�=i�C�Ke��ɶ�]"�>���?�"�ia�O��B5K�+�о4�}��k��'��'��'Qc���4��AׁB����Xrct��s�*LHA�� n;.�O&��?����?����?����Ε�]|!5.�pe��/Fy↲>����?����䧌?���7��@!vH�*�o>6�	�p�I[�)�Ӝ)WI�l�<AR|���+#&Ybdޝ$�~�WF$�"D�O���O>�*O��fg|=Z�ӗO�M�B��OF�$�O����O�i�<9�U�@�Ƀ)q�H(���4��r5f�9�5���M3����>����� O�>�H�ρ/7��sKU�ĉ�Ԫuӄ�58�`��3J~��;�E"s,������V�z=:��o���	��L�I�$��՟$���e &́@S�Qk�|� �]��?1��?q7[�P�'.�7�<�D!Z����$%RZ4��I�'&��O��D�O�I�7#�7�-?�B���^�;�ሥ^U��*k���i���'�D�'���'���'_�pCA֫<��D�G�ƹNk꼹��'=�[�h)�O~��O0��|��ÚL�r�ZsjԷGp�M"�[@~�B�>!���?�L>�O.�i0�ʂA�Nm���GJ�T��"�#@����T���4�� 	��-��O���ƒ�VH�͐fmT-P-B(Ј�O^���O���O1��˓{t���P>&�VH��-A^P$ze���<A*O�Mm�j��D^��ӟTQq�ɊZ�	QЯ�9q�hKmy��Z'xқV�����O��� Ey��[q��y��
X�5	|�p����y�X� �	�� �	�h��ğ4�O��\:�d�F�k7%^)�zARc��S}"�'��'���y��s���+�"4���>#9Rq�͖;B�n�$�Ot�O1��� 
p�R�I�F��p� .,�$�gf�G$�I7Xp�*��'lv�%�������'c�\��
�x&JH�C,_��h�S�'��'��X�<èO���O����;$ց	6#Z9LEȥ��3[G⟤	�O��$�O��OX}��F�K��Ġ�C"y�z�����l�A$G�'c:)J��&��>'f"�F��G-A��c�� @fٲ�&��<�	�p����dG��w���̶t�	�u�W6�tK �'��ꓑ?���/��4�L�DꐐqheɃ	�@4���q0O���<�vJ���M��O���E#����DjBxQ����R [�^dۓ�r��OTʓ�?	��?	���?���?�ֱ�ĥ�eMҬ��)��R����*O���'���'����'Ǡ�H��+F@j��I9L\>0X��>1���?�J>�|�BJ/��ɘ[�w����/��I�����C~��_�K�����>2�'���6���BC��2{I(Tv�ѝȤ������ǟ�i>͗'.�듇?��_�N����tk�1�$��
3�?�F�i��O,%�'�"S�hR��J&E�IL<��,���#~�6�n�O~�`��&��0��$�O��cA�D�ac���&�h����	�y��'f��'&�'��	O?b��ڱeg=ة�vd�:u��d�O~��F}�W���ش��!��Ts�g� C��P�P|[�8J>Q��?ͧ8�(��4��$H=��tcBޒ$Mpb��Q�Ufґ����?�$'�d�<ͧ�?����?��i��/�\9S��W,|(J5��H�)�?����ĝo}"�'�2�'��S��<kn�m5&�C���0��$��	ߟ���q�)���?@�B��4
�A�6}�����A�.�Mc�O�)҇�~��|��L]�e���9�T�P��"�'���'_��t]�hs޴x ��HCnR�>��%eLt�l�Γ�?I��x_����T}�'�P�`��oc���-	�2�	u�'�B��Ƒ�֝�ow������	�u(9o��r��h2�a\�$>�ry��'i��'���'�RS>���I8.Z�aD���?����Q�����O����OP�?�������V;�\#�l�,���"�M�?����S�'*���۴�y��̃�:l��IB��U�ժC�yb�æu��������O���RT�V��S��R�  `��K6�j���O����O��g��	П��	��P���f�|�Y�ܪb��l��}�����៤�Ij�	7q)����IW $�
�UON�r�AH^��]'���L~�E�O����<bޡ��'̡D�2$�ナo������?Y��?����h���$�Dh���T���i$mZ @����$�S}�'rbiӈ���I��9�#��Z���"�(ߨ�p�	ß8����e!�1�'�Ȅ��ʀv� ��T�O�W*�q �T�P���0	,���<�'�?A���?q���?1R�֚΄͠�fF[��y���DV}�'w�'�Ou�����ȝ��N���XqW�W�5-���?I����S�'Z�\qD��s����b,ř	GRq�hN��M{�O$9ĭ_ �~r�|�_���pdӊ'����N��<"Θ1��ܟ8��̟H��՟�S^y2"�>)�w�XQ2Ќɫ/��<`��^�A��0K��%�����As}��'�'䄰'M2F�>y`���T� e�t,�f2���\�t���9"Q>q�%K�B�)G� ��y���N�H���	����	���������G�'���.�&��U8r��o������?9�>��i>��	�M�K>��#ʸ�.M���P��S���䓐?Q��|��II��Mc�O�n�8��95�V�T�Z|Җ� 9p\�l��A�Oz� O>�(O��d�O����Od�r�L�F�BF�ߏvd�yX�&�OV���<��R������	x��)��4�4<�Q���:�$|�A ���d|}Z�M����S�D�M��5{% �v�r��ʎu�@��Th$X)�����#���=��V<� ��޾��lHQB��R���O��$�O���ɫ<1T�i�� nܛ/�"�����^�*�'��ɖ�MS����>��{\�!S�F��A�f�߬NK�����?y2���M{�O����"�>��O?m;����{Ep�)mN3y��`a��'�"�'�R�'e��'��ӑ-��B��3%�%BrL��at�Y�O����O���)���OX8oz���k��\E7O:�ĀJtL�P��D�)擙	n�l��<��"N!�y��A��z{�1	���<�"�'S��$����$�O��d�
9G���D�k�~u`U�'K���$�O��d�O|���	����ޟ���BH9t�\es�J�,D���0CjJ��:k�Iџ���n�I�z�$Ec�m�%{����#kK3�K���S��E(��|�,�O<����?�p����I�R$�3)�<|.%��?!���?��h���Q����#�I��0Q��e�Շ�O�p�'_剻�M{��w
�y�N�d�>@)�ݤk_���'K�'��� !W@�6���Bw�d+������h�X$̞� MƘ��'�����$�'~�'t��'�V��A+� >�
y�5FO(B�d8p[���O����Op��6��@�^�2A	�#fv'�	�.�ic�Ox�$�OL�O1�F����_5}�d����(\�*}:�J!*�j7m�~yB�Ӊ@A�������$.|���d��kuD�!ܖ���OL���OF�4�˓��Iޟ��$	�(	D\1B�
-� �@�!���4��'���?���?A1㏘)�d�Ǐ;C�u+EA<2��ش���5$�x���O��O.�DkU� ���f�ѱF��,�yB�'��'���'��I�8J�����C�:�k<R�r�d�Oh���]}�OI�}�X�O�XI���`��!�h��/�d��)�d�O��4�>���q�b�"V�|�D��.�ޱh*�S����g$S�L�v������4����O��9["D�c�-W�Hp��B����O˓S,��֟$���|�O�8�x�[i����"_ dtZ�O���'�b��?9ѧ��$VD;��>� w�}<h��E��D����$�Rџ��|b@FQ��C3�y:�R@bQ))>����O8�$�O0��)�<�!�i[�}�%MT�'����j��Z�ZA�'���'�|6�3�ɪ��d�O�LH����\I1ϛ�a�Y�˶<���V��M��O>И`HJ�2& �<��$C�?����;t,�z�l�<�+O����O"���O�D�O�˧; ���-�Y|�CQ-�$Њ�2S����ʟ��	_�'3ݛ�w��`QO���16j)Ex�m�E�'p�O1���{�ja� �
=rh|"���\�� ��:!���'��tٵ�'���&�p�'���'w0�����4,�� �K�4u�-���'�"�'��U����OT�$�O���
XnYc���h�&�P��O�,������O.���O"�OJ�i�_9.�R��jA&P��۔���Z�&T�rt�#�B[��ss��ɟ�w΅�*�5��@��وXg*��'���'�S����d,�=�z5��Ѓ����p\ɟ|X�Oʓ7��V�4��e	Qn�� 0PT*������<OV��O����(�F7-;?�����;�j�iE9[*`K�"�ci�p
�-�1U��M>)O���O����O��O�3�#�<q�����*�����<�6T�(��ߟ��	{�ߟ�� .
�?kؕ
	���@������O���,��i(TF�Sѥ.�`�;�Q�4�1GMn���DA<��4���p%�T�'�r���] ?���ڋVq�my��'p2�'+�����V�h �Op���"cwЙ�G��o��P�j�9#�d���?)gZ� ��ԟp�I @|h�H7�ͯ��aZ¥� `�V%��E�'���`PA��?�is��4�w�Vq	��9�2u�N5���!�'�B�'���'��'��~8) �7zv��p#`�h��qk�<A�w,�)*5�i��'#�8�I3QZ�ig�C�.�
M��yb�'N�	%7V<lZt~"�
>߀ �C`�K$`ÎԔ[��-`RiA.�?�d+�ġ<����?����?	S+�$���0լ�<? ��3�@�?q����N}��'�"�''哱T<�A�ɖg�н �[����$��I����I[�)
�f[-ٖ��0�.Y�\��3)�1l�rC�#C�����Vǟ8#4�|Bd�&B����፻?	А� Y4&_��'��'3��Q��Y�4):�:1�X�+)8ȁ'oԳC1����?���^��F�d�|}"�'/�d�ˇ�^�萢�7.l�)��'�r��O�&����A�׭9q��i�f�X�|�Q��[,��d1O�˓�?����?Q���?�����ا#W@�����7?	03�C]�u���'��'�Ҝ���'�p6=�2��`%�H��d�P�F��Q(�OB�D!��IM^�6-w��(q"׮>>P���,�4A�(p��� U�z�I�Q�	Jy�O~bJ�/�Tq�$hJ�T��A1F��B�'��'d�I9��D�O��D�O����3Ŝ����K �&�,��3���O\��5�dT����"L�4
�M���ù*��	< 9����s_�c>���'U�i�	B�}��C56A�����X[���	͟���Ɵ$��Y�OHRL
=ͰQ�
"J�1eʗ\���>�(O}m�Ӽ붂;J٘A�ʍ�]-���'��<���?��]�xP)�4���Wn�H���'�Fh�%�� d�踶�*Hj��dO$���<�'�?��?���?��eˍh�X%I���F��놻��Cz}�S�h�IK��/"X��sК� �i��8��R���	韸$�b>��W��r���R���j�K�@ԅJղ�nZq~�.�	Q(Y������$C>N�	�p�[�F1���2g��?K
��O����O>�4��˓?��Iǟ����+0�z1ZF͉ou��c�g��k�4��'����?Y)O��[�f^>���hխU�~Ota�Y��耹i���.,�!Q��Oy��&?��*^I��5"�7<�f����2����	۟,��������O�(!ٗl^�qJpI�$�*
L����'��'%���|b���6�|B
�9c�(�C
W�L�bl(�C��v��'�����Ԭ���V���B���k�.T�gٯ_G%	R#I�=}�)���O|�O��|���?��?>�=
A�T�5���QtBZaĊ���?!*O
E�'=����O�*�ÎO ̆��͛!����O9�'�2�'�ɧ���k�uA�9RX�]0Q�O�@�Lm0$-ǒN^ܙsE���S
%�B��|���Bt�D�2����"����	����ǟ��)�SNy��g�llC7n�-���ѡ�ék�V�p�1O|�$�O��n�h����՟�F)�)G�P�+��uT��BL�ȟ������l�P~B�Q-T�H����$�z9��3$J3O��|��h����<I���?���?y���?�/������� =j�u��Gr.�ծA}�'2��'��O1�}��.�:a��% �?E��V���o�B���OēO1�Ę3�D{���	�jHu��65���Ù�v`�	�;�8[��O.�O���?���G��$DLݟ8���a�@��jB9���?i���?)O.��'�"�'���	�F<�;R�:|@�9�A(]��O:�'�R�$�)�Z��w柧V4R*�"Q�g���?O�hhRF통Z�6�&?IB�'�6��ɉr7�ybM�y�L|��I�@�����������O�O$"F�IN������X0@쒢sirG�>����?!q�i�O�NT�Gd<�A�J	����E*\����Odʓ|$VȻ�4��d�*d]H���'Edd�d��*;�~��Fυ%\r�*�i/��<����?���?����?�f.�	s��-��)�5J&"(Q�Q���DUk}��'���'��O�rh��,����\�H������>�l듿?1���Ş1�a3&D�\�t��㏪'*\�� �Q6cV��/O���s���?	Q7�D�<�boܡE]���GY�e��5�Uπ��?����?���?�'��D�{}��'k��*�h�^ݻ�B��8����'�h6M7�������O�ʓ��y�,ǣ^�lU"k�2_��5�Ԏ̥�M��O~-��,B����>�	��`a�"-�%SoĐ /g�D��2O`���O����O���O��?�y�Ï(lJxc�/�O}6%�!'Eݟ��I��x�O�i�O0�lZA�	R�PP�A$�0 �6�����*%����̟�ӧn�I~҄�((��Ę�lHHp�n�9D�t��@�IFy�Of�'H".^,_�xs���@�H�M�'��'��:��D�O���O�˧3Y4��1+T�s!rPW*�3q})�'�X��?9���S�ďU7��j�i��:�f�A{��!Q�
F.N�F���O�iW�?��2�_!�e�:/^�z�+h�2��O��$�O~��i�<	ķiD�u���6x:dAB��h�<Q��'��	��M���B�>!��Th��j�}hr����.#K�|J*O`���b��*�z�������r(O�
�/�k���C�'�5��h�9On��?���?���?q���מG�~%�A�
ܸh5�_	e-�'����&?��	.�M�;0ذ-4�ǸoF��3�%S�����?�N>�|��%�M˞�� �����-�f��0葵�&tr�3O�p��?iQH"���<ͧ�?eB��qD���@��"Y���פ�
�?A��?�����$]}��'�R�'Q��PB�O8@t�c�&�d�IA���o}B�'��O\�Y��W���&�5�f�jb��4�EO@�FH�Q+�D�Y�S�GM�D�˟P��"+\��,�=C��V�M����O����O���1ڧ�?�w�J�>�0�\2ܭ�G�����������<饴iL�O��0f��h`�X�rq�e��W�*O��OH���O(
Dm���gP���#Ꟍ-��C�$p��@GS�/`�q���䓬�4����O&���O.�䌘&������}_N�#t��	 N��sg�Iiy��'��OG⡘�,�Z�bN��.P�1��'��!X���?����ŞV�0r�~�ء�钗x�&%�gƃ"g�@�'�Jb�Ɵ�П|"_�@hდ4I����M�Q���r�'NΟD��՟�����SyRh�>���'q��r�����T��owF<q�"���D }��'���'���Q&�B*��k�/ǖu]<5�Ξ`��摟p��lF���'��@�8�2�&�"Fd��)R.	����Ǖ;=sj\�����?�zU2���BL$Isr$�(Z!�Z#*U �� ��Ő1+�<�2K�	A�L-�CE�$��a��0��~�$̢<#N�0aT*�(�#�7 ���H�aW/n�.�@�HŠ�::�����Q"+6EB񈖏^B�C�L� @ƕ#�%N3%b�C�Й�ԁ%m_�j��D�b�4~�X-�q�GB��HW+K91Z��vח�Dt��oZ	Y�h,R��>j|(X��۞:q`�%��6-���'�B�'0Bʥ>Q.Ob�䰟 `C�$%���I���	WonE�"��c�%�`�I۟X�I�w`iP����>�xy����9�ߴ�?�����d�O6���O��Ok,Q�&�$��6ђZ�bU�ӡ�'O��Ec���	^y��'s2�'y�'�l��$�Q5��P�[�Z�@�nZEy��'��'5�'��'N6�A�U7�P�C�T�DArț ��12��'q��'���4ן(}���S�M^� �4i�0:!��×�i���'B�|��'�l��D\9'*������YU��`'N��Y��	������*L|�-�l�d�
yP�	 1K+qސ�9���)1n�qm�ݟ(&����ݟ|�u�TS���I�ƙfZ�t���&g�5mɟ�ISy"�'��ꧤ?���?yR�C,z���T��$X�كs�S�NK�'H�'����'��'��	R"X>Tg� K="ȓg�Y)B�[�����P�I���ɟp��5�@�:o���B�L��pX�Ƀ��M[��?��@�����O��c@ F+���cl�4,o�I�ش�?���?����?Y���D�O��DBz��A�5Ō��Lh(lw֜��?E�D�'!X���Ã�Z���b���*Dl���M{�:�d�O���O,d�'��I۟��{�TX!��N6�Q7��(��qnK�I�lb��L|Z���?���V�[��+r  � �G=eR����i�B�'�����OV�Ok��"U ��C�Ѻ3<�:wnۧ8i�I- $��$�h�	�����y�� %x<yc���$~1l*�C�7ě&h�>�/O��$4���O��d�8s �t��X�T|pA#�4U�<��� �$�O����O쒟1̧<��`��N'ڈD�Db�a�˓�?�I>���?�A�B��~��ܴx�`�$6U#�&R��d�Or�$�O��&>�騟���Q�5%lm�q�Z�Y�@pp��1�8�m�͟�'�t��͟�z�o�Iܓ'�^�z�� 7��  R�S7G�2mm��4��Vy��'GV�>�d�Ok� _G�%�C/[�pqsW��.S�'���ן@��T�s���
F�zP��9�Jb��{Ml6m�<��f��&Ŧ~"��?!ᛟ��G�Z{ry�3��):l�*C�f����?���76�OP��M����8,e�4�oM'Zܬ���G�˦���)�M���?��?qҔx��*�)��9jX�i֝^��L`$�i���'Z|ʟ�I1H��5��N���*I�lȑߴ�?�*O��d�<�O��*h����Pv����[��h��cP��O���~����~r���h�����(8$�#�C��M���?Y+OFU�Oi�O�5����m��V���B&?�d�'�4 r�3�	����'��d
7rczġu��"\@�#�I�V^���	ޟ��?���~Ri�v�m��$�(w~���R���M� �\��?Y)OD˓���
1A�xiFw?HJw�ك�M���?���'!�	<MU�6��?�����֨�T��\.�')RR���'�ş�A �U�q9�cƨ�9��m��B���Mc�"�'��	�FfO��{0O	~
�T	��W/7��=9��i?"\���'������9��$�@���<�`E;�k.��O���<��Fx��u�өC�
(i�ޏ%��Ad�V��M3-Oz���mڮ�����ON��p�_�v6d<�[�|C��GXh�f�'7��'��	-�9OR��i@4΀�N�6Z�T	~r��7$�>A���?!��?����?�3�#T�v�x`���\�k��*���D��b>���T����ЂY-g�J<�a%�O�x�A�4�?����?A��Ik�����'���#� n�J3(��\���O>��!h��iD��'!�� ��9OD���O��� �F�9@������ *��5m蟰�	&���|j��?�-OD��!C΁C$����ݰe θ9Nͦ��'��T�,�����ISyZc"R��do�������3��\i�"e�.a�'��	ӟ�'�b�'MR͎6;�Ց�c��_DLk�k �z�\0�'1���<��ß��'�"Ih>��
�$9d4  5|w�HD�z�D˓�?!+OF��O��$F�#��$�o���0�M����ȵ�G6C���n��X�	��8�I_y�O-^ꧺ?�1"8�q� ��B��W�XSAbxnZߟ��'��'|���y�\��y���#DFm�&�ܳ�Ƙx�ʘ�M+��?q.O���Q�d�''��'Ǝp�D�^�"���Y�eV&�LL�5j�>a��?!��HJ �����/G�,i@���$QeH�VjK��M,OT����	� ���@�O�N���t�B�?8��m�L?���'s�� �y��~���OY�-�t�O�|���+)NL���4�?ib�i}B�'&"�'�J���d�q��)���M�bH>���J�Qt�lڋv=P�ǟ�'��z�䖲l���1F��#��hX�A3G��l�����Пh�������<����~b ;�f=�ᮏ6x��d�чE����<	wER~�O�b�'��s��� �̷.�ܥ Ɛ4V.<7M�OV�DF{}bR�(�IHyr�5F��*D{�{q�]�Z�^u�VBH��ď�/��D�<����?�����S�/���xE����H�2�]&7��V}�Y���	Sy��'b��'��4�c�U�0�bc  ��|��ю�yBU���џ��J�8���@5玔B<�1f�!J՞q� �i�����'�B�'���]����A���J^k"Q�i{�����	֟�K|��V?5���P"�|)�N]3��)�"�7f�ă�4�?q+O���O~�Z�L��|�Q`ȣpV}B0�̪T|�2tB�^�f�'8bS��I����O���O�MP��	�s�~ڥMg�U�R����Ov���OD�3Ol�'�?��O��P��oΞ�c�G�^��;ܴ���O��n������Ɵ��ɀ����2��ƾ#�d0��O?1�P��i�b�'����'R�]��}�qcƕz^��GSЋ���6M�O��lZ�`��ퟨ�ɡ���<Yp�3`�D���E�`��ʆ���Q,�)��yR�'���p���?هk�h���&�R��Wh�y�6�'�2�'��L�>�-O��D�� ���B��A	�Y�2��+�>*Op�ǚ���ޟ���埸�s�+E�R`cF�I�h�e�Mk��?�6S�\�'�b\�X�i��!�FŢ5˺a��)�
����>Q�.�W~"�'U��'��P�֝�4�����B�bj�0�w.	?"�~6m�S}"V���	Zy2�'�b�'@ E�Q���%+���׍�}
@� �j6�y��'��'���'/�i>��OA��CqD[�PJ&���*�R�z-Rٴ��$�ON��?!��?��o}��D�7�0��t�v�@�J��Mc���?���?�)O��C�D�5�g��f����PB�t�h%��� �M{�����O���O���5O�'S2���D�VH���D+!�ڴ�?9����$�O,��O��'��Ά�gl��y��9b��]��ɫa\�ꓘ?)���?�$(d~rZ�|��>+xؒ>M��Ty�D4��mZOy��'J�7��Ol�$�OV�Dt}Zw��	�ԉ��F�l\�e�ٴ�?������'r�Ix�'VB���N�KL� ��ܝ=�x�0���Ц-����H�	����O�˓L/
1;�O�
T�\��3�ȼ¸l3�ie���'vrS������)���$Q�Q@ŋ6.�$��i���'��'����O*�I*3h5	�/��Xɜ����Ƿ��c��D�+�	����I�L�UJ2/~��N��'�( � ���MK��?q�T�X�'��_�\�i��i��!w�,U�ǅ�^�2I�c�>9@c�p~��'@Zf��'��i݅����=��4*T��;*�B�By�D��'.�	ӟĔ'/��'M�6]�:�	\ QBq���6���(�O���O
�$�O6��|�B<��H���Y��V��:M��R���ɦ��'=�\���	ϟ��	Tx ��g�H���@���N�X7,W�#�P�O��OP���G��5����O����/JTx��kR8j�������e�INy2�'��'��q�'p��O��I�̌=,�խ�&�!��iO��'���'8�y�����O���O2<S3������T�ѩp�v�)b�ͦ9�IHy��'	����O �X��s��=��]�9�씪��<i�$*��i��	��PS�4�?���?a�i�i݉��脵d��
�Ε�0��]B�i����O
�0�2Oj9��y��I�8r8�\�pͅf�z(�����=֛��'��7��O��D�Oz���u}"W�p�a���X�q1��?gt��&���M�Wύ�<����"������U�J�en]���Q5����Á$�M��?)��?Q��x�'���O��9�+U�.T�1��úvx`��iD�')�H�!6��Ob�D�O���Չ�>�(+P �@����S)����Iڟ$Z�}��'�ɧ5�oTSa���#�ܨ/VP�AF�C����Y�1OH���Oj�$-�dg��j��÷*&b(ъ��M�d�$�O�Oj��O0�� py�u@5F�@��!�O�}���XG@�<Y,O��$�OF�D1�i��|"A���+�D�K2��$+��Q/�E}r�'N|b�'O�i� �ybA&@��]�2H�L؉�d�'�,��?���?Qg��Dj!�)ؿ��ũ�"j:���W1O��$l�Ο�'�"�':ҍԎ���>!6�_�$�3�Z�^kP���ɦ��I̟X�'�rA)�)�O4��]EZ���S�И�rש5_��$���I�Ċ ��x&�D��ESL��D��54�`���^�Z	o�iyR�'�f6m�p���'U&?9�%*4J�cwƕJ�-�ĠT���	�d���W㟘&���}���׿Tl��1t��?�0���G���I�M���?����?�7�x��'��¢�	����1Ǉ(*�ac�s�.�0a�O�O>�I%'Ƕ, ���6�+�ȟ�2}��J�4�?����?��#��'���'W�dӒ7D��ANĹ?+���̇
k�֖|B��yʟ��D�OP��_�J��O|�@xrb�5N>-m��|�	���'>��|Zc �=��
�&bJ�$�?j�t責O�0@fN�O�˓�?���?�O?�Ha��&P�Z���� �hav��#	r����>������?���u�N�h��W�O���ٓ̀v�v`���?�,O��D�O��$3�I��|r  ]1F�� n9xm����B���'�������Y�㟰�j�R@�(q'G�?q0h�k�����O���ON$>��K|RPʖ7)Y�T�E֯M�^ �თ�6�'�';"�'̼@��d�F�,�c�U�O���ySɂ�ab���'O�Y���I��'�?���#��&jn	����# p��i�Y쓽��O(�֝�C�!��0oLm�)*�@��񄘓U�XIk�E҃j���rюcЉ9���|d\�H+	 �0pPp���|��X��8+�r�Wn�9I���)�W�Ow�8�a��z��s$i��HM$��5�.�"PK�l�3]��h��P���9�!d�A���� 6�����)$*Y��)ʚ"xP! �فP�Da1!��]���9a�M�E�ւ=��S����oϬ	r�|���̇7��Dإ-6��|��eʊg;�����J�G�J\blȢJ�ܘv�ɍ#�z<�P�_� 6�YxfϷH0��V�q8�g+jx��4�?���?A/O&���O���!	�"�J�qӃ��]�4���O����, �˰mⶇ�w8��k椃( ��!�p:�yڡɃ#'L��7@a�|��
߆k����	*�`����Q*T�D��Ĥ�BlP�I$F���Ot�=�)O��jg��K�lE����.i�X��R"Oj�������Q����<�+MI@���)�<i2��-Z~���H�v۠��a�ƍ�>e�4JT�c��'C�^���I�̧g��)kv�%�J���A�=~�P��$ �$��0���ir�@����i�Ӈ@�ZR�3������9`"��gD�S�* �ϓ�������i'��IB.Ş1.���l�q�'�џ�1����w��qԢC;��)��3D�h� '>("t"�� ��P��q���Op�G��3P���	H�$��n?���T��}�X�z&۲�y��'�r�'q�*�-��~@@t�Fo�F}*���!�9o��5 ��xcƤړ�I>
=�)�"-� �4�)��t�5����7H�v��M;%ɚ��(O�%� �'��IS0X�(C׏�py���3 "f�$/�OV���G�+�b��!gީ="yk��'�O�h�u��.��4Z0EG�_��E ?O^%@��NC}r�'g�O*��'0�EB8�o_	/��p��p ���ƫ1�:��$DV}*��c>�����s�X4[��H�z�#��M�N�VeBD���6���X�"~��!�t5�BGA&b�X�xWM�"M{ܼ)�O�����	G~J~BI>��5�Z0�T Q�І�a�<i�d��j�4�QGϐ�\;t����Q[�'kH#=�O�<�TCY2�^��8"2�@B�O8�D��O�p�nZ4�I՟(�'��'?h�b9�`�-��X� ���'��	tÞ�[����1Ov$�F@��[˚#w��9��D��O`�E���S(LL!�8�4��-^-|��C`P�a�pd��,������O���%ړ��� L\�9�)/t ĺ�aG�!�,f�L��)˼T��Q����@�~=Ezʟ�ʓ[��i�5�a�U�"�蠳m�)�>�qW�'���'��IƟ|���D��d��9D^��ܴP�`d�F�Kd�ܡ��]� H`|���NR^Ȩ�O�(�v=J�+ r�1 �%�{-���r��+$�H���ý��'=t9�3&X�,�l�`Aj 4�b�w����<�����2�ӧ(L�{��Р[@�X�l x�C�I5xt޵�C&ٌ/T�J���=� ��঍B�4�򄈦,��n���It��B�VFm� !E*Hz��9�ş-�y�'��'LreC��'1O�&a�=�$Γ�WcЕ�'C�(Ӏ�<�����O�9�A
z�l[��UjP	��䕱"��dLȐ��hi��a��)��"O� ��;��^�o|(t�I�����'�F�O�W�ؤq��)�$�K<G�@Pz�'"���֏��$�Ot�����O*�d�4tE��P�!R������GO�Q���$�ʧ���?!��$0F�8�.ȴ�bI!r�1r�� C�ɧ����;1݊�J@ע_�6�iYhԼ��'d��'����OH�+e�W%;~�d`���>F0�H�9OX��+�O�E�ՀW��H8�h�b��j��ɯ�HO�S��Ѫ/�ҝ�u�p�
��I��$!�M�9�M����?�������O��0$�>p��ᚠm���h%��J���Q9���3׋*lO�T�p�_�)�M�#$�w�%Z'�O��1�� ���D�,��,Д�A�h��uH�M}f�L�Mi���O��ԟ�ϟ �'p�����Q���Oü;� �'�Bt����*5N
��HH�]�Ṉ"�;�S�T��O�VT�P�E�u��ܫ� ��KC!�$��]��y���Q�nq` oUo�!�Ĕ Y�2�a 	�7:E�wn^�&�!�A��Urۓ���]3�p��F]�<�G�^=��0G/8(�"`\�<�f�Xò	���7!�pc�f@�<Yt�`�5�QD�7Gȭ;0TP�<���.J��cg,^���D�G�<�M��)���F�=
r�tk�B�l�<�2�Kz��L��j�~���'M�}�<�Q��(0����B�?	�����u�<�L�$=�&�St`��wJt�p`�Zy�<I�e��Kt�I$␗[=X�(uCM�<1C`X�B�0i��
�"�P0G�_�<��`��C\�d�C��v����v�<���37�����O�'��5Q��J�<Y�c��ܡ&�SUvLQ�I�H�<AFK��2L�7'��?�DU;��j�<)�#
	:cL��(��`��B�<� �<BZp��,��]@�J}�<9�.&	��ib� RI�H����{�<��(F
��(���@{"E@a�y�<!��X�8��q�C"�^iz#ŀv�<�̝ 8��(�buc�Dz��L�<�0O"p�v���K�"[�0%j��[E�<��'_�EB�xAꎪ�칱�g�E�<9ʋj�pv*ՠ��=y�k|�<a6�@g�4X׫ GJmz��x�<a�;d�2tآ�ٙI�$Y�&��M�<9t�����k��Z�m�8�9"���<�2nFC8Hȃ����N�� �e�<���`�썚�c�t���ۦ�Of�<1�g_�G�04"�"W�{G�6�"T�H����"yBy��iM�.�Aj'&D�@� ˈQrHM���8a�Q��"D�t2k �qr�ݛ$�zBi� �?D�����bD���AK1W���"D����"S)@��Jqa�}�@d҆m?D�����Eh�ܝ� M�8@*`�>D���f�v��9�O3f�0��@�&D�P�G��)5��S�K߶5�Pe�D*D��ir�c���1�5Zph���'D���⦊2h�M�B�\#JmV�Ke+D�Ȫq�ɗ.�v`ñMY�3�2x�2�)D���D��*ЀK`�U��$�`��'D�`� �>M ���"*U���$D��s ���əd`I�V5�dB8D�d��͗�L��M$J��LU:@A9D�4Y�㛩ed2�!&,��O~rd�$}�L�Ȓ]�S�'0'`ax�jT�hN y �$��r+݅ȓZTD�g��X	D04h�l��=Y��2v��� ��H�EK�n��e ��xK�aj�
Oj���#����GH/���񫜖oȞ�q
�'�©�"c4"�J	�B.J>��Ǔaؘ�j�`*扐o"22�4Iޞ0a1�� c�xC�	�3���a���8϶��f�$�nO�Mۗ(�|�S�'R�D勱��3(�5���;-�,��C�,2#e�m]R�	�m�TU�ȓ,��Ҁ�V|p��%U$j�Q���B=	!���7�!J���Y��I�� �fkХ{5P�� zn�U#�'�A`���@��@PD��c�T���'S(�0�ذ �bt� �ڿ?�ݓ�']��зD֗	'��s�n�+��<J�'{��A�:MG<��H�F
tQ�'���� ��qL�i����'I�����'���!�ǀ-;���
ŢڔK-ؕ��'��H���[���"EJ>���'�p '�x^�u"" ]
Ut����'7E��(N�O��UZ�-ƺI`�l��'�0� 6��5	�Ļ�����)h�'�\�	�<���20�$� ��'�Z�*B�E�BikT��6z�~<�M>i����j�6��@��$m�A2�� �!��D���C��Qclx3P�H6��O�;��'���b"x�� aaCU�4 �'RR ����|H�+�hF�{�cu�xh!�d%6�}� �)צq`����DyZw��Sf��
�@!�����!4WHx��D7�nm`��2�y�]c�)C��W�Y �:Ui�99�D3�c�Do~��AH?E��'���:�R!�(d�জ.�9K�'Q��C���e�Z�C��A,vW��I�'��AR�� -�`s���0<�ʏ!��Vmzi�4�Uk��h�C��}$Jp[��@�wSt��fX�*���ɒ��dy3M'�Hæ�L�/6<���,�υ͞&�O�X�XT�%��Iy��|���&a1�`�b)��6���CL*Upu��"O��ذ�E���10B���H[B�]�McJ��u/�>C�T0�h��e��n��C'�:�@!�60$��xi��􍓶Xp4qB�n�7?jp��+�_8h��O`eF}���J<�?�a���S�
�T��S"f����^QX�b%���o&D�p�퓝b����Ζ?c�H��v�� ��+סP9hl�1�$�O��q��9  �P�hҽE��dc��|�`M�ea��=M~�@/�?%>�[�'Ԉ\H�z�L�|�^-��O-D�ܣ��·O!dU��AA�E�$�QBF�Zk�}�JF��X�O���H򧌜�<��]Q�
�4Y���RH<ahY��jG@�	��)�d�S<d�D�6� e����V<�A�闗(��Z��M�S�N�J3�M=L}^�Q�2<ON�H7�]�^�S���Oة�Fٚ^�"	˴��[�d3a�.Đ��a&�Px�14�A�9`x����&Ii�Aꖧ$���	��@蒯�0�e���/���|r�2/1.�E�Г:��ѫ���D�<	�B�' ��[R��� 3SV�0��]sJ��e5Z1˥�P}��d���y�U���Z�
j��@�����yr$Вn��Z���  $)	Q��-��$�l,(%AY�2�n�9`Y(䑞��\0J@���K�0M����+\O��q	\�<;b��V��/0U�$O1v��/B�a��q�Q-  ra3�>�O�`���S	CV}���'�,�Z ��K-�r�-N>�$[�-G\��ԟ�u����vY6A�&S�9�d� �A�?�pC���(�z�HADզ.s��;�9q��X���G�T�Tl�6��C\`�C���,O�����W�׿[ᄥ�G��/F�~�Sa�<q��ѩ+�j-j�EH
,���� 7��lZ��˓h���5�yZm�&�]�L���#O�J��o��Qޤ	�i-�O\��"eX��U�&�!#�!)%D�.=�X�X�Dͫ*9�6���$�̓�Խ��+,����9ǧ�0�@4 gP�Fx�*�4�w�_�q�`�['�*�M�矤Ia��u��	�K@<eN�y�\�T&L�S��'���g*�O�μ��f�* Qp� �O�:&rA���܋��� *�M�g���� R�ZƤZQ�9�!d�>�j0�"Od�����:4be�G�o���HVMF�y�0BT�SC�i>�	�j}!�T��y��@�O?��EҲYo܄@���x��P��:�r��D�k�>����t8@����0iq�4�@'��g�$I�<�l:몴�nN�=�L�O���f>?yF)�
4��T+��̾�~rțKb�%�"��>2�TM[�O��� �Ll���'(3,O��;Q� Z3���$��Qeհ]�0D)OH���W��f͂�A����.O��؁)b�U��g �8��%�j]'V�xu�<������%)��:lg�T�$��m���*��"n�����]��]�BA)?Q��ܹ��GO�pqd=�̸q�g���f��Fj^t� L�eY�̺1��sqO��̹s�o�r�hѬN�x��H8��4��'���� J�E�G_9� X7`��
��O�h���9>�U�&ݶ#h@P���x�!\�-�Ё�'8��c0�z݅��
j��}�RmU0q�����U����Q�'��c(�(^4�ԣ�@8�D1�w� ����5;�;�I������V��
 �!8J�ط�[;��a:�n=�韔8 �-\�k�IA�Q/�����	�/a"]�4����袓� $~<�4��E�M]2��^B��׀K�Wy6t� Mםc�R���?;�V�J�F4��O����h ��O��i�IS�@R��JD'�D����=%'��#�&��;�N��N��B�����(�⟄���5 �t�ɱ62h��5CJ(!�.qY�]7��>�e�#^���{#D��H9n\B���$��8�1��w�$��Ǔ_�.#^3����L�[��=SaXo����YF�h%�"zN�g�
*.^����$U�hY�qF k�Pp�F��֏@�?�L�ZpBº(��ib��C��0<�b�ǢS��D��G;]��l�C�����Y�S���ߖ�z�N:VZ1�'̤<��$�7���ւɦ@��+��ĝ�P�3���B��0J�;(̙q��3x^ *�@)c̨5�ʍ;CP�=y�¦x�xH�	D�f�8)���7p,m�Ç�+a}�P�w.�R�݃�8A#q�F�%
�����o����$ϲHB̨PA�J��� � �*��խx�� y��B��nU)�R%!t�*�E��<5������#e.���IlzL�E�G<(q���8s6݀��*�I%jX��`�\n1OX���`�Xf�,���R�PФ�'�fQ���ঙɄ+�c�BԱRH������>���jT#>9�d�.8Q���I�xmt��N��T����x��WN�Y`��S�E\a�܍�iݵ��o7�U�R fFـ1�@ !���K^��&���'ސ�Pa%�a�gy�@	7�Ay��Wk-BT! �O��~��C=������9zZ�-A�E�"m@�uaB�H�`X�1#uT.6���vf9�S�\i ���&	�x�Ж`��pm#?I�O0g�4�?�2���\� ��D�5o����4��YP���H�tX��A��>�[��r�,�2N��PѠ��S�L��'��p����f�S�OB$���V�>�;����.�����4�0��$K§>'�z�#<O�]�7�E-G4��e�P�FN�1 �x�ց��>�O�H��s��%�VH��'Z��D�R2��v�l����-1�Ь�4�I�H��Z��]��52bdϜ��d_%B�Ι���#��4b�A�pџ�8c"SD�O*\��M�.�Ll�]���U��'�� �i�)]k�d0�ޒ�0��'+.
橐'+\؋DHQ~e(P��'�R�26�`X䫞+pOdu��'��BS��"`�)ಅЄnr���'����Fԓp��U!�C �i��<Z�'o���S0{l�E�ma ���'��<���!W��� ��a*�I��'j	���?&oT����X�l5r�'�`�a"JW����@曹Km����'F��:�C�#��y�$#�0<5���'~�æMȅ\'.��3lB&7o��y� ֟/8]x�H�=R�����9�y�N���ܻ���#kΊ`MX��y�++>z=��&��g�X�R�Z��y�L�?[L�H�D��<d�tl��N�yr̀��4��$ˡ��X�����y2mJ�"�X@QM $>��j�lʎ�y2%G�_P�˅��f�P��Ҏ� �y�("{�l:6n�)?�	IN��y�$���2�N$~@����y
� ܌��G9I1C4�U�,��"O��QV�յm@��(C3��	c"O*qQ�2Ȋ�� hN�s|j9�"OA�D�0���H���҆"O��x�۩l^H0¡5k��P�"OX��FB�&|����߂m��t�5"O@��Iτs#�9S��
&	��'k	����	�`�8��U'aT�	�'�F�(�K�VRw+�#�Tu��'�� �*���Ћ�ˀ6!tx��'�*y�K�8M��	f@S��\��'/Z�#�cÁ}̸�p�R���̉�'��ܐ��D&w�"5C��`�=a�'�� w��$Zm2�G�3Q0		�'5��c���3
����A��l��'B��h��N���B,M�P��A
�'� ���
c��1���X���	�')�	�#H�*YA��Y�{����	�'�n�"2��L��R7c�(�0��'�T��%�j.��Uf�t���K�'�xkċ��"�v�"V.��Z
�'������Ў�zgh��6�����'mN�k���?V6����L��"��`��'�����#Ƣc�^lY����H�R�'���h借�Lʜ����J #�p��'���j�j�'�T�(�(U�x3p��'�dI��8|{f��>�H|��'Rn��gOܚz� ��R�5�`��'l��X��ڌމ��W�5��yB�'���2WZ���J�Z�.,[�'�8qÊ� ��� z�I!�`�<�q��R��<�%�*~ ���\�<�a��3.� ��㊋C�yǹu�<)�#���rC�w攑!M�<��J<����eOq��Ã�Iq�<iG�B=]xQ:*Z�p���Մm�<�e��3�,�Cu@ϱ9�<\sBM�d�<U��+a��K�D�za��G1D��37 �9S�0̑�5�D�J�.D�T*��ˣ?:)b�Kʣdp�I��>D���`Y*l���r����\�*>D�88���%AVxP� �ߔ:����&�=D�|�Eʄ4r����dߐ�3�'!D�4@��ND@���cH���^���?D�@@�H )�
�E�/�HxȦ,<D�8I�	H[�$�`��J�$�kUb:D��S�fXC��4�p��4��i5�"D�<"��K�b�1�BI�:o��X�/ D��!��Mx�B3'ۆRr��3$�!D�l��X4>�
Uɓ��*Zz��em:D��O�0;aD�F�D|��Q-.D��bP)�%�L�ZF"�Kƪ�h�(D���B�U�\����_��FS�:D����~�Z�P���ug3D��(a���r���%h�
��QN3D�֠� ���Z��g4+u /D���!S�< �{�)ׯ �V(�. D�4b�nG�K ���@G�L�f)"D����ϙl��B5D�2I�����!D��kDK�C2�t�"�0K���a��?D����@�� ,��.d;��Ԡ>D�p{7%��u���"5G�I�d�=D��QSe�b��Ф�sWz���:D�t�� �w�V�pƄ��v�:��"D�� �����Q��0�"�>5��t�"O���C���L�s �D�*@�$�O&�=E��+~*�#�23a��x��W��y�\�&���P���%���h���(OT����H5��#&iE� ����� ��!�d�%G��e:2'@<lrp���3u!�d&#riRoڿʜ��GB$0\!��>���2`��O�����*i[!�D@�_Ø�kY" .����d0!�DkZ^����0�@�1�E�<#!���q��]�͋9`��p�$M>u	!��8m�����
���#�@��!�D�	��Q�d

�2�f0��a�!��[�,�|��UĊ���)�t@(�!�dͅ_�Z|[�K�a��Y; �Х
�!��
�(������
-����&>�!�d��'�z�(�]e�T� O���!��'��S���.",���aV�/2�C�I@i�s�J�4ev��T�ֳ�6m-� )Ȁ�z"	qa�"^,v�a�4D��3F��h���I
9�V�K�J=D�D(����EHZ\�4}��d'D�r��tA
��7W'�,izJ&D����M�C�q$,�f��9��%D��*��S
��\ �	ʩ
h�����$D��@���U1xM�rg[#6h�ѱ�!��oZ\bԀF��B�t0°j�d�B�ɞ9��})BQ�vn�
��X4?u
B䉚x��_>�� X�m��C�	�;�>�ڦ`G91�I��!Ԫ"<�C�ɜQ��pi� �$s�� J4 R�Xs4B�I82A���[,`W��[E`��gH�C��N�f�K���#�|�x�02�'�F����P�X��އ����'��5�F�]������Yr^���	�'(h����!5ָ�'�F%8�� �b�fA3�k��D�N`;�'��D�ua�3je��h�CB�0�	�'�t0'�r��� ���MHp��	�'��M��F1A���B@C>.P���'hx �O]&1��ͱ������r�'n !��D��@�
肥�'&R�Q�']�|Ch��G1~�z�#�'���Zc�-�ɚ���!o��)��'^< �ïH���ЁiT�w�P܈�'�P�c�d�50oBd���s"	�
�'-*����H0EF(m�� �FQ

�'���eO�8s��`�6o�6��	�'=� ��,E.)(ٰ4�Nn��X	�'��ͩ#��&B2p��m��z�͙�'�\�!�ķ'�:�r"B�zn2Tش�Px� �)h�*=Zv	&�6��'����y�G���%Zc7$֠�k����y��F3:�� C���j�(i����y�5Dn�qTy�r�[fm\�y��J�,0�)R��d�r��`<�y2��d<(�,]�%�<�Ł��y�n�5"� �b�N��v�c�o��yK4"� �N��daq���<�yRD��V��<�rc�(BK �Bc�5�y��g�r�Q��٘O������.�y"�ym�P�E��{����sH�yboE�xqysA()��|sI
��y�j>vF������.Q:"J�;�y
� J1�vl�F������1%^�l�"OR����A�U��L�1R"O��;��z;~�)��Ė+�T)��"OF�ST�ʈqd�Q�.P�hҞ]�e"O�X��	>1�,]��J=mĸ`"P"O�e�DNQ&3JL�*Y�I�jT��"O��WA	!@|���G�1l�r��e"O�1j I^)]��R(��1��q�g"O���o��,�ƹ��ĉ)����"Op}�Gn�*(Dx��`ŭCo��W"O��fFǾp;���&��pQH��"O�����N�t�����J�	8>���"Oia*1n��M(���J��h¤"O�$�bɉ�V�x��jW8ḧzC"O�� ��:1,��Y�C�zXr8�&"O��P�#5Y�� 0Ç�fh�2"O����-W2:89�� jL"Ը "O8�PVk��r�I���A"l-Ј+"Op��@	�<V�갓�F	�v�y"O��@�Cm$��vc�+��I#�"O�P���I���8c@۾`��'nqO�ţ /U�X²U�DH��{+�a�"OJ$BL�}0���eI�"�=��O���	�'X�.�r���>:>(�E�C9C�!��=,�8�0nZ�;Y��AC�'	�!���B#4$f�y��N�iNL�"Ob�
p`=�(��`�y���@"O2i�cl��M�D���(��vRhA�Id�OGB%!D �8����_�~��91�',8\`��G�w��2�m�2le��C�'��x*��8F- |"#�׾d�B���'�8�� �F
:T.T�uEǣ+"�!P��(O תR����QKɯf,�#�"O�U.����5�4�rMC���:�!�<"T��A5�H�ȅ�Q�|�!�dN�5�R� A፯�$�HA[�k\!���x�@Q���M	\f� Ӽj@!�d�	kW<���a����A@\�D,!�D�&���qh�9�	/��X!���+xl�˕�F�
:ҎҺ!�!��Gx��2f �~1J�-G?4�!��8%�\�⤂+o0�Q���P�n�!�S�}D�	Gb9�HM�K��!�Q6UL��;�hA��`�IF�Eh!�$�1��Y��,��ՅΉ�&x�6"Ox9*P
 z�3�䎌V}�Q��"Oа��̜�q�@�QiN�	���"O�
g�U�k�0�mf��ehU"O,T��vT�eJ�*�d�r(a�"O^��D�\�b��=����X��M��"Opi@��I�4$�ے�&twtSV"O���R*N�:4������@q.�!�"O"}z�)S�|�2	�ȸp� (�"O�q���'+Ȳ@
N�:�Y�"O��b#/5p���҈Ѿ60F��S"O!S��B�� �e(1|,@�"O8X�C�A�޵%(�I���"O8�㔮�!D�B-�&G�\�̡�"O|�c�U3C76<����[�4Qb"O��1��OGCh�1�&�&��(�w"O8��um�#m�$���D?X�TKV"Ovh�qc׎~ �U"��L��� "Oљ@�ʪk �2��5�JD��"O`|IpCJ dj����!C���1"O� �� �L;Z��1e�!�☁�"Oz��3�2y�1�Bǟ����"O8����A�����H�/l����"OX�� Jא1�N4���gdtU�6"Ovx��R�@��d�&�)S���"OJ ���9�Ҵ��f�21V��`"O�m
0!��u�� ��D(�	�"O��9���*V�Lb���%&�yu"O�p������R�n��Hr�"OPm1��U{5�A�pM�7c,�RU"O��C �
�!�,U���!e(���"OL��kV����4L�ZF"O��X�\1Ć��M�hs�I��"O�ő�&��?�e���$�3"Ob� ��V
�jŢ�ΰk�!Pr"O�Y���Ӆ^��3H�2P�L R"O���
PF�R�h������"O��c �J2�A�!�9-��+r"O�!�MLm:	�ao˭q����"O����J�q6~�SC.��\%�`0"O�M1W�*}y� rM�	����"On����y��q���߄2 ���"O�|��R5�n�QM�
Iy�Y�"Of]�b��m�&՘PM��q�ʑx�"O��2��;����N�u�5�E"OhPy�hް �mD))����"OT("d(��b�1ɛ�Z�2QS�"O� �r��<�,��)�t�U:�"OjMCVʆ+D����1��SE@�[R"O�Hs��˶*��X�AN6-;vqi�"OJ�"��9J�+��$�d��"O,�s��ē>�$�@��>䉈�"O$�@AO�c"��Zbi�6Nd�g"O6\�6锿_�ѵ�1 (8b�"OP�BG�1�4�Q��߭]�����"O��aH�	�8-��2��ȱ"O��ʴl�'a��� %��
��7"O�9�o�6`Ű����чwMp$�g"O���4i� 3�:�Ic!��xKpH
�"O�0:��F�tDi���Z6�1`"O�c#ه.s��˅M�f'L�;B"OH����|�aB��,km��)W"O<��%n�LM�M߆$^R0�#"O*	x@�٨�Ĩ��L�>y\N� �"O�P�-[�2����]�gW�!kd"O�%M��|�px{��A� j�ՊB"O�E�g��%(�<�"eF>	,nl[�"O��"�N�T��H��i�b��1��"OU��G�1a2����ڬH���P'"O���7+�(I�Xe��t\�9b"Ot,��צ�y�"X�!ǔI1�"Ot��ë��8���;�g��Y�HEI�"O�0R5ˁQ���Cv��7g��	�"O��82
]�mD�` �N����9�"O `�&��P2��RT�D�E`��w"O�\fe_����k�O��/�Z}�"O�\�C�ޘc/�$��+S�V���#b"O���.�p�O%�hIx�"O�H!�LS)TIE�WB
@��q�@"Oҵ�&t�إ�@N~U��"O�����ݻV�����HZ29�\Q*g"O� H�M�00�ǇH� �N�A�"OR$#M��$�1�B;x*�-	�"O*����4^uP���
 K�"O� YH��VqQ@�`�l����"O*�CŧQ�<i�Ub�2�(8y�"OB́�oTTߔ���G��jX
�"Olz�Ē����2g�+�� 1"O>@ �GO/�$s�5B�=�v"O4�w�[�7�ػ�b�E�HH��"O�Æ(�nT��;�a�QJ���"O�����\3 �3�J��34�I "O`H{��L�E��43 T9 �"O�ē!��D�l`2%L��u#�"O�9kG�~&4*�-��(�"S"O�P�C�]_�E��"8�N���"O0�X�	�~����L6O �-�&"Oz��쟞 ^`A*�4[����"O�<�b��p�.ءI� *W0qc�"O��rE(��=d$鲓���Bl�4(E"OX�C�/�B��(1�A�����"O\̻4��% ����� � yzL��"O�,��nV�Xc�[�w�n!�`"OP�ae
��b���P���u�ba�"OFx@���9p�UzR�U�JM.M�"O��)�C����! H4^�h<��"O�ܱ$j�X�^�b!)ޔ�Q8�"OРP)��/V�� ��_���"O��ʣ$��TMp$C�\��4"O�dZ��N0'��h�i�9b��"O��Хd�<w�L�#�T�X��;�"O� SG�ػ(6h�#�@Q|��"O,��A	άVH�$+3��0FN�-��"Ot�K���A�4���I<\5*t�"O��SFI	N�P�ǩմ$'
3"OxQ��	�#5Ь{���� �K�"Ob%DOњT��E�0p��l��"O�ԄJ�!������5�n)�"O� ��	>�� �V�=	(�%��"O��A�UBz��'$�Ql9�r"OB���6>-��ɗ�ڨj7"O
!�TĤL�J�A��!�d|�"O"��i�=���>��p��"O�11KA0V��a�OZ�7�xe��"O�T���)�D�"�M=��,�"Or�᳃H~�P֍��k�
�J�"O�-�Re�Z�T<kЌ�>��]7"OJDk�;4`j	xd,� Kt��"O"�;�7CY�|�P��<v���"O>��e��o{�HX�Z�T/x��D"O�`�"M�"����T@[+H \�3�"O�$�1)˗y�s��շF㨠yA"O]�ahL�Ѩ���.ćU�Ь%"O*y+7�_�	����P8��) "O��Є0�N��Eh�U�����"O��c����3��J�f�-V*�00"O,̢����4��,y�σ9ɀ�"O�A���F�2�ع��EԔI߀��t"O�h�K�]���N��Hbj�"O
hȱME�F9�%��`P��@�"O�`ՒM��]Y����V�ܕ��"O���Ehĭ:�����A'2�ȡ�"O�e5�	�`��<�v �n�h�bW"Ot<5"��q^h�	��H���ɓ"Ozy���=��E�2(H�.���f"O�	���h���ض&P�U	V�"O�$�2OZ8	���F
<L��"OX��&a��Th�����U�5� ��"O� �d!��-��a��ܑ�T��r"O�ʠ��oK֑��Ę��8D"O� ��Hک<|���L ���6"O��+2@'+*!;5K�`�6IK�"Old2 �w"P�s���>llɂw"Ob��͗7����7i�`/H��R"O�X��7|�JyB�匞l8��g"O|1��LF�d���z�Z�M�d� "O��`7h�=DkZ!�O�O���s�"O��Y6���|���"%�z��lʥ"O�U ���Y�~���D�##�hQs1"Oa"���Q��\��
^EA�"O$M��l!����� �ru��"O���'���]fN�����l��["O������ ��$�'�ު;Y��YU"Oh`�@�X$v��DАFO�OE�S""O�Q�qb�8o��z�EY�U(��0"OZ��A�Z�,*E�BF	��"O�L���U�*����㐍`�NM�"ObX��c��~,p��~bL�"O����.5i�,I���AV��A�"O����H��.� )�A�A PLYq"O����N����G�rk��!r�|��'�ԩ�r�Y	��I
#��#&�N1��'�z0� Q�{8"" �7����'H,��mS�rBvAz�'��,��-B�!�4O�63��	�'��t��m��=}F�@�R>�]�'D�XC֡E�)���g�ݗB+0��'P�z��O�:i��f�ˊ4@(���'� <
��͚F`R9{W�\�%��U������5Ax��c�=�Z���Cv�!�W�~������L�4���
�!�Ē�i<�l!�J�"I��pG�B�!��[�>�I�6�7>~a�V'S0�џ�D�ԁ�9��		��ȡx���)6�y�\+*�<�&������W��+�y�2�*P�a�OwU8'����yr��d�B�	cb	�Đ[v/�y�٠K�P F@��U[�mӥY5�yr�����[DgA�N�&��R �$�yr%=r �|SA��;N	,���T�yŧ�V����oڙئY7��xb��v�t)cN�s����u�F
ZV!�d������P/�z	.�*M�'�ў�>��Ɗ�1"$� �֟4o�e�%�#D���&+Ԗ,0�b�-.h�Bq�"D�(�"CїE�(�C R."g�T1��!D��Vfܭ_��lp*�"n
��$�>D��3 �:#�|�SJK�|���s�9ړ�0|����+�� �&`�p�7�o�<���C$`4�d�!mz�:���� m�<YrL,,�1��r^f ���h�<�T���l��Lu��Xc�� O�<1FiO�^<a��\6��%bI�<Q���("���1�A	K��#cI�<I��H�{�2 It�V
	S�aB��@�'=�	Z�Oe���T�)B��e�P�o��T9��x�iG��D����-�Ȍ:W̞���x��X�=��������y��r�
��p�!��X1!�f|XaaY-1��s�(Ɲ1�!�DR�R��*�M�G�����:!�߶@�t�y@�8`*"쒐늑c:!��|�MB�� ��YB��Ζ(+�'���5�)� j�S��Of��8�	ч1����6"Oz@çm�9+P�qF��HE�2�'���	}Q�h�2���\�sn�<B�8C�I�+Z���[X���"e�	�C�I9L����d}7PH��`)<+C��?F��!�f�-��l��V�B��,(ҰI�����,4i�0I��B�ɤh}<p�ԧٟ�9
���}��C�	�~������J��g�Q-r�v�HG{J?�K�CW2�,�e�+T!� �C˷<��_`��#��]�~�L$#6�JI��ȓy��sT���tE��_1|�p�ȓ)@��)���P�v��ti�*�ZɆȓ/l%9�KT(,`����h<p��	���d̓m��dY����Ro6|�sA��bN�����	���O<�b��>��ȓ$��Bd�%p����6�Μ
RE�ȓWў0���G]=��icb5-ά��j�n(���30�$�)�b���W��0�D�e�Zq�C!Q/��݇�NR���&j¥~�B	�e�Tf
���7�����	Q��8YE$XiG u��i�p;���U��IX�I�	bI�݇ȓ��Y	U��3~�|��Gib\�?I�Z��0se��7H�b��׿,O:��ȓ��B��́LF�Z�D:;�>���#� �IMV�gR��2󋙲%�rq�ȓ�b�
#�\�b쑐h�?~0E�?y�Y�dŘe�5�^�9Qi&h����	�<��NF{(���BX^A�%�Cl�<Y�1K�J�,ߗC����TaL��<��~��j��~�?��q�q�Ņ#�b���*�yRL[S��]!�$e��C�3�y��c��B�.�8n怼�ă�y��/>*�L �A`� A�b�F��y�πj�: �3U,RX� R���%�?Q/Op�O?Q��H_U2H��e
.6Hiw�h�<9���M�����N�x�c�b�<�ABP )G,��	�%�b�P�jCu�<Q��? t�Ҳ@�9j�X���Bs�<�����(��&��=JwAům�<�cI%o��[U� ��0���ZOy��)ʧh�T��Gꅤ^�0����)!@xɄ�Ix�'��y�S��): ��+4�Y�,ٸ(O��=E���!q��xJT'�6 
}�G"D�h���z��4.K>'iH�hB�5D�H`GLT`IҗJ	�*&HAs�5D�̓ᧉ�g;�9�a(����)��2D�d25A��Y����Do�8�9ʰ<y���ӯu}���
j�F(�1�֔F�.C�	#F�Z�saL�b"��+��N�C�ɷF�I"$
T8���.�'��B�f-�qR���&_�8��v�.�xB䉉GƦ)�%GDx,�1���TB䉍s6�2�(��ww,m�e�E�R=B�I�İ f���0|�vl�r�@C�ɢS�D,��#�>hy�:C�B�I&+�����@� Y����旐n\⟈�I[��~�4L�b�c�����ѭ'2Ѕ�*���QaJ��Lq��2�*]����ȓ.'\̨c�?NΌ�6Û1�|�ȓy��� w�V����$�01y��ȓf�~t��Yn���&��R,���Ɠ>Ќ��v��U����ȮU{����� ��I1�ͅ7s4%�'d��D5HW�	|�'���	��a�)�nI�Z�#ۈx�'*a|b��%�J �Mߢ���B�_��y"N�����;�&�� ̛�ْ�yr��*��T����.0�� CD"�y�&U:�ȱ�&�*-� �a��_��yB��5�����B��#0�&�y"�.��JcB��"�Ǖ#�y""�9*��$�0�f|s�a@?�y��N�>�Y3�ވ!:v�z�ꖂ�yr��������: W�U;�k���y%�/��-�ņ�-e��;4��y$yf��pk�I���hE���O�㟢|�N�j�l����Z�l�XiIE�<���U��(�[�.b�@F�B�<!�M 2�޽A�!��(��k�z�<A�Ŋ8{"d���=a$�(ÊJu�<��i2�C�ܻb��b��U�<� �/% pr�Ahzd�"P|�'?}00N).����t	(~�x���=D�LPp͋�d"b�SL��|�p|���-D��s�A׼3��Pf��VD���*��0|�Q��6��U�T�K����TkQN�<�'��(a�u҅ ��v��`'�Eb�<Iu&��2��@�!Y!�$���M�`�<YA�P�zX(%��)`�}е��Y����<���3NTUs���5A��Saf�S�<Q��,C�>1 l�Yl���e�<���O�+%H���? ����'Dߟ$��	n~bC\�4��ID'�r=J<Y�*�>�y"W<Q���k�>!+�)К�yB��'($�Kp�Xu�"��i�4�y���N\�̴֣r�Z!��QG�<9��W]8�ݲDB�[ZH���Wy��'h
�R��5B���ۢ��5&�M�
�'�^y�R��>!��I�I�K���
�'�f����MH�cG�Ld�X��'���:�IE�Er��ã!�Q4p��'���z��ɺ/�֡����)�~1A�'��0n�)wS��pԎWf�x��'k�8�H	
*h�Sϙ�Vy��[N>y�����O.���eۀW�M"g��w?� �'�tU�-ԃh��2S7��@���8�� �S�5�T����V��y�h��^1��O"�=�}ZTB�+[�xH��_�mb�&]D�<����-*�8�/<_6�Q��[�<Qw��N �E9��2F�k�k
ş�G{��I��k(C�Ḅw����h�v$ʓ�?	���߶������ʼ��㘿2�!򄋝����؝��iQ���{B�$G�����УNV{r�F��3�!�DZ�i��`�H�"U�A�NO��!��Y�2�x�`���sP Q��:�!��?#��`���N��̋�b�!�W0Ly���B׶��RK�O�!�ЋQ�d�y��%�\=C�/�
+�!���c��`�l��2���;�U�W�!�Ęr6�Ia�"������f�]&u�!�$�6�|���`7��D�g���'�����.^A�Ǉ[�C�ֹ��'�Q���" _��`���B h��'&f����ޟp�%Y!&�/���M>9���i�4_,,(u��A7v�xen��O�!򤖓�z�I��$8T��B�!�� ��Ha��%[B�9�XG2��"O���Fۏo��T����7;��if"O�Bt��	�`8��_OV�
R"O^x�sk�?H���Q 2B��p"OV-�Ca�G�>�!�i�#AC�8��Z����}�S�Of�}�W���LU�D�a\�K0�I��'����̐�U��l'ѥG�����'?�Tq����3o�A�D�c���'��ĸkY��Qs���4@��'�`u!�D�oFx�҂��FR�m��'�Ti�S��2��1(�#�?�)�'f���'R4A6���������'���B�T�85����u^н*�'��X��D0)�*��$l��' �J5�=+�hXq$��q5����'��k'�Г��ѵ 't����'qp��w`�j�#�g!e�|�+�'��y#�!�z* ��ۈ[T�("�'Jt ��9
��'�+��QB�"Or�#��zg����L7�\�5"Oґ��Ƥi+�q˱�<7v���"O����
a���D�O�Ҍ.�yrM�ր�:�GU���\�%^2�y�*�TQ�����c6t�F��?�y�a�{\(���8Zl��p�Ί��D%�O.iK�`�(�"=x�JxP1�S����I�,e�vH�V+y�D��-LB䉊y4�ѥHڿ,������� �4�=	
çK�l��n� 9\ɹc�I<]4�ĕ'ua~������r���*$@�mK��y�ļ0�-�s��Bi^v��,s�'�N\1ā�)x �`�
ͅf40yK���'!<��`�aXp��LUp��:
�'��ch�	hV%pl;��x	�'%Jh�q�+)��8b��X�Z�8	�'V�:���&3�U	ECzA�j��y�-Ү^�
��`F\*9��%��y�'։H��*PX4,��4{�)D��y�k�#Y(�u����U�4��� ��y"�(!Ib-��P4=����'É��y��V��f{K�5S�]��bC�yҦ��Q
�牾A%N]���D-�O�@�"Զx�Eᅎ�6;�T�A�"O`*f��y�@B4��v�lS�"O(�06EZ(W�~Q��_�@j��A�"O�)� �5�@�
6C۠S�P��"O�XV� �p�P�p���&,��9��"O��
��ɨW!�4�A�U(c*H�d"O(���H��T��,Y��D�F:�AG�'�ў"~zj��?:�E���O a\}�׃�����0>I��I+
��xW�Ĥ/P�uK��XA�<��Ê�R̢!�� [�Q�^{�f_U�<�ů�5HU���� �V���"�c Q�<�&M�J�ְ3囋�L�2�M�<�D�4�dE1v
tp�EBV�Do�<��G�4e��ik��W���)AF[d���hO�'�n��i �?zJ�i��œ���"O(Ab0O�D�����d��a1ڽ�U"OL�Qɓ�R���ew.Z�ٖ"O���"힆RʌJ7�S�> 2�%�S���9���gi�.�� ��!v�!�, @^\��a��G���񀍮M;!�[5p��C'�]�'�V���OùzB!�'&t���TSo��)�и!!�� �|�b�K(5�Q��/XW��xҔ"O�I8ӯ�AҐ�ⴎ�6Z���"O��X5�^�;��q�%�+57�eJ�"O䄫��.PWN���.t%Dq"O��jD&�"�&R��$�"O��H���Y�HYW�ץ5:|Ò�'V��2=��`Sv)6W �	k�	��H�$B�I�D�ɠ#Jf��Ί+S�B�	�!���s���h҂$�B�V�r��C�ɿm�:Y̍ ޘ�c��Q� Lʣ?1���V2Y�%!$BY��4��0Ŋ�`�!��9��I�F,�m��JVC]�]!��͠4��HHsO1P]�|���J��	^��The��<t�q*J5�����'#D�0�嚉͒�`e��"HT�Qrj!D�y�dX�`��DHDf��*�+'�=D�0��◸)P0����61H�iG*?D��7eF&C{�@�:i���"D�0ر�^��3���//��D�#D�,��صJ�J𤤆�]%����"!�d$�O �0�%@������&Hc�d>LOF�#w��J��y(f�2i�N��"OR�f�����*D���"O(���jP��NP�.��k&�� �S�	K�����㝏���r�2C!�dێ`�6,�B�Q\�r��Ĩ��0!�$� �p���D>z(h�Ʃ�/j!� &\���E数Cg���Ǌ.d!��YF���は��do��C�gL�P!�֊�$�f���eq�E&%G!�DF�,�k��B �I;V�:wFb�	o�'��@äU�j�>�����(l���
�'��4+��)[����fJW�#�jD�ʓ$��=�	W�+���#U�Q�	�'�ў�|bCjG��: �K<Il��@v�D�<ywn�b�J�K�%N4r�|�%��H�<y$W�H,���{z(�-yGB�	�UOj�`�}:��Q�H�e��?I����.�΄rx^�8�Q��!�d��^$E�+؜k�ś�AL��!�D��uO�,��&/�5g���[�!�d�*�1@Zl.�A�v����O2@H�j�U�ZD ���%j�l͹"O����ǔwC؈���/�N�"O<e��-C�=������3r���"O�uJV)L
<b��$f }}.�x�"O�}ѧ瓧B��<9��c`��b7"OT3#K�u2�;��]�(^2��b"O��I��V�iQ,�s" �3�����"OVli5��tL�F��&y�V�Q"O���-V77Ѻ�3O��[ q "O`���`�~�
}P����D��y��'��,�RdR'���pPΉd�R�j-D��K�m��tL�Պd%�2=�"�%.D��P�
�:�L�d�͚9���K/D���);��yD�� $阦�2D����$֬]	���`�W�y���0D�L&K¹sH<!҇��>o�䓑�*D�챵��l�Dj�'Ѕe�FE�fn)D��0vn�53H��Q��;YDDY���(D��e�N�<�(i���Qb\R��1D��jf�Ʒ'�|���m�A���/D�K�$�!l�s%��/|��h*B�.D����Ǫq�����N�LՌ�P��!D�� DhC�"1x�Y��/q۬]!�"On퀂�عBׂ���D�>�� 6�|�V�h��S�~<����#IY�4��a��A5�C�ɜd1�7�O��詢$�%�C��LE"�1��$�x�i�iީU�B��(�U�V�\�a�����(���B�	�*I���HםQ���P��{��B�	=u(da��[[��(`����B�	
V�~����˔
}�`A�J�DڔB�	4�r���l����z1MA	h�����	�Q>��uC��A}j�x��P~��B�I%rf<`���5$5Q�?q��C�I5�r��c
>h�
	ؕ&_ �xC䉭)�F�qLX3uc�0����5ybC��+!�����W[��PO�1C�		zb� ��lB"��6(�	B|
C�I"��
s�	
�f�@��XJ�B�	u�ع��
RI��M�IQ�5xC�	�nY�+3�A8t�^	"BE�{�C�	ɩ5�9a��4��.H�S�.C��7r�����͙M��GO�U��B�I�M�b���@+.0P"1'_�B�I/J�NlHBц^Ϯli�.M9��|F{J?��
�R|��`�.
�ÈP�f�>D�����[��`�"B����"��&�;D�pУ(C�Q����Nŀ7��S��8D��Q��@���Q�*��k���b�+D�4AFƐ?a�p��s�c�!$D��"��*��RR
_�5��%))"4�Haw'�VW�b0���������DD{��)p�`B`���e"w��,x�ڹ��'D�d�vo�_��bE�:d}��J��$D�P���<0*SF�}C�rDI#D�h!	R�*ֈA���� ���5c;D���"NL��jK(	<�I��/:D���#j�Ot�U�'H�/S��U1p�6D���r�²tXk�n9��M�T�(D��S�'��Qi�K'���iG8��d'D���nC�7sVA�b�H2�T9D����\+U�M��D��c 8D��c"Ԇ1���4�Q0��X2�!D��B����+8�i91h��wȆİa.>D��8�G�kW&���,�i*'�;D���qk�#�|8��Ԩ{2�c@�7D���3# �Q��"�֬x�E2D��B�F�RW���V�Lx���0(4D�ȨBI9@������&0:֐��4D����`ו'ð�P��M%����.D����/4A ��X 	�,��K'D��ڇ���,i�h�s
W�_��PB�%D�X;�`y�j�S���A�l|�@�=D�����f�Y�7�k� ���7D�`�AI�p��1g�W8ZT��;q�'D�غ�)�(F(�,Sӆս*�(8ƅ/D��[�'C>Mx��r%M�<��T1�b#D�ȋ����⨉��8�� �bL?D�;"��W�&y�2+�\y�i�c<D�h�!�ɴ{3�]jw��Xi��#ï;D�r��9`�(��\m��H��9D�l����`�c�.P�BQN�M6D�p��fݔI�H�U�Ln���b�4D�D�S�BR�q����o�x��4�/D�FH_(��	8�
�Q�z��8D� Xfj*Q�����0��!E�5D�� $ū����Nz���"C��&�T"Oļ ��"5q��� J��~�"OPeq̒yd����RZ�N]y�"O���f�*�J�%͋�k$PmB�"O@���*�V� �K�'A���t"O)��\�@�޼Y�IZ�m<�DJ�"O��B&�[}*��ǿt8�y�"O,��V!ǅp���@Wn4�6"O��
��?�J� �o�j�e"O��5���T�$M�Bn�?
(5��"O�`��2z��Ԡ�M[��[�"OrY� �Y�:��㔁��a��"O�jW����u�dkJ�#^*|H2"O����En��c�o�x�S"O)�S��H8; $R2�&�;�"O�}�"͇�Y����6cݜY7N���"Oh��eK;#�z���"�-yF�:"Oވ91C�7cP.��D����@� "O6U��`�,"b�l	")� M��l�"O�� &�E��AP��6,�> �"OF� �_4Z�4x�� � ��c�"O��:#I�Mײ����"���e"O��#�R�G��%@b��?||�Aj�"OԬc��F�n��g[�L��HB�"O�X���.��{�G�s���f"Ol���ǡo+�E��  c�x�"OȘ�C�tE���&ѴU���c"Of�ȁ��+UX�2% %�	w"OT���ș�`��de��4�4"O܅B�d��7gX����	�B��"O<MIv����ċsE�0l ْb"OB�� ���4^�Y`p�)U�>��g"O~ (G���X{����ă��d%r&"O�d#�j��-�]����)��|ɣ"ODY;�2d������;��E�"O��Tϥ<�xP1� ���HT"O��� �V�>�#"��M����a"O��"�n!!$ô���#��p@�"Op�
�A���h @�i�4X�6-�o�<�a, %�0\��+��${�)BE�<�1�8Z���e�B�1^D�ʠE�<�� �, �t���$�&���j�nD�<y`	 >��	u戮R}d1�M�J�<I��Ԡv��
,�n!K �`�<��)]�:�x��3!�: ъE�F�<1�W6Ph#��8����m�N�<i¢�Q h���@�C�r�h�H^L�<���&��i�.S��иA	AJ�<Y�`� � �ѐg��@C�(Q�N�^�<	"�G�A�c�&��S��a'[W�<Ad�[�Ba6H��ȵ�� ��DM�<���S�N9X�y�� .��e�v&�H�<qd�ͷ<�Ö�&�k�N�<�sG لqQ$l&+��ʰ��F�<�A�P�b��Ea^IY�p����/B!�D \���d�9@��3"��!��ޣ%�6p�f�>*>�)�fօB!����`�6.(�Zg�D�a�!�$\�<�帠o��j����Hf!��P�-J��(�Sx�D�d��;UW!�� 
�@��ِ	��Pb��P�\�!�^�; �u��D��,ٲ���Oz!�* ��)�C������4Ӛ�!򄔭��Q�O�,-@��ۄr#�C�)� $�KAڻ/��Q�<(��$"O�]20W��bU`N�)�	�"O$I�녜&�Ѣ�G,JE��"Oly{ �ħx�& "V��k�tx#"O����U�>��"�?w9Z��""O�M{�j0a���ǇǠ}4� ��"O^QI`OE�5@� ��k�-r�"O.86A�1>=0�ɣ%"�ؠ�"OX<J�I���F$��.� IS�"O*�`b�ɸf �H%Dح,�4;w"O^j�'�%���1���3}n� �"O���`Y'Ak������teb�8�"O���0l�*����j %bLA�a"O�`-�<x"��7I�h%��"O@�Q�X�eq�a�Ɖ'=�AS"O���!��¡�wϑ�s΅��"O�tR68}ȝ��#�;l�T�5"O�:Nr�T�N�B���J��y�)�_bj���K���rσ'�y2�/����jR�}&�	�0�Q�yR�Q671Y����K��`&?�y�m�MxΔA'A��E�~=q�5�y2b~��=��&�=CR��N��y�,!$c����m
+��PZ��	
�yB���̙&�^uG`�	��?�yl�T���iP�W�ZX�2���y��¦�$�����}��1
ѧ��y��I�,�R�@QF��q ����Z��y���
DS�����J�k�V��Gf��y���!%�ɩ�h�f=&l;� ��yr�H�
�=�7��>^�t���H��y�j�,ˮ�zb��^Tzf��6�yr��:f�ŠVD�V6@@�/���y�$	t�. ���8LP��"F���yƖ4^	@�إ��ѪIGpD��'�h�:UFR8�I��`FI.f�p	�'�n�*���6��	���	)H0��'r�!ۆ�H:g�V諱D� r�p�Y	�'dF�2UϞ:d�ޑ1`��b��Q
�'�<�B`J�Y���bT�m����
�'yT��U�ɘ	*�E�a%�/;���3
�'�h�nR�T���F�@a�`�	�'��Iv��>q�$�q�'61?�D��'�BH�w�U�-�Р��ΰ. D��':-�F��n�V�k�τ1(�"��'�.t�#D۾����K������'�> :Ņ�uƴAu�IX����'�r��f�C/�ĩu&B�VnF1	�'fn���1f��l"q-��I^VL��'^Xrk��.]��\0Pc4�'�����hg�qb��F��Ia�'����d+�2J�h��W�\�M>j�'��8�HY��@%Q���6����'�8�W꒝0B� 0-��1�:�'p^�3A�Ց0��ɲ�_�%��	�'������ɖE�RqүH.,$����'*n,	g�е@�V�a����r�pP��'���H7��1s⌝����$�����'�$���0E��03"l�#X<q�'�8M;w��V��Hv"��(��1��' F�4cs��ē��B��	�'���ˆ�N4%�5ڱ,��\�	�'�.�!B��� M��ƛ� �]�	�'/n�� ��-<j ��ҸK��D8
��� ��1k�L���ʕxw ��%"O�����?y�h�J���nEh��"Ol|Zf��,��!��Hb�W"O���$���/��jœ�w���d"O�\�"N	�R���cU�W��V!b�"Oi�/ؼl��lQ6F����"O��C����FB���fKZ�Yc�"O��� ��;s��X1c*˛Pd��"O�Mz�c�>Z�.��JF  ��{�"OfM �ϙ��N=���SN�2U"O&�DڪY�z�Ѕh� +�0�B"O�@
U��x����*\����t"O���&�^�+^x�A!�*�ِ"O �	��سb���Iv��&pz��z"O*(@��_�_�)f�W`o�A�Q"O8 ���}Y ��E��(��Y�"O\0�Ӭ�k���Ҕ�M��[�"OP�xD/�N<<�t"�`O�@P�"O�8 E�-�Ȉh���%�&��"OH�Ц�dm���v� 1�P��$"O>� ��Q3ܸ�u�M� �h���"O��!��Fd��	
�5�f�[U"Oh�[w���
�J�FK7V��i+U"Ov��� ��ơ��G�J��S"O`}@�k\2*5+�E�=Z�ɣ�"O�9�A�*$�r�� .�4qPR"O$rAE�2,"4(�'����p"O^`yǎ�C:����٦SR��P"O vg�/'��1�ŏ/����"O�U��R*^rR�0 ��	S"O�Q��:�1�V�/!�N��"O�p��2���хB�ppS3"O����A�j������Z�cTa��"O�Ъu��6r!�r�A�MN�#�"Oĕ���ŏg߂�0֡C�e�X}c�"Ob0�#,)0~�����a�ڜ�"Oj�x'<��ʂF°xp�i�`"Ox�&�݈
�ĵ�+�gf����"O�j�JH!r�D�	i�4<c8�P�"OH���J�O^�{MP�9^���"O
��я#��5����=芕"O��J��W�f5\m��+��L�ܹB"O�1�O��&Gt]�P!E7x���"O�U#C�O�z�ȂU��(�T�C"O�2u�
W�R���}��ܢE"O2��bLL��
��‏��R�ha"O:IA�EP="����i�60e��2s"O�����4bp���]_��2�"O� C=n�P� ��AO5<q�&"Ox��G�#vzl`�k
2%� �""O�Ⱥg�!{�\�8�ꘞ2P���"O��3�ޝ0*�\�����\��"OJ��R�W�7�)TIP��@�j�"O��bu�߰|���z�X��"O�}�%�X�-��<��
�C��%�E"O
���!!��a��bH8q^�� "OJ�``lќm|�s$�F�Y�	y�"O�PGl���F�3� ý �:�#@"O*�zc��x����E�BG�80"Oj��Q�9�.�7�ЌD�B"O($Sf��� #���8�0q�Q"O=��BǕ)�<O�t��}Pe"Oh�3D�#8Tp���%?|m�%"O틆#�6���	��3�"O� �|�a�B(l.����	�" ��"O �q#ڱG�pYBG��S� �)$"O�H��?WV��t$ݔ@�|X�"O&ݙF���*]`3��eE���"O�pha���9yX� f^7X�l10"O�5R��Ј5���0EN?�$�1�"O�P#R���n� ���6��)"O�CS �>`�fK3�ɷ)��x�`"O0�Q���H�6��G��W�q%"O������G��r}�|���B��yb��2,T0kpc�D�QA�lY�y�?~YN��3��&hY��KX��yP�QT^�I���uL�t��J�4�y���7^�z̍fT��K�y���-��"V`	c��h�m��y"kD\���9����b稱�eB�y���B�$'�XEHL�E�S��y�B;dđx0lN�J*HA����y�ˑXh�+A$Ï?�jT���y�#�9I�Z��#��&B\
��H��'" F�"ov}�V��3g�X��'�D�+��6r��(��[�a����'�&)9@+^y�е{�GLf�]��'6|���
,vt�z�#�����
�'���(ׅ�P����9�� !�'�Y;��Kj���Ӓ�F�+���K�'����b/~�H1#�)�5 a��s�'� ��`NZ'^�!a���,.`x
�'tVQ�`��*��]�8tHl�*
�'PD���߷?�Rh��
�zWN���'�ly����b��C����@K	�'�����O����Kv�I�x�nEx�'�Ha��C'Ө���X"rblQ�
�'���*�/�UDР,B�x���
�'����Q�0M�,@.�|�� I�'���p#ŅE�D��G�J#t���0�'PHⳋ�8&�&a�W��b�����'�
0��b��,x���I��h	�'�}Y��ͪ&��d��s�L�)
�'������6 @r@c�qG���	�'�R����=
d�-��
�>!��'�1p��;�ll �R%�H��'���。y��ܛ��� n�\��'���@D��E����iM�x����'��F�݈L�hkwm�m�@�x	�'ބ��VK_�CY��yv�>q�B�C	�'������4LB,�DU��X"Ox*¬?#�`H��A�bb"Ot�{�/�҈��'��UZq"O�a��A�*�HǦɱI����$"Ol<��� s[���bOɣv���B"O����`�5!�0�%N�9<!��"OX=*PNGN���띧W�L��U"O�!�aLG�N�lp��@�l�Q�'"O,TP��_�Y
�����)�J�*$"O�H��.Μ7o 9JaA^�����"O��jF6$r�;�ϟ6	��y��"O�8�FI5h� �[Ce�%t|��p�"O���%������0Ik��"O�Ak�I�WB�<(�IL+Wرcf"Ol���͗0l��ay�bӧVP�"�"O`AD������	!��D���"O�+[�@�K�%o���W"O6q�ѱ"n���ʘ=g�l���"O� �ҡ�T���F�Y�Mj��"Oz$*�@A� ��q�$$��"O��i ���Ur��ʜ)>�2�"O����-G����[���"Ob�c4!I3F�lkE:GN�xr"O�dYR����|�cP��|;�I g"O�L)Q�Ԕb�Z*Uf��-�`"O��HPa��,�h����#`51�"O0ݫ-�5]l�p ��J G���"ON�ҖEֻkJ��b[� q��G��y��X
&+�,Rn�R���h��yB�ڪ!��@�X/R�"��c���y2#����τL��mA����y��Y�P��Q�΄@	��t���y��+*�>]Y��%K*B���_��y2%��k��x��"��R�L(r#����yR��6v��qĀ\.4R��E�M��y��Q�
*!�蝎|�Dp�c�1�yҫ��1�j%��ȯp>�t�S�Y1�yr'��m����%���a��+�>�yr�ƹL�"��NT�Z�����=�y�F4"zX�x�C�2W4�l�@m�y" ��kR����JCHբ6���y"�L�)���� �)E�
i��k�y�!/h�(�a��@�J ��ش�+�y�	Ԝx�?;�|�d���y"H�(GLU�Ö0�bx�T*���y��^��5��N�+N`c#&Pn�<AïW&o��8`T�>�Ti ��M�<�3ڍy_��GF�Q�r�1�*J�<	�`��Pu������H��Iq$�}�<��lFSʼ�V �t<�q�D�m�<ْ��+ �VQ��/�Խ Ņ�^�<Q�@_X��հ�ê_�e��l�]�<a�蜕/n9�O��]��0��[�<�,��Y�|�R ���>�ْo�<eaN&�(�!�
>�̫q�@c�<A���E4�]1�ڃ><�xC$T�<i�ߧ0�}J�N��j`�ea�d�<Q�K>\#�S��3qn�I�X�<��=kR�uKS%B�,�z%�MQ�<��,�3$��mF���h2b�
M�<Q1,̴c�����
�q*B6��S�<1R�ѝW��2�e[��$ήWܤC�I�.�\�iDx�:��@���C�I2Nz����A��6dv�Zco�,HZB��8M­p&)� �P`��q8B�	��eK1�ZY1�)��#]�q;B�I�k\Z0/@��b`{5%�'�C�ɴCs�f��}�U��lݯG<�B�I�A2�9�g�(�*hRS��=u��B�Ix����̜D,$@�Da�E�B��3sb |�c�[ u�M�T(؍r�C�	��gE�j��I����&�C��.M�8��0�N�@�D����F�hB�80qh�	4&ƚ}b����=%G�C��.[�� �/C���F�5��C�ɕqU�y�Le ���cE� � B�=u��i`����B�<�#c&�:*��C䉠t�ʨ@W�בV����+I�|B�	r��+��C��J}�ui#`B�I& �D���ɼj:z! F c*B�� �^����$Kݲ����
;n~dC�I�?��=
&�=j2�4�V/<)�HC�)� T9�	����T#�l$�s"O$B7c�2}t0��BC�#xW����"Ov 8$M���#c��JI�50d"O�Qi�
z�6А� ��gH�ę!"O�m�"�35��Z�A!G�#"Ohã߇0Y�Q�%f �);���"O
��p�Ȫ/'x��Ve�w�,�QD�'��d6d�=��W- ?�d"��L�SF!�J�Fh|��c�^�^:" 0�!4On�=E�aҸ!���Qk]�}�Xٲp ��yb��,zrD�$�(wc�dr.:���>�O��"7h�!z�lĊ��_���0�'T���&N8�n�9<��5joD?I!�D�+S����ŬT��.�mY:,!�d��d���d�J{n�[��C��hO� )I�m�:��#�?d�eK�"Onx%8�ȡ�5�م.��9��$,lO�xQ ��	�L��5�>$"O4�H�
K+@��(�D�j��݃4"O�+K�6p ��&cE=��J��'�\�dQ��T�5-t�z���2lO����V9a���S�A=����h+���S����d�%l�\Ls�)�"(ZjY	��!0�O�=��j!�D�D�=e��'�J�!&< riXZh<q�`��F�|yFG�[x�#�Gmx� �'���{�4#Q�F�C@��dݚ^�C䉛�E���ۑ#�:H*�BW�Z��C�I2���s�Z�~y���B�L� �����X�t��h%����r@�*Z>!��"]p���I��ZKP�w�K �'=ў�>=ZDM��z�\��愺VB̄�5ʔt�<����t���V����5bTg���'���p!c��VҔ�C ���7�D��e�<D�$���K�3���)�զ|l"�zH-D���2��>\��T��"G�F-�$"*��1�y��i�"��Z!m7��-���K�'l!�dɷ#�zڡ`K55�Y�tn(�!�	��RS�$]��a5.�?M!��Z�<��PN
��$�n�/{/!��A�+f��@Gc�~u����͝�/!��T��A�F�W�$̠��R�!��X�2(>+��P�Q�<��f�ȿ~��yb�;6���Qc#��8�d��@�12��C�	�(.t��'Z(��2@��kª�O�=�}ZWD�G�:y��6`ڔɳT�]i�<	#�
<8T��pO��C_�0pF�j���=�B"�B)sq��	9/���C�c�<��� ��,��E�	V\9�%Ǔܟ,���$QyV.�;IX�s0�,8 a��?��a`�5f��A��qE~���`��1 $��*�{eGTm�����Y�F����	Z�E�
��WN�)�����Mc�.�^�d�@��/~lH�J�`�I;0Q��>��(]�8��iABW����ۃH!ONb��ɹQ�L�a�h"�~�+��B��9r���Gy+G<�J����� ��c��׶���HO���< �	��[q��1gn��f�t:�A)D��g!�d,�E�Y�k�H��',O\m�~�>D��Xs��=_ ��P�,�=[�L��<9
ߓ[SzDJaK�/r��B�\4X^J�$��A��4�,1��C4(�Q�T�V Z�0B䉣[���p�,=����G�$���?1�Ig~�`��8��&�3.R ��F���?��n����k�&z?��#�ʀ9 � "O� .	��#T�69��C�GPk���1�	�P��>��wh�9
p�	1 ��	�`�k0D�t�a)µ.�؊��	����6A�<����Ӹ+��a飄�% j�q���یUSlC��#4s��+��ѩ;�����a�P7�#�S��Mk�H�I�>���гM0Nܺ��Of��'�S�'90�F�e̩��U)zҸ���4���ʕ�E�֤���(-� ���u̓[$�=�R@ÆDӼ}��ܤQ��L��*jڵ"�g_D*x���8(^�&�|E{���oK�D� ��䞾c� 0i��yr���:h���d�׋Ym���F�̲��'�az"��a=ƍb��A�:�q��С�y� �n�4� ��}}�d:�B5�ybI0�>,�G�Rrs��H�#��HOޣ=�O}4-�Qf�+������3�R���'H���0䒞E��)\&,M�=	�'�<�¡Ɨ��=���_x�8;�'%��˓�Z�*��Fn�<��ы�O���d��7�Ј�6��'��I)�C��Ug!�Dٱ	%��zG�V���l"a!�dJ�m�8'"C\��1�֋D?S!�>?�ne8e�œ�H5�p�[�!F!�$A-P	��&��w� P�BN ~�!���eS���a�7q7��a�.'!�]rv  s��M/�J}	���1�O ���/z�����6[_���e�!�d��KN����#P��85�R�!�$�3GgF1K�̈�eL�XJ��z�!�ԅf�P�����v>-�b���"!�$ól75�낻w������=ma}r�>��)&����բ�K����t�W�<�Ɂ�~QP��.:x1it�T�'��F{��n���4���o��XOF�zu"O�YIV$ڜ%�f1[� *LZEh"O�U�&ܯyt�r��s,�z�"O �� �Z��-�0��M!��"O�3`ܙ;�1B�O*l�%"O�jqDŶ,����e�ܝ}�P�J�"O�`s�L�>xbm)�F
�E��Ò�@���	�U��A¥OuR�x�LχC!��,y���Br	��6l[�L��=E��'@$i*@�{��u��@I
Q��}��'a�}�D�Q�^h�ipr�3n���'�p�C�k zDűA��;#�5#�'ɨYFa��;�U��/R�:�a��'/�!�QF�*�	�$&�83.b�!�b�>qI<a���'�uPSHW$Wk�u�� ��l��y��'�O1��4��d��
dq@�'�<���=|ON���CX����/ʰ%ZF+�S��|��'���M���HbWd�~����'�
��q��5o��qBw�L���	y�O�$#<��+��h$�l�����%YC�<�4.�!J^t�x�@أ <�K��@�<�fm(sK����
�4�P�C��y�<�g�ҎKR��5��0;d	P6�l�<p����aáE�l(�!J�`8��$�P�
o͂��PM�7T�$a�W,-$�p��%t-@'�X�'���`m��(OT�=�O���� �
.M״Pņͽ5�9�
�'E�#��Q�8�X��Q}�m�
�'Bb�MW�y��؋�FąLU �8
�'�\U�Ҩ�4:RT�a��M������'�H]���[�p������a��� �uQs��0Y����
ʟe�s�"O�[��H�r�.Q��韊V�t�2"O*�8W#�*u���ʄ�7q̭��"Oƕ���d�"]x������u�s"O�-��U50fD�x K[�n��"O�]H��9_�B����9`6��*OP���ρ��pP%!4��
�'ȰP�e����G�՜��LH	�'v0��I�
�4$1�n	53K�,P�'TX<�B�!�8�ԓs��3
�'Ǝd"�a�
��i#m�$:r�9H	�'D�Sq�(X��ybrh\�+��p�'���Z�@O/$jH�K�#V�'n���'�v��O���h�ۃ���8�'��0nF�^�R6cU,����'x���dȊ6[�8��E�ڤ`�'�̙E�P
&��|���9q�$(�'w�x��� 2k�@�.���	�'���Z�̀+z� ՛��4 �1�'���e�G�<�����˸bX%"	�'Ofi%�=Ԕ�	A }y�]C�'������o$0���ؾE�X�
�'��Q��ם����T'؁u6.�Y�'�H��b�'.�t�r�`ŖKb��'�^m�f׼dC��y���Aˢ�J�'���{���:�����8E���b�'U~(#���f�1d閺?ߞA	�'g|�!@	�8X4`�0��I-/$��'Ora�箍��蕘���1'����'冔S�N�`���D��vyS�' �5��ة�f�Z"�?��8��'� �F
Й5Q�-���/� P��'�E�7�7�D-�q�Q,�b�B�'�X���bC����wG�� �>��'�r��Ad�4Z��w
��$B�'��@��D$ත�yb���'b�������k�l�rh�~MnpA�'/D�� �P��qS�(/v��%��'�v�q]'U�Z�` ES�f�^t�	�']
إ�:0R�����]��9	�'s`8d�� (�� A\�P-4Պ��ty��#��5Ǵ(�tO�u��d�*�u�lu�ȓa�N�q&�A=]s&��K�2�ȓ�t|� -�.����� 豇ȓ1rAa�CB�� ��D��v�"���`wҹ�஘ ��l�2U<m�؄�r�pcX�`K8��H9.L���_� tc��НFB�5��١=��ІȓH6�8�!��:VTi7�4uP����!�t<�d�JܬI�k�l�Bl�ȓm���"�A�l^\���Ð�9g�����m�F �7j6.�M) ����t�q2�<<j���
����ȓ,�\�I��4�F����Ue�2 ��Vg�+�6*�J��&���Jm�ȓO&����M[(&y�l9#�]�Y��фȓ8�Ҩ(�C&;��)�2��d����ȓ{�f\Z���D���ռ~22��ȓKD�&��390鋗�Z;}B���h�řq��\aE��D�ȓs�� ��-_���K> ���ȓ�T�JfO�{����d5&��<��c��8���U36��K�/�,'�C�	�;�x�ju(E�d��p`U�x�DB�)� d�k�ɜ��|�Sg	� M~d&"OV�P���8Hu�䀖%r2I	W"O�����v��X%��o9�(�"OPp���H�lđ��� w�%�"O�����-[� ¡�34��XQ�"O��Ad(�SSd협�؝9�XY�r"O�d�tE�#�
	ڔ��=.�X�""O<�@����F���j`�ˋWyF0Y%"Oΐɢ'�7��h��~T$e/$!�dF�b�z�x�W7Y��Y�R���P�!�$U�"�^A����%�b��!K�a�!�H)I*"��uN92�ഹ��^c!�Ě$zʲ)�Tk����cV�9r!��+�X�*5�'G�`�Ҵ��fz!�I	߸ ��$vi��B&��;f!�@� X�l��qa��k0�.*Y!�$���mN�3��1m�%4!�$�%�R�Y��̜v?F]�Ṙ� !򄀡lM�щ�
ΌA��0�@@��O.!�$S�U��FGO�wc���ӯ	4z!�D-8�p "a�F���(���54�!���q�8���!�;Zk��Y҅N1Y�!�$�|���PS�)X%X�]!�Ć10���&�ĻL����2,!�d��Q�ْ�@�b���hÔ:�B�	$B�m�sH�ø�J�O1#�B��(7�M�C�Z�I�r}�#��ZC�D�4�wC�
+�t��1,;J��C創|�)��M�e�~q)�:�!��k���)�b
:"�lA#��A8!��ع^������ĵIc6�Y�W�k!���1����!�(x�d��'�0�!�$�t�.�³�P���a�Хj�!�F��a���J�'���3��K��!�۫=�M(4ꙏ]�`-��"ȓ�!��G� �h(���9-���aB+ńC�!��1+;�\ [7D���6��\�!�ރ^|�]s�!�v=vij�!��
1R�V���č�PJN9��S�au!�$I�*���j(��ev�C
�!��<e3���R���H�E�9�!���&r,<���ĺz$���Q}�!�D���P�Ё	�bs��*!���<4�ܨ��M�$6��CZ!��"_� )�lCT�Q�[*20�	�e���r�'by�6��}E0��U
�Q�	�`�VL�E�ڎ��A�T��M���ZFC��T�8��J�<Y�"�y�z,ׁ��>�l���H�;��b�4uS������2P��8;z�L�ܺ���aW"O6�Kb
�3o�x!B6k��HT�$�9&�)۶/�e����I1O�Q>7^�pKHM)� ��XBV�W�+<`*�$K��x���Zz>=+aDLd!���Q�=Z�0��GS�A�X�!�yi�I�aw�L9s�|Zw���*�$�3e!������X&,�
����h���=(�h!&'Vay8=ㅍΣB=~q�w���
u��
��S3_��(�׆~�<�O�#}� hƝ#��)��oߙ��ՙ�%�d̓�����%��
�r�ybݓX���9Q�:������(�4>ɚ�A$����Ѯkz�y#ɹ.axr ��5��I��ǧ\�`�Q��$	 2�	C�ɓa%l`��6�r]���)פ	:�9��
��9�T�6{����u�T��2hl�Q-Y�Z����g�L�����Æ�݀�AaE�xw���,L�_5lX�q�\�ّ/Ozŀ�%�bu�)6L��(��QTfR� �V��dC�*��qA����NmH�'ܧ�� ��I%�`��$JzU
Q(�pd��1B��L�T˓?ιi��4 ���PÂ�	����O�b��'��;���?g�|�8��	�
98(�@�ؾ�wfYP��&I��-�+=4��ʓ�*M�G Ǯu����Ó ��� ��m�t�CC�1**K)�<T`�v��81��$���!�q��9H��Y�K �� ���#Ĵ/Wr�`�T=�Nl��	�81��A9�J�+�(��ET��[ĨP���#q)�?�H8�E��@�m�K���N�;a(��d��p!$	7��-�8�"�F6�&���+<O�0�r@�2�2��s���t�0�%�tTi`G'�}aA�F1]�v�1�A�r|x�H���3BC�)��$?�����b$����˗�V�.�q`��N̓W�&�A��	u��i6YZ�vQ(u������'y���+�X��X�o����'�
1 �*�9/!�y����Lz,�Sh�<����9L��t��?�ZȠ@��.|�3Dʟ͘OȊD���
LH<��a�q�pUI�\�en�0+�'](������9���7�.)Is%�+>.�1`�_23�fl�Ш�7]*�����Oh�W�V3U22���l�59���@��')�  �N�t0�9�E,�"�<���ǟ�fuʕ��M��K��0�iS�Kq�i9&�i��	DlQ�Y����e�R�4��!sd6�	� ����G�`=�7� I=��SRG̐��4�؆H&�,BF�]�M��⚃�yR-<jM�U�ٜr�������g���ړ�Z���m52}>!C�lX?[y>��9��i�@%.�qj�KF/�NC�	>7gz�`5�Bz�j��lM�<�[#�V�" ���VQ?��9�l�����_�TJ������7,�~>�{R�J�L�ٷ�K�����H'c}��F�&r���an�O�|"����>�������c6b�ʽX�� k̓b�ȱx�΁)KV>e��>qɟ 8��M�p�Jdhħ[�s	
��R
OQȷ�	�m
�QCF�ɭ)X^�����,cϒ�f ��gq��'Ĕ#}�ep�����J?"�S4.l�6u��/I� ���B
QU
�  4���<�h��A0Ra{ү�� r6eRXQV����bC�[����d!.$�em��M��̇�G�`PS��/�jp��Q�<!j�o�ȹ2$�*P�4�;ņYv�{����n�$ �2#}
w�܁Y9r�)&I!H�h`�C�XH<1g@�z*��D ��HIt�ӞQR���"�IM �I�E&eEj��~r��0��0��*9� P�C�;�yr�Y!N�^p�C)u`5���	�'���l�:ԀBGV�zY��ir�		Z�=�E��n�գ�`+�����V�l�TH
bbaN�ժ��H3f1yf��:Z����D=R�����V=-��9w�_��APDF��j�G}��w]D���(_�S<(�hT�p�[+m�(�C�f��X����d;�ɫ7A X)E�(�0�EG��˓I]-�@CA�pҧ(���!��<I�L"��G�tl�B��4�S�~V4�����xB\i�G��*���O���@��}@8'?�p�3���@-B�2-\�f=��c�d6���Obe�
�"tsX��L��F����F�B�"���4��?Qg`���||���|��i�f*���)F|�,�>��殟`��r�v�x�L` A���.b ���$$�ɛ�t��1��5�4\�B�Ʋ�{���� �H�ҧ(���A�c�*���A����y
0"O��3W喭&�:]��ɕb����Ti:��I�`����t��*;&h�U�[�j.%j�K

M���dݺQ�g �B^۲*�8:r���훅�x�^��(0�I�!���`!���S���O@l��)�~[���aɏ�lft��'�� �l�UₐKФ:O��0A�t���I��1@��''v���L�xˤ�R�-,w�aӌ�$�OH�����mڦ��Ν;4o򨪱EȦ_��+ab�	B�!�ϋD�p�G	U��mHsA�	��������q.�B��y�,��:�l)x��Lw�.IB'�:�yRNJ^�ݺ4
ޑru~Јaσ��M�«���'���%��3�G)��2��\2��dw���'q|Mdc^Y�LA�� �2�4�?�	�sb �	�@�zU��ˠ����=D}2��x�}�桛��r�*Q�C:I!�d���x�<1a�a7\���bң:p"q;�(U{?�����&��e���ٱbwD���"�B�ɩ^���Ke�1O�$�ӆ>
j�B��,�,�Qm(5lM����\�*B�Ip����F�"��%B�Z �C�ɿ�@��V�^�.��jKA��C�)� da�q��=�D��Sh�(&"O�E�!\�,��,R�00nF"O|A!$��ռ]󵯀�A3��P�"O�G�#��l�2kL�X,���g"O�PI���U�a���W�d$��`"O���2��}L�<A�AI���D"O8�G�Q��H2� 9n�9��"O|�jT�� nV~�#�ǩy_�L��"O��J$�ڧ1����d�p�]�"O^�����4��ae"�o!� Y�"O ���Ć�͂L�҂^�k���{"Oܕ���	�y����%`A.B��X7"Oօ2(D'h�1�7��>��훗"O�3G
�7��[�/�=a#��&"O*�0�g��:,)I� �"OhB��Q��`��B#��h�"OP�1�Xt��]S�C�*�1p"O,�cE�]?���c?�Y�F"OpUP��ޞ-'��ّ!�9�5�'"O�0��G���u��.H�i�"O<Ћ��N@�#��cx��"O�٠�^�A���BA��<N����@"O<dS��Y6�:$�� �6<���z�"O�QH"�_�,�y�o�J|Vp5"O&����<�Ps�� �L(�d"O�,�0�y�N�"��A:��5�"O�6/�8��x&�ݘo�X�M:D�xAWgEQn�2w���5E� [��-D��`P�Xx���M�������$D�����,�����l���lps�f"D�D�B%�5�\q�t�P3r_�TP��?D��ȆT%[j��]?�h�Rf�=D����E��p���+��7?@$óI8D�8���'��a�CP7����cF;T�􈦤�=�(�^�/"�a��"O��0�L�77���M�7<,ly�u"O�i�CF>|��1�B�I��e"Or0�q��[��+��ƈ,e *�"O0i�E	u>���E3��]�U"O���4-]`[Z1�6͏ fH�""OR\he�VH��}�w��eD����"O�؈��C@���7&�>����7"O�h�A��ڰɧF��<��]�"OR�	#)Q"E�j��`�Nc��D�"OtD��HRvؽ�֭�)䨚�"O< �T��K�� 2�ö?�}b"O� ;sɔ!:�3D�ƍR��v"O
����ލE�
ԹkE�g�>��1"O0��#�2�y�e�ܖJ��d�Q"O����O�*0�6�a�̸�0�"OZE��HFwh  @�k��܀C"Od�`�U�h�R�!uΟ	�.h�p"OtCF-h���L������"O��h#gSN�P�!e�%Py��p"OR��R�*iC���.�5I�ލ��"O0	��j�)#l�ܣ�n	��͋"OvH�s��4����@ʘ�M�.���"OlIc\�d�P����JU��)C"O `��&ߕ<e�M"���(�{�"O���P' �>?��QF�En�̼��"O�}3�e�6Qx�ͩt�)q��<�$"O�M)���/B
�(6b��0�,0'"O��xΛ�_%z�� �n?p{"O�M�݇#f�a�&[�eK@�d"O� ����HϾr)���5b��"Oĝ
�Bn��	��#ڨU1�8y "O``��B0a�v��6c�!{[����"O��Y��1�`��<�|��"O\uX��}�,)��C�X�*�I�"O�rue�w������R��}�""O&� �cQ����d@ߪ{�B�r"O��)��!W���T�WB�h@"O��{��By���B����`��"O2����Y31�L��!�>`�"O��P6ꕷ4�DX����K�*T0�"Old0��J�%�z��q
�z�|C!"O���e�T�2�բ�Y�!���9�"O恰2i31�"�*P���u,���"O�!��ETU��53$c�"yzpQ`"O,�q�R�2��A$6�ô"O�1(��R�;q��GG^Y"O޸pr��)?0�H��m�B��l�<�C�E�8DDk��^�\�BjYj�< ��'�<bb����Pw�N^�<���7�p�6�NK�I8��U�<���%*��K�۷��k c_�<��¥\��a�d��&&i�e�D`�<$J�YbS��Pj��'@�<�c�"�NMj�hB��ۀNKy�<��݂.�<Y�`�.H�Gc�m�<a� } ��Q�J	k���d�j�<�QВ;���0� �bMR���x�<�g*�>_��z�Z�l�61���Q�<YO�Ts~�8�e'_� �+���D�<��C� x��M�f��[��G�<�c�V�[�u�@�F�t D��ERC�<iUn�9�LثW�܉�N����t�<9��ɳ#�X�c��H�f�E���w�<!0�]I�����0p��J�<��.�#f�l �m�o�L��fA�<�s�B,Q�0���
�1G ��4�YW�<C)�%Y�p�NR3~�xҁj�h�<Y�(P��p�H�-{$)�*NL�<���X*�$q1	E�*,��!FS�<���R(�f<h��'��q�t��k�<�1K^�F8`P`�,x���#��<D��h�C�\��:Ti�7Ӓm9��=D��0��O,_����'T>SLi:T@:D��e�F�F%J��S)ķa������;D�Dy%	��:��بT��Q�ԅ=D����K4d�8Xr˖8q�"���i$D���tbP�1���(�dS�g�z4#D���Dj�(v)XE��d����!�#D� �"i���pA8A�բ@k"D���lS)
RnE�WM�
�P�;q�'D�(2T��+ϲ=㲅��0$�"D����m�� �.����ǖ(=6İ�#D��P$�77w<\��V^�>����5�O\�pd�`���F�1F=��Q¯�9`���a�'��A`�N�W��uo�p���Y��d�IpP��ӈ-�Ӗa���H�AR������3����DN�`��� &�@$p�e�΋^И���)�c�
LWڗ�P�%�9}�SLW`4� E vtP\�`H�D5�#?�"#�)-
���b���&Ŝ�[���o�-X�)�(u H�kք��U�H����.=�=��![#|�U�@��-{<�Ɇ���m��|����B�/}2Ā�(g`P0��T�F��c��+]�T�Z!F&��(���gg΄cEk	�঑h��a���+XM��P��"E|�P��04k֥��T��;2�V4Y�ǟ�q�8�JT�A�I�F����:#܈;� �%��M	$`�
����L.l��E��A[nӊ@z�,����vX�Dr�q��h�!�a/��I��!�D*G㜱j���X3�Z��4lt@��b̟(QrP�	r�ƥSC���!�m�]��2��q:� ;�a�t�jV(��P��*D�s�h�5M��$����S-]�[ղ�ns�'"�je3�(�#k�L���dΚ�ʄh�a�7q� )�hԿ�x��1	�҄���<���С�)A�	�Po��q��A޿F* ����g��I�a����k��I%�ׯ-m>��%gӡ?p����+�O0��b�U\�؈C���3@���# �10d���iM9��9S��; r�'��C�4s�O�����C�EN��]�@a��	��8"0
X�#�z��"�
"��4�ӡX����(�M��g�M�����F��!��,<O
�R͈!\���1�9?��"5\��J�ԜB��$��ճ`�\�}�e*؁2B���E�D�d�DlaSh�PΰQʳ�6T���5�������G� ̠2��K*X?�Qy0�>Q55�gy,-/(D�&K�0��=j��^/�yb��u���� �ë�,���KիD�$�b����2�*�j��e��%�Y�(A7"2`��	;Z-p�ɇ���#g����
E���1,�*~�!�ݭ!̀z� �#ka���1���
1���	�$�Z�.�q�NV�(��N�3�"H�N̆}����$���y���y�P(���"Xa�-)��:+�ٹ`JP��=��O�QͧQ �<�dj�zB�YI+x�x�	���L����WHGSb��t�i��h�m�!������3y�0+�<ӢBq=�O8�;P�U�b6�� ��&Tp�[�DΡCX��`Z��H�^��☡s��q"V'+8u���"O(��oq�B݊aI�Jq�!R)d���A׊Tm�D#�g?Y��A�<;z5�e�Z�z leK�g�A�<�n�
��Q䇂a>��I��8��m�Ij4P0�'.1��M	��`�7���\$:A�x q��"B�w*7Y�a�¤�9��� w�ɡd�!�$M4X�N��W�0!��H

h��OYq�m�$��x�����<�@ܑ�d_#bN��F�E�!�>Ss:=�a�Y�sd�ZgF��;�l�EG��*g&��tg���p��ؓB��th$��`R�ȿ�!�d�Z��hAu���x1�T8O�T�DV���N�J�Ӕl%��gR\8���X�ab�4���;}���	8��ؗ��I�]c�!8@:T���:�΍�]�@S�aOx؟HB *N)�	HE�N?;�p�Y�2�!�4� �`�9���`���/�t`���`��_���"O$�3!.�D[­	�MB�"A�ܙ6T�d!�f�5%�9S�>E����\��H�0����녹�y�)���9RT$D�b����D���F�'�@�S�E�H �ϸ'o6颥�ֆ	��q��[,�r����>j8��u(�����o��K�d�� �)z��!� �+�O
`���6 hћ�N��{��1G�	�8��o�;��O���"�@>?F�ţƭV
����'�65�B)��P'L)vly�!+O@�`PE0nv^�J��|Z��[#�X�2�m�2&Q��P�@QW�<q�"N�iF.5Q�ϫ5�d��'�����5�l��w!K�g̓e��pz�Dý@���0���z1���Yy<m[R/	���X�*�"�Q��I�$��B�I"�l�	w�r?��Zpo�_�pB�	�^���@��T7jfp��\��tB䉀��D_�L�}�����.B�	&I�bC�!�c��V*[�pB�	�L층�2�[l�DS2 �'[�C��5Q`�����СH�Kr��C�Ɍt]��DO�t��
Ө?��C�� *#<�{�'Ĭq`��cȝ�N�B�_~m�҈A���S��X�,*B��pZ�&ݧ<���'��(�,B�	�G;�l�a�X�(QщN�2�C䉼.�yA����98%�6 C�C�IcA�%�d��69Fy�t��
�C��v���'�=�,��S�N�B�)� ]a7���$%h`�fg��WP����"Od�SAŉZD`�藇�kS��f"O�tK�)WR,��LM1!H�\K "ON8�Ѐ��l`���j�{��E�"O�U��l��oF�<����h����"O�!���.R���qt�@��ۇ"O�0If�*qA>��F�M�_��yg"O�l{Q�Ҥ)tA���B~kF�ѳ"OfL+��L��R&!�@�G[��y�&��/� �)��aIb��!��y���PX{#��*QԎ�3��^0�yb�q�n�F�šO�<�`�^��y�B�X*�ٖ��6ikb�����y¦� 	�I�7�ֳ?^�"g� ,�yr�_�����SA�^�̜���L��y�	9~���p�^G&�jE�ѵ�y�����5���"�0 �k\��y��I7逩 W���^m��R��y�B�y0����	<�<������y�aƸl���{U)�1-�5�y�HN�_@8@Q�<kZ,xҦ��y�e����ف��]r�̫�HG�yb'ֽk�T2�H��V��~�n\��'8,u��$��,L�`��qX$���')�5;EB/_6$�3/�l���	�'lJ��b�:I*ĩp�ڥY~]p	�'��9
vhR�}{�i�a�j�03�'�M��  `��]AW%W/o���J�'Z*)�l��? ~�)�&g�n���'��9��V6f>���&AߑT� �C�'2vd(U��
8���[��J��'�6`
e̝��ƹѰ#�9<�,�3
�']�=Y�	�`�q+ЂV�<�x��'0l ��ɏuu�͉w�D#0i�I��'3 ��9?��v���0oz��'_���0ѹz�:��d�T ��'��03u!_�C]PPE�ߨJ>�A��'�����+/\�H�T�B�NhS�'�L��'mO�6�����Ak�&m��'�����	{�v<bQ
d�f��'�X�bF��Pwv��3Gd�����'���c��!a3�\�'�\K��a�'��`��&��R��2�.U7C^�|��'
\h��#BJ	Z4�OjW�q��'�$s5&�
%ټ(�fcӮ��'C�H��{���ŋ8�� ��'��mZ�&{@�Fœ9'��i�'���k�#*�&}a�,p�'��tBFF.��v��u�$��	L����Fұ4@�F�G����L�7LI���ȓQs�\��E"0`Xv�| �M�ȓ*8BC��F*��t�!�]|\���qb��Y l�K���A�ȓlR<}!&Ţ{���H�|��Նȓ|�jIA�Ϫ��ɗH��|��\����~_� �b��?_��X�ȓ6�Р򧏕eO�yiGȍ=e��8F��S9���H�Һ�U��bB�#���}�c�5��O�R\�ON��Q3Ո������"|!^u�*OV��JN<���XM��|J��W����G��|IT�[2�AΟ�Pe�y,��ה>%?���4a*4IP
Ox��ç@G��@�)��@����g]=~�II>�꓇�(�P���ߺڞ����B�<}i�R� dy�ޒ�0|ca]����6/�9�r��� 2�K@���o�:����+���|�H~v.����a�ٟn2�����S8b�j1p ��)ۓ͆�l*/����� \���a���i�ǃ5��J�O�!mE�|0v��$~�I����ʧ;�zH{$�7I��%	�H�0p��+g�l���'T���Ԋf>	CoωH\|�%�)T�Γ0v���I-k���M��?��BӃM�bM`'+�,2F>��P�1��&W�-�ᓼ>0�M`R�C5M���{���g���O��[��-�)�+8F�Q�3�Ly�\$�TR��I�c`�؃���S.u+�q(�%�j�e{��	�/���r�b�0]�ɺ?Jh}a��7�g}�T9&fP�Z7��8B���q���s��#<�zV�λ��<���BR�5�`�C�e⬫��v
� �&���&Q�a	(��[�X � @�?�   �	  �  �  �  �(  42  =  H  3S  Z^  ni  �t  �  Ɋ  ��  ��  r�  ɰ  ��  پ  ��  l�  ��  ��  5�  {�  ��  �  R�  �  - � � \ �  -' �- 64 y: �@ �F WM �S �Y �` *g |m �w �  � �� ̖ Н � T� V� ��  x�y�C˸��%�RhO5d��p��'l��ɶBy��@0�'�F��L��|�t���pd��46b�Z�4?NNqhs��|`I4jE�M�6��"-_�7RN�wk��uGjY�7���
/Y���F�6=b�l��wm�u5�@%=,ĥ�t�X*v�"@�#�0 ��'��O���]37�,����M3����U�̳��A#['�QrDM[Q��=�2�I5'�lÚ8+J��E�Ql�6�\<9I��d�O����O����.~� "G�zʤU ug�%w�����O��Opʓ��d�Ot���OL�����Y��Qᄡ	�Nr���O��d=�d�O���ª1��I�<� �����8#�� ����â�o�<97g\�^�rZ��]�H��f`����:� �s���7�x<�O�)�	>t��Z��w�$���*�R !��WIL�w��O����O��d�O ���O`�$�O�'%�y	�ǎU!����:����I��M۷�i- 7�EY}rf�P�nZ;�M/�h}�@�X���M�3���A�W�'�a���S/b!jc�k_����lV���<9����*A����dƹA���ˀ��*>�R�)�^G1���)L(�� *�:���-O"��d��\������(H�Yz��#џ�'1�"t�M�4e��`e�?h��3d�'�ў"~r�7+�j����$%i�pA�R��hO��܉�Ƥ?EY���&�J�!���;D���K�O��O��D:�3}2ꉜWP�X�p �&+p}�7ˋ��y�h5o���f�)10����P��ymН�	KgS�>��ٳgKƏ�yb��q"1�N�>Y��"�(���?i��'�i��~�12�[!��X�����8�?�
�%�*&"̼*PÐ�}}0=�ʞʟ,��o���B�ɗ�Ik�|�� P/z��� f�#D�8bwC��H�8#���6sND ��#D� ��`^T�V�0%I�\���G�"D�@��oD�`$,<��다h�,� � �n^�>�q&��r�HV-	�B�"�����ONЀ�i>%�Iʟ�'`ʘ��O�� L�=p�lǇo5����'?Z�� �R]�q�A�	��hm��'I$�bc��..@hP ����a�'�v���ϊV�d����X36��1�'�VA��6?]JE�88����K�<	$�)ʧ%R����f�p�쳂r4�'7�=j��'4ҝ|���$޶^���q��!g�,"*0�y� Q�H���e�M˔�_��y�l�!uup0�擪d(�E�y"��\I0�(n��8�@إ�yr �/f�1*D5Q�r�g�7��z��O�����립�	ܟ<��ǝ��U�3��Q�/�џ��'R�''�i��箱v��Kx�.Ց$�͉;Y��b�ax���X�`h�y"�	+j�3�KGwi��`m�0<Y��ƟP�	����	� �p6'A�Xb�(8pa��i̪��'����v}��p�m�0.�]
�U�����R�䛐�شt�$��]�c���O�OB�N�^������y2�'��<KA��m������ӳ�n�E�'��j��,���{�𩓫k�
�!�@XS�)��(�.\��	��p�z���S�h"��$I��d7�P��F� ���g�nH�	؟�'?	�|M�i^��Cv�E� p��EȇW��ϟ���	�,fr��wK�6�j��עgʣ?1퓝_����k߯�"��� ҝ���D_�5F�������I`~�nWNF�B��:�%:�IC,�yR��1iw�1��A�z(0|)��T��yb�C#g��"�ŵH��T%��&�yBg��;\X`���ҡA�a��Y2�y��V�H9I�<�������RQ���J8 ��!C����)���@��e@8>��D�O��O&�O�'Q�g��s�@���̅T�����%B��x��ԛB����1_P���n��Kj�8q�'���Ƨ���ʰ15E�Fͪ1����?i��?a���?c����!ЁEy�2�"8��5P�L�g�<)�R�\D�h�CIB#�]C7L�{��M����d�fi�;�Ý-���[0�C� 2e���Z$�`�I�|�`e��� 0�e�Ki&h��abM&#���'����D^i:�Pˤ��S�Ib��U�L�ax�Z&�?�P�|"U�#�����-~:uI��U��y�o��,�VQ@V��BE~��`΁��?� �'^4T`��5@���v��bD�iQO>1�N�cE��';�d�'<�D�Q�!F;ǭZ�a��h���'tb+D�B��d��l�ܤ��#\96­Z��O���.����[?x��1k3$Rm��W�4���B���[��Ǘo<J���)�ņZ���ck�Bp��(&"ȩ)ò��'�� 9��bQ���'�����'�,��5膰8�|!�,C�~�>�cu�'���'�2�'�̩iD�h�$�j��Y�[�ls��D�[�O���%. �V�j%�D�@1��i@2X�X��m����4��q~�X'l(Г�F��V���u'\d�h�O�%�Pl@0�1�1O8p㣃��`�>}	�
	��
X��c�+���JTnű�)�3��G��q!I�qJAy��M;���O��$QW[~��'�<I�	Az�c���a��	<0d�	�'�P��R�é}		�"ĳ��݊(O�Gz��O�Q�<HT�\�Y��9S�N%ZW���ӏ�?N�r��ݴ�?���?q/O���O���߳Yִ�;��Sk�8p�!���d�i�I_�c��� �Χ55LS�&�̰�S�[�"����K�2��k�*�0 ��i�

��,pR�	:6��,x�NˑP���U)�����F��OD�Đ��m�	Sy��'��OD�gA�2E�Z�Ӆ悸@Y� �#�(D���4��7U>9BB'��.4FA�V"�<��~W��djӂʓ}]4uaeU����J��	u�h�&��1f\����؟��'@��'�Gޯ�\��gCː���O�i���8��Ɠ?��cF �:F���$Λ;Gv�`cc�/0��H0s���n+�=Q&�	+v��p��iՙ*�ȼ�b�V�W�x�=�ъ]����ɢ�M���sP���K�
N�2�g�U�)O ��4�)�'|�@ �V�ۖa�
exTCm�މ��I��Mc��Q�qup$���ţ��:�e���?L>���T�x�B�O�l�
�d�38�F,�bE!l�Ľa��'.��'R(��#�YԹ�EJ�F��I��'\*��P"�b�$�5���P��
�'�,y#���9B��M"���
�R�0�'W*�	�g��
Z�\)V.�E)��ć`�O�|`����wF�HHe#3��\@�� 4Dx�O���'v��� g�
��I�wOt�x5#E��6B�	�N��+wC������C|�8C�	^_p��4+F�Dp��&��)C�	+F�<q���Ǻ���q��o��C�ɻ]���'G#R�jtK��O�$K��cr���|z�dKQ]��Iqe	������Fhy�*%��'�ɧ�O��0�v$_E��A m�)c�0�'���PhВBTFms"�\�5�8���'����ؤURN��.���
�'��	����?��r&�-����'{f�Pf���BT��T�J����J>�q��<�$�I?`�٨��.0���Ta�/>L��>�D�O��?�'F���ȉ8F�b�٥��:�� 
�'�PL�Ь&=�]��@�x��	�'İ`�Ή�{gʨP�N@�{C����'P�qp���tI$�J�Q���(���E�2�" ���M9��H;#���hOfq���S�)$&�d��?�R=
Gk�vu���I؟���I'�Pa�J%^�H�Y�j�L�B�I�	�1g���0�����B4�C�+�h=Y�+޼Q�fM�R�\>Q��C�	tz�SC0�3/�]_n�?���	x��P�u������FM,Ƣ���'����埴��^~���Rc ̑��I��N-AP �2�y������!D��u�)���S6�y�ퟂ6�1��R�
\���
���y�.�D<KD�ژ[fF�1w 
�yb���Jn�aU@^ �(�֊���d�~��(������ݞz�!�OH�/2�� �_��hO��H��{�)�S�W��5�B,�p����,~�C�)� DU2U�ŝ_@pQ� b;w~�k"OZ�@��*�l��K��ڙ@"O�M;�H�8)蹨��]R�0!�"O�D�֍[�dMH`���d��Ց|�*(�͚�u;X�HìH,xۑ��
ID���q�I�p��O~L���=g��4�"�G�2����W"O@%Q��u���ǅ�9����yr.ÌP H���A�`�uA��y�힀=�X|X6(Y�iv�9E���?�5�'��y��-��W*�s���I4*�)��DSa?us��4�0�Ng(�2F�Uҟ��Iw�� K0d=-X̰r�KG��,r�K+D��Qp�.J�(����-n9�J+D��s���~��M҅%��y�@) �>D�X�iϫA����&N�9o	0��<�BP�>K*��$+j��]:!R�����O�4�E�i>��	���'�� �6��}Iq���Ϲz���'�:H����&a>M`r�I�5\��'4�xQǋ�,��U�p��4�>�Z�'��3�C�W7l��OF2+�]�
�'��+�Ċ	��
ぜ�7�`-O؅Gz��)M1h�x�Ϗ{P�x�E�ABf剃@�D�	ɟ�%��>�YW���&Gԥ�t'�d���)D����t��u⦋ԍ�0<��,(D���� ).��I+*Ѿ`��Q8r�;D��S��E�jTXs�	h|,�Sj;D���ڷ�}�e��H�H�e&��I�'�ڌ!�'D�2P�����QAhN!�F@���䓡?���L��`*�+b�L���� E*p���3D�\�����I�vŜ	�+�+<D����M�Y-�I�C��28��SB�'T�X�V�ޒw��8eB ���5�'�����-`f�Q��J�s~��!/��ў���4�0N��j��8��y#%� �������?A	�'`�[��լ�8�v�κAL���ȓ2��qGA��y�N����*�^Q��H��5���O�ibJ�CԾ�����k � � &�)"\�Y!��!~��DEr=ڧ��bG���XԘc
ql�	�	��#<�'�?����$�1y��Tb&'��k���ϢHM!�U!R|�I��ɚJ(��	�!�$J��^,�N�E%�����؁t�!�$��T�����H��~A��$*X��!���.�`�XVJY3L��bcU
@�剖�HOQ>9�e�D�V��QK,��.�[B��<ѱ�?y����S�'?c����U9V@�9�
�6-�T��Hr�%��䔤i`�8"M�c��чȓ�X���'B>F�"AlY�S�Nd��ln�UҔ��_&�I�Ub� �̈́�tHH��� ^iy�ǖ]�X�$������^S��;}��L��Mu ��OOYy��|��'��J߼ɲV 1��!#70��ԅȓ4r���G�F'�uY��0Gm��ȓ F
	����,nvm)�mL�/�^�ȓN�+C������1D��$�M��	�?1��x��U�w� ��L"`�WI�'ڲ�Ј�)�(�H=:�$V$]���B@ ˟9�B���OB��$D�].nh���]2���B�
�;!�ׅ���B�/NDS.�;���y�!�䈂d�J�Z�_2pv��T鞄i�!�Dz�`E�"I1i����A�NV�џx��i��֦1{�$ܹ���t�å<�����O���O0��:?a"7����_�R�h!H�J�<9� �� ��D���D�Wz��#�B�<� 
0�T�̾q� !���No�.�S"O�A�S�|<j�j���6�
��"O4�Æ�+B4�tQ#i�qDr��X�,ˌ��" �$I��e�h2��q�Ǹ`H�b�^�����?�M>�}�ElL����J�`��  DZ�<Y��I���L�e pp���^R�<��BR=d��񪳁�C	w�Ww�<)���@&����(T�e��ŉ�r�<9���
�Ȑ�a�F�WD�Y�A	�o�/��OR0[s�O���g�Tg�t�@�V��$	��'��'����>Aү�y�����"PP-�',�z�<Q�'�#�HH0�%�%dP8g�GA�<)#�: �y�@��<%(�CFh�<�B��6K���;�vP�7��h��py�C��`�� '��3��0�QF{�&O�͈�2)P�(G�O��@�`�*�zU���O���:�O���
��R�|�$�O2V�$�"O^Eئ�%hyL�IČ�$`>�J�"OM�7"�)|��b�D�d\*\��"Ol`�@`*8j��^)	L84�'��>�h��c��ijcl($F��i�'���ʉ�4� ���O���X��ML?kH�2�[[����ȓSa�1c@@��U*u�oR�@��7�P�%(ĝna�Ya��G�W8��ȓ�B�Qv%4�8��$'O������ɑէ�L�$!���U(�'��"=E��Ƃ3
��
w䅊#>𱹧�����.hՌ���OғOq�*�
5��q�ASF 6�XM�4"Or�ؤ˛z'����疨A��U"ON����?
8��晒g� ��"O\��D,�S�0Q��N�*�ޙp�"O�(@� �z�8yծ\P�*PaP�|"A#�;�V��_��`��J@�Yx ��ҋ0TH�	R�Iޟ���O�ЁC��6Uv(� �)s�����"O�����W�Tr4ώ�L��"Ov�w,�j�� Q���]R�A!"Oji8���r�<a�s�S$}��=��'���� ]��!�E�U]�p��c�<m\ў�Zǧ(�D����V�G�hl�����-��ݹ���?	�}��iU�D���ģ��DB�H��.Z��E�^ nx�0H���Ms�%��D�ڝ�ƀػ6��(H��Q&K�M�ȓp
9�T�̉O�f������D�-ڧ�x���S�S`\{����v��	�S��"<�'�?����]�WT�ͩS��D㼹�C �`�!�D�$"���� /9�p0ɑ�#�!���V�S��V#�������y!��؍]���7 ԁS�X�v��:!�$Ls	��l��D���4�ڈI���HOQ>ՠ����_��b�P�O8�{��<��e�;�?�����S�'|`PѲG��/G�ٷ� s~��=��(2�ԔfV	�JK�<Rr<��	!�0��<�r���Ȥ,n|�@�'b�c�d��aֶA�ċ�+16���'�T-J�INL �1R	ς)�HYIK>ɥ�	�9[R�	2Ln�����+���n,3z��)�D�O~�?�'OB��!J��f�P��S�?X���'{�1��*���GJ.Y/܅(�'Ƥ�����3"�:4͒;U.�'g�)Q��aպ	�D�Q�r��X�J�2�_1-��`��Kpf���ȓ��hOxp���:x���XT�P@�A�k	�������	m�^��vc�E�çv�Bx "O�y���?��4�f��a�|�CU"O� �r1 �h5\��-7iX: E"O�|��*5�r4�,M _MPh���/�h���9Wd��q� ��HhŬo֟�bT�#��|j��?��O�=*�E��%�P(E��I�"OlԘIJ�S�����́>k�&á"OJd���y�:���LDUY"O�Pz�G�����&�ٍf;<@�"O`�R&NF�1��V�'9�،CZ�8����'0�6uy!�2�+�ݯ�L�x+O���V��O���/��)���t����9�Rl1 `ǝR�!�B�hcHP�1$:K�Ɣq���d�!�DF�D��!%Y��<��A9�!�ܐO�����@����L^*!��٪U?�����D�+��Cs`��t�'9�"?�G%�E? !͖|�L	�&H��Щ����ٟ,%����A�g��E�;��,i�*��Fm2E�QnX28!��H���y��G[`С�^�W�!���m�L5�a���lz`Ƌ2!������I��ɂ��̙L�2k�O&�:�A��g�*�3B�[�[���vF0#~�@l��>M�5�!@�N;z�c�H���?����0?9n�-|��hR��.C�J)y!nu�<Q��ҕY^�Zp��k"�<��	Qq�<1B@�8�$�r�L�,�mzf�m�<a3N�'�P�0h�.
Jb-z"Bh�'�b�}*&���_MlaRaN� �Z�2��ܟ"+)��|����?��O��jac�
7?Ti�r&F,Z���"O��V�݉��q��	�8�v��p"OT|Y#�.��u �M�<H��"O��aS�+^c,���1�h�`"OVX:mD8o��m������^�HVR�!���5+Q��*�i)_� �;4��~9��ɕM��i�'nB%
 ,��3����y>��H���m���kN�)�נ����?���PDa���.<�`��"Ѹ~j�Osj|kD��7x��Pc�ќ>6l��d��U����)�N�R��0!�|Bu	�(L�4I橇���e@TMOy�'�(����?a������მ;T&�0{��#���'�O�-�GF�yp�<����Q0��'��˓J��a���?B����_�R�ɗ'�	��'���9O��G �u��	�z�a҈��i�X�$SX՜5�L�6�bL�J���"~:�,U0��+����>��͉E���<a���#Ud���P�h8L4��I�^X��G^ �Ta�&-F�4+�E�_��'��)�):?)�m��y�.-BSF !)��%Ň�]�<A@�	�6������fNx¥�+�P�?=1���8#%�33�6%Nh�;D�ן4���(;6�:�Ms���?)�����O��f2vsN%�i��6�TL�  ��:
��I&�TUЪHHh�g�'�pܣg�z��u;4䖐q�,\ڇ��']rW*w,��a���7���I�s�2A�t�U5$�F�U��a�N�iK�����XF{R9O�9���G���H�}{�pj�"Oȹ�Ꞓ~�l�i`o��or
�S�'P"=ͧ�?�-O�Ѩ���=阩� d�!�p��&��h���o���	��'�b�'��	�/g�2�I6j�1>*�`�cH�J���N/.ʘ#��N�"TH��D�4k "B�	�{N��cR�Ӫ,��5;gMD�q�V ��b�����󤄿q���D�s�H�2S%XZ�pM�񭝑z���If�'J���cnE9DR���L�0�h͓�'�6(����u��Tf�i��q�.O(�oZ�,�'f��V)�~*���dJ-Eې���	D\��c�R ���O0���Ol٫l-SC��C� ���4�n�Z�CSP=;`��OZ�{��ɹhߤ�a莳wJ���K|�A�ǟ|���@�J/^��x@���o�'3n�����?y���Γ64:ϟH���[�ͺ"[�����7b��Kq�=C�fe�'h��6�2���My�e��:����7Q�|93� ��dL�i�FHo�韀�IH��ퟜ�I�j[�aSE��C�D��Q����	2=?,C�M�-�:eh��?�O)1���5&��Z>rͩP�9w��Tٔ7O�v�Z�*�3�NDyL�c�
`
@ ��1�4\x�'��<�0� ̟�II~J~��O� �e��oT���q�,]��H�"O��p���p=8��Bǟ��eP�퉵�ȟy#S��1�ո��:V��u�R��OD��O@:�
צ��	�$�	Ey��'�Hi`QcՅl��	P�^;����N�^}Rh@f��@����SۖP6��v�݂��HS$�8�O�H�	������0�?#<�W�:=��b����a:�FLW~��Ŷ�?Q���hO��I�~�1��,�/ef�󈆲)�B�	�������,欀�wM�B�
��A���T�'�	* C��I���
@d�U��6�D-`%/!�M���?y������O���i>��T��)
@¸�@E��+�"�hYY�"a�);L�bdX��&lO����ԗ�F���o
`IJ�"��<&Ȁ�����O�b��ɘQ�z��YkX��T��vp6b[�0�u��y�'��h3�ͅL�(����o����.7D���G�x�ֵ2�(�<<,��B�<� �i��U����*p�x� `8�kHX��AabM�]� ps(	���?q�#�VH��U�/I2T�O�əR�H��,&e�m]���t�ͽ:�ja��C,Q�%��Ϯ! TJP�Q#)��t�%j�O6���O��Dr>�y6�ó��@y�D�!?jA�F�O�-�)�'f<CV��Pb"X�p�±U�B|��*7��:b�t���"�k���WD�˓�?���?N~������V�(��Pl�]$�MP��ɹk�axR�'��O�<��ɳ��$c�&#-?���Dg�\Ot1q���Ï!:4���2���r��R!U���D�m?�B!�]�T>��~���@�6�t�퍥e��0�L~�%(}�c��	2��'q7�X�s!#�8"ƍM����3w#5}����G��'2���ߕ% �i��&U�X���ԎS
��	+��
Wh�'}|�N��1�d["x��A�̴�	2COH�'�i����
�x8��d�;���;�C�\9j�d�!+��U�S	� �O&�oڟR(zIFT¥��n8�*�,��O��E���,f`�R!˅�nE�)4D���ɉ\.�ҧ�9O@t���d�����S�~`y�E�ٕ �h�ф��Qy¡���DH��H��-��S�D����KI�+J1���'B I�[DZ���9OH�b��ON%��2�8��T(0���X��'��}����
��� 8[V|�����#�PB��.��f�GdE@x�5)ۀR�F6m�O��O �����|nZ�/��tYBaX�(bԡ�X(d7M�O$�OR��Ϙ��ܴ&�Tu��K�"T��H]�V$�HD{����[�$����$��_����",���y�(?K�t�	�g��Y���yBE���D1��ח56f]�QǍ��y�H�6���3��M�:�bX��Z.�y"M_1s�& A@�ͧ[�j�s#�$�y,��	�q���+	�ظBI1�y��J�z�(���T�U��:�y�P�Bs�7#��Z������y��/w[x�ALȐ*�d��*O-�y�	�{���P�uJ�E��C?��OJ���O����O��DԽ|�� U�R��(�aJ^5R��=lZ����I������p�	̟p�	�����!Z��!�Ke� �!�b��hc�!�޴�?���?y���?���?���?���o����28���D�!����E�iv��'�b�'���'&��']�'l�P�gg8]������3�ܴ���'}2�'�r�'g�'|2�'�"�'��isJ/
������j�1P j�X���O����O<�$�O ���O��d�Ol��A[�lN8�e��Q��8������E��ȟ��	ҟ��	��t�I��	꟬�e�3G� ��J�9}���A
4�M#���?���?Y���?!���?1��?��h5~�q�Ă�&�4�RK��y��'���'T��'���'���'�ɏ�I���H4Sk��Tr!&�5grv7-�O����O����O ���O����O����l��`7�����1�I���Qnڟ��I��I�T������	ן0��,B��kW��I���حWi�)��4�?I��?����?9��?	���?��p�0ܠ��ۦU�=ˤ��1.�:x��i���'���'�"�'�2�'"b�'���TiM����"P(�f���%nӤ��?�-O�"~��gQ 4��D��ԩZ�Ɂ�����<�����O�7�l��(��'��dQ��ƻSrF��w��O���l���'M�O;�	�úi��$�0:D�q�"G��
�'��9b3O(�	� ў��<a�F�6^����VbȎq�B0faCȟl�':�'�c?��	w�? Ұ	�I�|�^�1 �T�L(��`���V}�'�r3O�)��Y5LH>Ub�+uICR����?1��&AJ���d��ş�s?ODDQ�#�z�I"N�{~YJ ]�d�'�H��-z�UY�$������OjA�'��I<�M��r�O�h�Ф-� ��u	�ARk�X#�'���'
��	������'6���� �a��$6:(�d��.	i��Iߟ\�'�1�N,���(M�Jl��Ö׸��'\�4��O���?A��ħ� 5�*����*L&����F
�_����?1��y���ҫIġ GO�c�}b��@fW�q�5c�rT��(��'䨬%�$�'j�A�H�L���HV�i�g�'C���y��A���swÎ�@��	�PN�$�?ɲ�i��O$�'�B�id���*l�aǠu/*tHD|�xeh�i��$�Op����
��*#d�<��'�y'Q0U��l� �QIV�����?Y��?����?����?9��iY,�� �c��:�(�V��B�"�'5���>���?Q��i�1O��*��G� �܁���C~@�&�|��'��'����i��i�e+qhH�
��B��@1o62���ȝ��������d2ux���#\�8uhQ�bKѴ#Д�?�wW����ǟt�Iu���Ȼf��F��O��m��G��Đu}��'*�|J?�Rŕ�s�:��DV38�Pm��N��U����q���'i���v?�M>�7z�n�A' �J1�tg�4��?��'R�`E�ã:����)=4PxX����T���?��\���4���3v�Y�x0�X�� �(M��AӸi��6� �T��7� ?V�J�w3��) ����Լ*�zl�&Y�`LR�+)3"Q�t��ڟ��	ʟh���,�O�ʴ��,ʵ�\yhD�Ŵ#7&y0�X�4���8��I�s�D��4�y�ߧ^qIq�ʁNf����B%�?������3: h�ߴ�~RI4K�8Pu��sb~8�G��?��HPv���S�Iiy��'n¬@�z��Q�fJR(��"�+""�'2��'+�	 ����OP�d�O@%SrhXQ����Q��V`D=��7�	���d�O���?�d�#�&���9P/Bb��\!�w䜽��(�M�Ő�MQ?)�'�< d��)�<�%����?���?����h���	)o�lHXS�X�V,(tb A7o<��d�H}bQ�0�4��'U�DA�'s$uA"��A+.}���+�2crӤ4nZ��M��$S �M{�OZT*T�����$G1 ��A��h\ xg����\�yr��O���?)��?	���?���r<���7}���
��b0`t�-OP4�'���'?2����'`��bb�_4[.���#�r|�B �>����?�M>�|�fa���戈l��! ��4��%JM֦�S)O��a#/�~2�|"Z��0B�U�
���P� ,Җ��Ǉ�ß��I����� ��LyB�>Y�wL���7GB>쑑�Y����%�f���{}"�'f�:Oz���,D7 o��`sᚑ��,�!bW,2՛���sR�F3^'Q>�;iQ���]�-��(ԩ��>6�$������ȟ������e�O�1�eH!MeTx�Dp
pI����?��
q�	G���l�.b��g�]��z�8UCH�<��)�@!�D�O��d�OU	.t�*�I���P8���F_�]Լl��K�QUڴ0�Op�O���|����?y��Qb�1bl	�!��-��P �hqQ��?+O,��'aR�'<b�?�����:� ��r�*~���<��Z���IަRO>�O�Z���jքb��ի��\t�̔���Ȯ��6�\U~��O)�A�	�*4�',��b�@�Z�Y�����`�'7B�'@�'�O�
�?IB���Q/�u��Hɸ	��`Q������ן�j�4��'�^��?��V|>������8��ຑCZ��?���V��02�4����X����?��OטH(Ռ[\DBhE���̑���$�O|�d�Oj���Ot��/��aЈ'�4���	�VX�q(�O�����O.��OB���D���;� ]�E-�;;�z�O��hA���M�S�|J~����M��'�p	sÓ7JĪ�H*��ܡ�1x��A�O���J>�(O����O���ǀ�J>�GA
j�l���O(����i�IUybú>����?��4a7��v
�{�g�
0<��2��>a&�i�6��^�	�Z������WFH�UɁ����ɟP8�lD�#��Șq+�yy�O������(��d��>��D�n9AD�W�!��p����?9��?���h���0/�<HPKë%4�uX�@81L����x}�\�p�4��'���c�ź!�-��e(p����R�{�"�m���M������M��OT�T ���j��ɨJ�Lhp)�n
T�&ڕ8U2�O��?����?����?Q�]�,����ϻ6� ��'��Z�܅k)O��'���'�����'��)���!
��B����T��9��>����?�L>�'�?Q�
+�꓋�;M*)��͑z}�q��
�M#�O��Q���~b�|�[��Y@I�9�.1�����Nɚ�G@꟔�Iğ����h�	Oy2��>����� ��t�(N��Q8qCQ�e�@1�'
*6m3�	�����O��du�ē@���%�9Z��úEP������ ZJ65?Q2�6W�"�|�w��[���{Qz�� ���� Y��?���?���?����8�hP`�ql�)�v��&���'r�'p듷?1��V�dĳU��tSd�Z�W�0� ^T�'}�'\"$֚I�����tn�&2
Q�5��.+�lP����)��Ov�O���|z���?���'�Z��D
r��qƑ�(�Ra����?�.O�T�'_��͟L�O����挔%9�8	-��O45�/O:��'��'2ɧ��!�,��)���e���Ѝk��q����7-Jzy2�OT�����z!�>2bѹ�ܦ`���z�#�O��d�O���O֓��˓d�riZ4`@P-��Ϟh|�3�+Q��?!.OlZY�l�Iٟ�@i
r��0xc
�H����E�ܟ��	0�:=lj~Zw��pCڟ��'1ERժ#���t��QC����	ly��'n2�'���'G��?��H!�I�uH4 -��K�@}2�'���'���yb"u���I=g�4��RO�x�~�z�%��D�O��O�����q�A|�t����%����T�qq�?�"�$X�("�'>�'��ϟh�I<QR�+��S���)�F
@L������I��'����?��?�Uh�.�h�����8��k����'5x��?���']
�IM!h�z��>O*�T����텆]�4��Ġ.?ͧ�n�d@�yҁʹ�p�&N�#���PdК�?a���?���?y��Ib�¤��5>����Fß	Q�8���O��'���']7�0���?b��%9dLzb�P�R�n�T�؟P��48N�&�t��@�*i���џ0:5�NB�$��
|�A&C'��\�a٫8N�x��|Q�@��ߟ�����ҟh��O�O1\�Z(O�y�,e���MPy�h�>����?q���'�?��C�� �q��d  ��sOֻ+�����MC#�iv�O1�H,���U0Q����FxpY�����s�����.A�4B t�	Cy��=?�k"��hF@(tjsA��'b�'���''�	���d�OH����n�4���E#s�\���!�O`�mZd�3h�	��Ms �iA~��/}(,qք�UrD�rѣ����J�in�	�^�i��OAq����=(C���7e������I�Lf����Od���O��$�O�$&§*=�ɭs�,qjg��(BG�'t��'S�듛?��Z��&�d�e"ɓ/F�>�҅����\+dO����OF�)Ә4|�7�;?1���8��A�r���_I����O�F��6������'�i>Y�	��I�3S�]�Go
:FF6�Hp&�	 <N��ן��'�ꓮ?��?aɟ�����u����� �W��[�^�`{*O���{Ӓ5'��@Rq:4�ՏE��0,�Y"n�
�%=R� I8�d>?���p�&��ȼ��p�9Ɯ`\�,;��-c�����?A��?I���䧷��hiCG��5�6�DEμ^i0z���Ob�D�O^�o�C��<�����M���:�@p��?�V�!��A�;P��g}��:dӈ�<�vq�k��B��\X�. �Դ�z�g�*���'��	�����џ��	���I~���=;Te����#^��b+�,=�I���I�l%?�&�MÚ'��c�c�;3�,�E D�e(����?�K>�O~��2�M�'l�I�1�iUZ�
�NĐf Ա����Ge��0'�ė��t�'<�$ڽV�L�(���$�P���'��')�Y���OV�d�OL��B+=���l\K]H�"�,h�⟬��Ozm�(�M3�x�O�n�~�j4d͜N�4Kf�	�ɑ5�:�R��=|$?�J��'8|!̓Q[��h2�g%	) )K�
��	ϟ`��֟��	�O��D�'y>b�(ւL�P~�I�eX�,�B!�>9(OrAmG����P��a �i��]�b�Pciև�?��?q��7� ڴ���Y"'��\���r �1��.3��PC� GX �Ɯ|2[�4��؟�����	��x��ė�HT�ҷf˫"�H=� ��tyBI�>q��?y�����<�$��=�Pb��OXh�`�cG�T ���|��Y�i>}�	Ο�����Q�pZ4��/n���P�G��A`l�mv~"B�)V����䓨򄓿{9�})�A�,+�4n�F���$�O^���Ol���O��S��ן0K��I��V���KQ�3�V�QPҟ��ش��'�.��?��y�<t5��z1Μ�<P����޺��޴��$ uD�����i�ٙ�-1�zM��mA�`ŖA@T��O����O.�$�OV���OB#|wy;���f�\5�&�ƅퟨ�I���On�{ԛv��'n��)�6폹yr�e��JB�'���'��O�6��D���۫ g8m����9k1�c �̟j"Pa�O̓O���|����?���Y�h�"!�3�P�bG!5��0A��?Y*O��'i��'���?9:�[.HaD}z��Αm�����<��Y�H�	ӟ@'��Ot��hPb�2�<��"��"R}�_>�{� j����V���T%�Hː �;B+h�p#��50��Ɵ$�Iٟ���ʟX%?E�'tR�� ��
�,��h0���ՙX����'�b�'^7�#�I�����ORU2�苋e��`E�C�R-����O��DU6(?��t6 b?�uƀ5y&ha�GɐR�i$��Oʓ�?����?����?������4U����=71<l� �Ŷ6�듐?����?1I~�b.�v2O�i�-n�T�#� W"���'pr�|��$�T�R���O&��Ub��Y�@Ңb�Ai�Y�g�'&�a�(Ta?AK>9,O�i�O.�h���)u���qU�j�����O���Oz�$�<wY����۟�I�f&��cA�&X�ʇM�4Vl�?�V��	ʟ�&��;/C�<��|��k�")j�i��D^y�m�1Ul��Ӵi��i>Ź��O�扥!C�٨%��T:��]/��m����?��?���h��	�H?.(�Fk�(.E���PJ��@*���~}2U�X�ߴ��'��T��v2���Ǝ�`�^��*�s"�'l�'�b����iM���G=V?�R��p�rHB�mZ%e�6e��d ��<��?���?����?1�L9Z4�x���`N��*����$�[}��'���'I��y"n[�a&f�󋍓&�Z��P�˿?��듿?�����S�'q+����� V���1]�V���1���&
8��'��*�B�X՚|�R��ڠ/��r0��тX�U�n�)2�ş���۟�	ݟ���Lyb�>�����u�y�̘#W13�lͫ��o��F�$�g}B�'&b3Oluc��V�*��eMY�7�Z�*�)�_2�V��j��L�[��)1�ib�i��A ;R�)%��}HCj�O&��O����O4���O.#|PБ2��=��cHj4��K�ş����( �O$ʓ,�6���1w;`�EBێ]����	_� ��'���'���c��i�iݥrG�C�<G(�T�_3~nĩ���@!>L������O����O�d��U�Z-bw(
n~�K���;����Oʓ?�I���͟�O�����	Ѥ4k<\y0Mƥ{��q.O~��'���'�ɧ��5�������A�BU�g^*{��h��8*~V7m"?��'R��	h��(\_V��a�JI�u��#�( �D����x�	˟���u��^yR�O�M!�+V�g�:y�3�ݧ����'��	��M����>i��nl�Yx�&[�<�� ��*hY4,��?���@�MS�ON���@%��Oю	��,�ԝ�E�X$*l� ����$�O����O
�d�O4�� ��oՆS��)0A�1P���$NG���d�O��$�Or������̓ ����쇉G�Z
R�T�(#�<���$��$?�Bsʘ����pcx����Z��đ�i�l�pQ��\I ���O�O��|��7E�WF]�!��Q�Đv h����?���?�/O6U�'s��'���6��=ʂʅ����m� 	��O��'�7˦-�O<��F�e�x�j�Iɣ~h�)cj�����h��J⦄�D�i>Mr����g;O�!x3(��)�@�8��˭Jz�'�b�'��'^�>-�1�.��e�ɂ��DH�a���<P�I��D�O���ئ1�?��'=�$I��F��i�'��A�������?1�^��F�Zܛ�>O���߬c.��'�u�Jk��b3KSz��y�I�������O��$�O|��OX�$|q��I�&_�O �I!�����ʓm��	��I���'?�ɫ��Y�k
�<�4AFHL I��5ʩO �mZ��MK4�x��$��,
ԂDdV�?P�	�g�Ce��.���ԑ�P'���ԂQ�|2W�y�g�s7�����X"^~ �Uτڟ�������֟��IKyR��>9���D �G�Q�Po�Ѻ�-V�$N\�1��R6�6�dM}r�'���O*HZEƫI�%{� ��X�u�T�	��6��L0v������i`�I{�LB��ʠ��h��쉀b�O&�d�O|��O����O�"|�#�H����p��52�ܻ�d�Οd�����Or�d�O�|l}̓ (
 �����z��sc��]��hH<	'�i�r7M�Zq�3�b�:�+f��H��(����Рֻl�z��Co�6!���D/����4��d�O6�D�"mD�Hp3@0�5�N�g=B��OV�)i��蟤�����O����pg	�K���t�j�A/O�$�'~��'ɧ��'R@k$�[�� ����ZB����F)���V�i��I�?��F�O��OL0�͔	�,���è[��Թ1k�O��d�O����O䓟��h<B�)�%i$�C��<���/�?����?ir�iF�O6T�'d�G޵?(qqe�ۜ0ج�����B�'ȖD��ir��O4P��*�7��s�l@dbH1�^��Q�`�	�՟ܕ'��'v��'���'���)h2�t ����I���k�&=,�\�'U��'���J�5͓j�Ф�B��/��3Я	\�u�IʟP'�t�	��P�I50�]m��<Iţ��3r����'�oO��2�FN.�?1#�{���y�Fy�O"��'�(��BbM�9��u�!Ǯ"x��'p��'B��'����O��d�Ov�ˑOƌ�8�ˀE��l8��M.�	��D�̦q��4Q��'2�cU�8���ЁM�<m��H��'%R��+�����H������5���	~�0=X��DW�)h�+�X�d�O��O�;ڧ�y
� �8�n��,+>}���˟KT����'�f����ZЦ�?��a�8#�Ί��T ʕ�Q6#�t(�Rkz�v-mZ��>�l�[~�kɅl*@p�Sg�f,�W��ӓk��;�Q�|�[���I�,�	��������g��-����bC�i��dk�F�Fyb��>�.O.�>�S6x�q��Y��<��Rb�5r��s�O
)l��M�f�x���
-9���S� �5� �5	���g͙1X�	HM$�G�'�`e$��' ���"��	 V���bt�'T��'�"�'��Q��íOl��Cz$�5���S�0L�A ��S�����æ}�?1�P�̊�4t��g�O`��I�`i^��6F��"������9ۛ����-��Y��$�X�Sܼ�gn�0I7d
T���Fy��ܟ�I��L�������xG�t� ���ʘ� E`&M��?���?� ]�|�I����4��'���Ŧ	C#�|
�d��X���J>	���?��%@:�Q޴����v��E��<��9R�J�,x��p�@�*�8��P�	Ty"�'�R�'"C�/����qꅑ����!�51��'��	���D�O��$�O<�'_tQ)�*њ �^4{"��9%�q�'=ꓳ?�����S����'� e�d�P�DQ"m�H��z�J�S�`�<��'S{T��z�I��0�PQ�0fe��P����T���ڟ��̟X��k�^y�(�O�)�v��I�p��	�� �H��'u�	0�M��b	�>�v�i5� �f[� Ŭ]��� �S ��"��q��doڊ~�l�A~�&ۋ ۪A�S�S
��/�l5A�o�c��H�FK^,'����<���?I���?���?�͟���G�p�֠�`���.������>����?q�����<�5�im�DS1t�,y��I�3?��t�mɏ�67��}BO<!�'�j��\.��ܴ�yKR��U��;0I^��ǎ�n�-��=x�����'y�$'���'���'����2�b�*�E�[�}_�ӆ�'�B�'b�P��O��$�Of��(0�j��CJ	�*�(��C�!u�
��#,O��DӘ &�,�`���m^�E�S �y!L=�È�Op�DV�s����38,���?A��'zX�ϓ|��4�PnY�S�y1-��g���������	��	q�O��D�%`#�_7~qt��櫏�r�"#�>�+O
�n�N����юC=B�8��
�4�n�҆#+�?���?���W,,{ܴ�yr�'a
WW���S�i�);q�ĠLX� aB��b���O�ʓ�?����?��?���u�j�I���Pc6��vE�,ɲa�-OM�'5�П�&?��ɇD�L\�0 �4��Nܲzc�Z�O^�mZ5�Mv�x��D G+=YG"�'Z9���s����d���P���Dď9�����'KJ�O��ST�w��!A��ɱJ��=������?9��?����?Y/Ol�'h�ΗWV@��+X�Gd0�h%
ϗL� e�h�pY�OHil��MK��'����oL9~T���fN9w������Ď�MK�O��F+�$�J��?�l��&��y&E�:��\z"�'�2�'u2�'%��'�>�4��9H0�s��4
?��Ȓ��O����ON��'_r�'�7�4�I d�(w���Y�B�B��}�L&��nZ��M�'�(@�޴�y��'+�"3R�	�"��Vd� b��1����!/&9���nD�'+�i>���������EÀ��P��^��	9Q�Go�0�	����'{������O��>B�(3G�P�������5�4	�'~F��?���S��ߞn�ڕQ�(A-#ڝ �ϙ�����6m �Y��2�O��I���?�eH$��X�!���,��?7�)���0�|���OF�d�O��=�ɵ<q��'RJ8p��(d�� c2@�;k�����dB����?)2^�\���r��Tౌ�S�� z@ R0o%���ş�ύ����uW��S��)9B�'P�b$�� �@�?������@�'��'��'r�'����)�Y���\+!*$4a�kTDli�'��'����'��6�r�<r��W�i�����W�q�N�O���?�D2�	�R��7M��hp��ض6+j C��U�-�6�O�m��G2�~�|�S�������si�1f��-��K�Lh�(�n�P���� ��Ayb��>a���?)�N�0��D"Bu	�E�@֘P��=��rϳ>���?�I>���JK��0��]��aߖ���`�|��=&?���O特�v�k�\�������n��D�O����O2�3�'�y2�߼G�X�pv�ʞ9�l��jW>�?I�\����ǟ�ڴ��'e��
�:Ap�;��۷?�B�N^�:c"�'�R�'���9��i"�iݥCn�o�c�|=uS�/͍f2΍��c4EؒO�˓�?����?����?��+@�#�- �e���6��?}%�:+O�e�'�"�'m"���'2�L`eg�k	2����B0R>И(b��>I���?�I>�|2P.�)�2qr��W�<�s�F�TI*ߴpF剝{Z����O��OF�';�A	��	�}�ћ�m͊K�԰����?���?��?�)Oļ�'@c��R����X�<�Z��ړ&2BmeӐ�J�O����O�N�kx��d�՜&������sT��X��l���-�Qa�l�?�&?�;k���떫��>���6De<��������	��p�	N�π h��&2G�1)�A�sL4+�'���'�x���$����<�"�@1]��+�
E�:><9@GBu�I�l�	��8����!��?�6��s����3b��G`���kL�~�x�I��8&������'�B�'/H�
�CE<B�8p�]�!��R��'x2T����O���?y̟P��CB�K�b$2��
y��U�l��O2�$�O^�O�3lJ<�s�J9TN�M6e�g���8��İ3���n�V~"�O�̼���pVl�X��3*�$��p���Q��?���?����'���ٟ4(#� 2a$�Xb�%(���²A�O��J��f�D�e}��'�}� �l8P����joD����'�ba�G�F��ತۆR���LHeB1F���
ِ[c\b��'!���p���x��ğP��M��a�Wf�i`C�F�0�02A8V/�	[y��'�� Dl��<y�/�Ж ��!|��,�f蟰��p�	H��D��Pn�~?�Q�����#��Y��s�ϟ\h�9��4�d�<ͧ�?����3%9�`q��&"~� q���?����?�����NB}��'ib�']P�`P&T���[�.M��C��dH~}�HpӰ�m����b|�CQ<�l@A��3�r�*O�Hc!p�$)�����?ɥDh����ۧ^S��ݡ`���H�L�O0���O\���O��}ҙ'��[a��9G���FLڅ_���� ���tyR&|����Sh`tИ�ܮ4?�M�lV(,cƐ�	�Mۇ�iѬ7-K�:@�6M3?�fMˬ_[����?�fd�p@ �x���J�HF@}*H>�-O���O
���O����O� �I)���" O$_�D��s�<iQ���	����	R�s������'4`��4	��M�	07LӼ�����s�4 䉧���OM�4��H4x��'$�y�E+�^܃u��w�q6`�c�'^�%�ܗ'}:l��Q$5��p��ԛe������'tB�''2�'��S���OJ��r�L��&,ٙr�.�[F�رq$�$�ɦ9�?yER�\�	�D���!/V$gT�BW��H���Q�+�ɦE��?qiw�j����������&�
����X��M9@t�h�	��I�(��ğ���o�OD@a0�nw2�)p�Β{m�9�,O���]v}B�'��f��c��K�`΄"2B�٣���/���VN4���O�$�O��C�h�t�Ӻ;À� m᜸z�K�g�8�������'U�'��	՟���̟��ɀS
h�R4 ��$�,�[�,�$!�I�p�'2���?���?�ȟ��c�ˡ`�t���!�09�WX��©O$���O$�O�b L�"d�s�9I��P�J�F��� �� C�iO�ʓ��G��<%���D�/o�`YY�/�}��u��*�ڟ��	ڟd�I�T%?A�'w���W�JQ��0 ��C���.G��'j�Dr� �l��O�d�++)��š\����sx�D�O��84Er���Ӻ�d����D�?��֪@ 9�<=A����qU��(��Oʓ�?I���?����?������� ZT���	$:6Ё�npO���?���?qK~��]	��6O,MI�o1w�Ygl(>�"u���'^�1��+�i�Zd7-����c�WD�|I��W���X���O~��ƈ�?��>�D�<�'�?Y�G,xO��衧�:L|��$�K4�?y���?9�����_}B�'���'�f-�����q1�(*?��I`�$My}�'�R5�$�%j�]�"gE�O��T $��BL����1sChL~������ٟbG6O�@5^Y��pv�7Z�x�s�'&��'2�'��>�Γ�8�Flв!n0��0�O�#վ�ɹ��d�O��$�Ħ��?y�'r,����|�:�ŧ�	A��1k���?��]}���4M��������ń%{�����`BfΝ�T�h�'���{b�a*'�|Y��������I韼������#eĀfP�8q�
!�@�iqy�ƻ>q��?y����<�eV&s�ER�h��.��9X�M\?R��2�M��i)�O1��]ZÊO7���+2k�=e�+)��g�$t[��<qr�_$�����䓏�`�������Bq��Q�\�u��d�O���OH��O�˓2Z�I֟�&ѫ��q��Mۧ1����5e�ϟ�{ٴ��'�Z��?����y����k��Cg��D d�důI�re��4���&�
�ی�)dޅ;dU�o8�<���9]�XT@�OR���OV���O����O("|ZFN�P��pӉЄRW�yr��ßl�IϟਬO�1l��D��WΌ¤(]�2�0�� �+,�'O��'sB!��h�V<O���� 4�ک`UAX9t#�	�LǾi(uiD�
�~B�|rP���� ��ΟX�ėsL�K���G}�����؟x�	oy2ʠ>����?�����Q/l��a���܄V
���I9#`�	����O ��2��~r���^ �z�S>�p|AƠQ�Ly)E�����/O���
)�~��|��	Z �q�$cJ���V[�e��I؟��I�`�IG��`y��O��r6�O!c}RqLJ�u3�,(g�'w�	&�Mۉ�L�>�����M�u���@����P������?�f�ŧ�M+�'�I�G	���LyBk+Fc���C�
9	�c�

Q�bV���	ߟ��	ϟT�	ɟ��π D�B&�.yZ P��$����5��N�>����?!��䧦?�׾i��d׻m��p��0<vT3$���t�	؟�'�t��������^
�@m��<cڀD��7�ֹ[kА�����?Q���}�j�	L�	~y�'�R��z�HS�G�,<�x�B3g�-]R�'2��'<�ɽ��d�<��n��H�P�9%���@��>�����"�>�C�iH6�M���%��E�Paڰ��#X�wfɗ' B�k��Ϝ^Vș���T�ݟܙ0?O��1�gOɖ�R3" 	R�E�' �'z�'��>��x�0�ѯF[�d@T��?hx�����O6ʓq�F����Hd���ڞ\�|p�C
 !�.���O����O��Ō�6�+?1�@B�A�:����CAF�ye���#J^�g�>��sD#��<����?����?q��?�"��p���9t��$�Pc#�܇���A}��'��'��O	r�jx���
�k��Ae�3'���?�����Ş]�!�0��?,4*�zU��:d��I"g]�M��O�ق&���~��|�T�`�s�[ #&�D��5�Y�W�P��$���`��џD��Wy�c�>���-s�њ��ŭ� ��DKKRM��'��&�Cj}r�'��7O4�ච�)����7bu�4A��ox�f���!�f��M'Q>��;I��z�Z�xaƌis�M�j&�|���$�	˟$�	����U�O�|H5F��@�n,!��^�P�����?i�0)��vyr�p��b�p�� ԲXi$S(�v�D�2�9�$�O�d�O�����l�B�d��0��,Bkqv�y�B�0�X*ecJ/Y�(�$����4�\�D�O��$�7�"eI��]�GW~��m�7<�8���OH˓P��	�������Oٔ����ҍt�M�p��Ac8]{-O~��'B��'4ɧ���g���������!���'�����O�<t�F��������y��A�@�L��D����-QH>�jv셬G�.��I�����럈�	X�S~y"$�O2�zr�Mݦ+����k�8����'���,�Mk�R��>i��J l�!�j4�Z���IӇo��U���?��ʿ�M��Oİ� ��'��L|�,Li ���#��n�-!`˟t�'B�'
"�'g��'���5J3� �#W��Q�N
$gr��'���'^2���'$7mc��I3�Ϙi����$��@b/�O��0�$'��I��P7ͪ�,�2.YIմ5ZB�+�t��j�O�V�#�?�m7�Ĺ<�'�?����i\|�jDB��:!yf�D��?����?�����$[}��'��'�M�C�,5��I[c�%c�M���Wa}aj�<!oڌ��X}���)1\�6�3j�f��.OtĠ5ǝb�X��a�:���?�a�{�@������ ��A�F�=����O��d�O.�$�O��}Қ';��.v*F��D�	Jp좐-�Ο@�OH�09�&���$ ��lV}�����`��D�:�`���O�Ql���MSA�iU�Pֲio���O�И�h����,�/d4~�y�¶)>��7h��O˓�?���?y���?���R�f؂�L�.d|�c�nN�,\D�.O�P�'[��'�r���'�@ �4���7*ݒ�?r^�L�>�B�i@^7�@�)�||��eITHP�6 ��$���rd�yXf��'c�X���
Пt�e�|�S������ M�@<��([j| Q!�ϟ �	���	����Iwyb�>9�ӂ�ۢu�� �̈́g2�XGϯ�?�s�i��OH��'���'��$BF3�i�g	ƨ0<¬4NɀJ�~]H��iU�	8%e*��p����k�X;L]�o��W��s�b���t�	������8���hF��,I�1��0�5yOX�������?���?��W�\�'p�6:扉xB�XEᙀ!����� )e4�$�P��4X���O>R�2�i7��O8����#"������Z̤*t���t5��]lx�O˓�?����?���Hr,�1��S*?���[����=q���?y+OhT�'���'�?
@����zi����`��� �<Y�Q�$�I쟐'��O��e� _NH��AHr�>	b�ձn]޴���x�q�'��'>.%p��0[��4�0�����',��'	r�'��O�	��?Q��TG�r��b��hZ��Q7 ��(��џ���4��'1���?Q@e��3��hw([!h+�y�.���?y��hR�s�4���M�"�Ҏ�@�.~��HT�˟Y#f�y���?�*Od���O��$�Od�D�O��h�R`�3-��%�P�vO��J�8�OP�d�Od�=�9O�\n�<� ��/a��HD��7���A��ٟ��I@��y�S�P[�ls?�@��6>�B�:��Z�)IB�qqe���`�3/(#2$T\�	iy�O�"�U�]���`g�;'���1��M�"9B�'\��'A�!����O����OPi�sG��sA|�y�ηe-�`;��/����D�O��d.�D�(�n��˛�V
�:��S�t�����O$9���I��>T���@�f��A�<A �)(��w����3��؟H���p�IڟE��7OP�7��4��(�dڔ^��1�'�~ꓧ�$�ʦE�?���h�����xn�i�m�"��5���?���?-Z�P\nZV~��6"Q:��S���GJ�L�U��5��0��m'�(�'���'���'��'�� �tJ�3@ā��%I�ᚣ[���O����O\��(�9O��I7-�a�x$RpX� a�_}��'�r�|����"p렔s H�.>
R�PU�\Ը8�c�i���- (p���O�O��@�F�*�ĪY�P��Ή7x:<B��?����?���?	)O"e�'�R��4��c��\�T���Ǔ�2�q� ⟔r�O���O��	�Ns"�Q�l#$BҼ�b-H�HQN�pdDr���!%�E��m3�'�y��
9z�ّ��=���ŭ���?����?����?���?���	Ա{� D�T�Q�Y)j�[�n��F�b�'\Ҡ�>I-O<n�B�Ј��R�V�����87�&�P�	� �I�Jڡn�V~��-"��� ­$x8��E���0��&Qz?�K>I+O���OF���OPP�5&V�gM�h����&��	@��O���<�RW�$�Iʟ��I\�T�T�,?�����;Lv�������R}B�'���|J?�C���V�鱧�NK�90tLI�$rA`��m�T��'I�+�{?�K>�U�sX X�b�F����4�Z�?q��?���?�I~Z.O"T�	�Z`�y�,�3x�d��*)\5>��<iG�i1�Ov��'��e�(5D6!B7���}; AԺ+m��'@�m��i��	�M������ֆR�=	 ��nR)�C"*ZcB^���	۟��	�$��ɟ��O�R��m��2\���ۘk^8B�X�x���H�IS�s�4I�4�y�AJ5�00+�M��帰 �1�?a�����?���?1���M3�'h��vז���Bei�0�j�X��'�p�8 ��n?�O>-O�I�OV�B�	Z���5K �L�UG쑒7%�O6�D�OX�$�<�UP���������o~��-(<b��-�|��?	�S���	��<&���dD^)�jI	F�Sv���`�xy2m�/����i}�i>92��O�牺C5z�j��O�x8<i�e�)7���d�O��D�Ot��;ڧ�y�$'7�rBܻ�(	���я�?A�R�d�I��xR�4��'���DN�Z+аcG�\�vhXǍs���'���'z�1y��i�i��Y7��M�M�7��6n��rA ���N@�����O��D�O��$�ON���E8��p���H�R�:�o�"�"�	�L�	����2�\'�r�%G�t�bNv������ɂ��S�'S�Иc�F:��������0�Z&u�t$�'L	#rl����H�|2\�x ֯�*J:X����}��C��S����՟p�I����ly�ä>���X�r��p�9s"7e���@&�S�)۴��'���?����yҽVgH�a�ۇh��ȂD�!\��3ٴ��DD�D��'��O2�.F�"���$gS�Sʂ�!3a+��'h��'��'�"�S��v$ZDi�-#^�"N6OoJ���O��Q}rR�T�شƘ'؈c�B�6ImX=K��y�č(H>I��?	��O���ش��d���ZjȪ8�� �cjG����яQ*�?�cj,���<ͧ�?A���?È٤N��봣�1X��!���?i����$�H}��'���'1��K̆؃R%��Ü���� &��˓cP����M;�iK�O�'�~1󕠖8@����tF�`H�����W�w���M9?q��\>��䚲��\ƚmx�'D�;�6Uj����B��?����?����䧀���|�C�zpq�+ɾr zȂ�	�O>�D�O(�o�N�!��	ן�Y� U�&W�80t��+r��W��ڦ�ٴt��	ݴ����kW�4�'�ħRB�آujӄdo>�BK	x(.h��my"�'��'�R�'�2�?ՐBAT�д�VK$]�xb��YA}��'��'��O�s���	�d�U���_�;]���SH��lډ�M�7�x���K����O�!�F@�	Nt�[1�^�)CLȪ��'D��Ć�����"�|�V�������{� �K�ꊡ0Ux��e��������	XyR�>�-O���'jy��B�����퀈|L,�D�O�|n<�M{ҟxR��icX�3p��,��%��O0��4Vݰd��G	m�D��|
RG�O��*�'��立�r|�"k�y�T%j���?���?y��h����+#��홅!�-�4ԃ��;X����R}��'�2�uӂ��S�T��y	���!)T��ѬZ� y����?�ڴ}9��f�0_$�֔���a�5~����H���kF9<t��h�.S�~�D�3�|�^����������IΟ��fL� �VmJ�K�i^�Bp��~y�+�>����?������?Tb�0� e���0&+4P"�1x'�	��Mc��i�FO1�8�!�G�a�2Y����6]$!��٪l�1HƗ�\B�"
5T"2�f�Iuy�iV�/͎�Kō�)/m���L�B�'���'i��'��Ƀ����Ox����4wBѸ�͏3}?�5�bB�Ob�o�h��s�����M{ðiZ��]�J�0E�E�
�_r�hVn�,m���a��i�	�q)�p��O�q�:杮V�aiaa��Yd���蔵Bd�D�O����O,�$�O��6�'}ѐ�Y�ʒ3����@�̣y$x��؟�	�����O��̦9�<aF,�D-Av�:�詡 �c�꟨���<Q������'�<Q�+�w�����o�1O5��`�T�а�����4����O��$>� �1려 �/Ɉ݈��4�����'~�Y����O�ʓ�?y̟,5�'۔N��pZ!F�y(z�J�\�x
�OP��O�O�*����HN�٢��	�]���ZA�J&�&%n�I~��O�h�������Ä�9S��8���İ'q�����?���?������D�័W�_�s�q�6�] db8��t��O��$�Odnf�r���۟���kHL���
0��^Ǽ��`����	8 qB�o�_~Zwބ�ӟr�iz ͻĬǼrP���4/G�l%�fҹA�R���D��G�LS?{\Nm�E�¶fx�9�,[��Sd׳K����<3Xy��8Z`�a�r�U+K���C$��e�0����32ER�6'pJ���6FX����P!P��y*�A��X#\�u��$;�e)��l|�)uCǤM+���CGD���jC��D,�z��*/'L���+�(��u��dh|�{ӇTT����\�P��Gվ!Qa fH���P�xP]�R�S|���و~���+éo4�iiC[h�K�M�O��Z���� �u�A�j��[(ħs≩�A^?8P
t-%V��c#�?V����K>x�}���2��*[�n���oҖgd���l6u�R�m�=!���d��D�f�� O�>ls#l՘{\�i�$n<a2B��hn+��肄eF�;��L�1x[+�޸"��D���L�z��Za�m�
̂Z#t�7 �I�H 0�U�'�����L�zJ˧m���c�4�?!��?-�M��T���'��1O��C]&�����1%��!���d�(p�1O��d�Or��7Fݜ,	�G(B/<��QJO?MJ���O���y}Z��I}�^�RB��r���2&�?[����'t	��|�'��'��6���t�����
�&Ɋ�\�D�O}�W���IX�	ҟ��	�3�D����FDX�Q ڢE�tq ���@�'���'����1�r�s��O� ��Yh3/r>�PӅ�'��'r�|�'s�MԻz ��R�f��l��.�Ng@����M��I�����ß�'?=�����P5MG��+w�Y���IA�_ ?q���Of�O��$�O��,�	�GGT��B�Ү�/r{���O
�Ī<q�!,��ԟ ����(�CהF78p�D+�A� ��{y��'A��'�hx�U>����[�<Ř��	Y�E��?�+OD�d�O����O��D�O�ʓ<��� �i��cQ֜����<Q��Y���?1��#4 \���� �NHSF�:3�ab�k	(�?�w�6�'��'�"��>i-OBZ%��@EB0�1�0&y �	�!�O�c@��n���?q�ny�D�;�C++�&��C7@�f�'Cr�' ��>1*O�dm�$�Ue��C�`�S��3H�����-���8�%�8�	ן���6x�A1�@:w��z�ۡQ��U�Iԟ��I���<I���(����eD#v8����C���Z*O�9��)�O˓�?	���?̟����+�\L`���MK�K1�'v�ꓽ�D�O��O��d�O��3�� W������<wD��O��O$���Oh�+�I��?��6I��e�C�\�j%8�0��O���?�M>����?a"/��y�.�Z"���+�ti+��>��D�O���O>��|m'>�peR�� IB����,�BHb)��$�Id��ey�O?�Y�X ��@���-���* D�O����O��?A!����'���
Zh��ʰ�_�xrXh��Q�*��'�	����q�s��)�E!A��#E"�:
�b9�c����'�ronӤ˧�?A��p�I�B��/��'N+��1�M�O���?�����'��0���P�\�L���ȓ�Ӧ!�4U�,O����O����O�d�<�O��9#�]�oY������KFxic�X���qa0�S�OFZ�ue�0-ؐ��V����< p�'g"�'��'��)Z�O4 #�@�"�z<@@ʍo�Dzw�܍�O��?��	�<����2�0!���t�N�r��@̟��Iݟ̗'+�M��w���Z�R�A5 ���m�5IL>I��A̓�?�.O牉zP��#�\D5�I�SÁB����˓�?�����'B7Oj�y�ö`���͆�?�A���'�đ��O��d�O�$,�	��?	څ�e�8����Sgtp@p-�<���?�I>�(O���O�����=/��"���pi0��0���O\����|���K��9Y�'��iPr����܂[�y����'�P�<)��>}��~�kg�D9Q�2%{����?�����ĵ<�/�p���O���|��P��$�;j��!'��$x/<�O�ĵ<!�*�l�'{.y���[�ZM���i�<��y��'y�	��ߴ����O���|y2�wR�a�A�3X��&�?q/O��d�O��Ȓ���%�͙z��d��E�� )��&�O���֦m�I����˟��J<������cn�)G��!�n��Iɟ��	۟h$��g~�������|�~T��@��7��'J��'H�P����U�
^v�4"�����1��!.��Q���<�I�OJ��O���`�� g(c6��'13bd��O��$�ONq&��'��nX}h4f�-w
��u�/ԡ�K>�������O����O,�f���&Cʼd���!��̅col`�� �ē�?�������D � �e�*KN��	��ܘ�"�'~2V��I柘��X��r� �������na�9:GMRy��'NҘ|�_������7eшe�:dc�i�s6�@�I
{y2�'m��'��O���'�?q�ܿR�@�h��  ,�*h
��0�?!����O����O�@ѳ���S�6��a��HL���bׁ<�*���㟀�IQyB�'0dꧦ?1��?A��T�{=t�puK�!n�T�Wm�4����O����O�9x�?OT��<�O��p	����9� -V
E�ԩ���d�Oj�nZ러�����I���������D�[:	� \�gl]�es�d�O������Iry2�	�	�DI ���p��u
��T����'�\7��O`���Ox��Hk}�S�t�\}d��J�gFF�z!
�����Ehe���	oy��i�O*h�pO�]�������r�� AA榥��ݟ��I���ӬO���?	�'	�aB�*���(s)ě@b����?)OD��E�?���O����OF�b�*Ɇ~�����P�T�s��O����O���'�������'��.��,S|qYR��Ql"��WH�4��I�\R�	}y��'����9��r��,]�a�`��".�>�*O��$�<����?A�Nh�����E8!Q�����%5��D3����<*O����O��$(����?�� `57n�!$�H�:��XU��O�˓�?!+O����OL�����DR�#�nUR�-+i)ޡZ`Z�89��'���'2�S��S0��	f��T�[�2�~%K�
� o����WD�O|���<����?��lAHe�O!��P&C������R^�\����Ϸ�?���?�-O8���k�T�'���'�Xx!K<��l��D�=�T�[���	ҟ(�Ɏ��Ix�	�|*Q�F��B�xP�1� ���͞�Д'/��o� ���OF���Od��'4�聴#h���C$�Eo�s��':R�'2���'��S��|�*Xc65(�	�gSzP�WٟX�I<�M;��?!��?IPX��'W⠚A���7�����g#���s��'�֍+��� ���H�@F�1Bሴ�����Y�č��4�?���?����	Ny"�'��Id� �̜1�hdS ��	��V����*,j�'?��	ݟ<�I��X"���Q)�0a-G?���	ɟH����ē�?��������&�0@^4t#�Ʌ��8�)O<��T��Od���O�'H��:��tK�3f� 8���ē�?y�����?q�TnE��-�=�`��M86�ҹ��ꅦ�?�)O���O�&���?ur&�*Ib�9��J3�����!�<���?YK>����?���_}"�ɛqҲ�Km��U�T���Xy�'k�'a�O�P�ܜ�I�97��u�+E�C������O��d>���O���D�P��:?�4�ͫpZ8E[G�ҭc����"���L�I��ؖ'�rD<���O$��W�V��0��.�>?N^��s�=Q�ʓO\���Ol8CGk�OƒO��S0$I��q���3�e���p3����<��Aۛv]>��	���.O�% �N�!8�#��EtG�d9t�'S�'#^��'��';1���Reƭ<pJ�X�MW7u-l����'P��t����O2��O�&�p�Ih�b���lY�Ge���`�<`$�I>�����a��O���?ـ@Ҿa�<��ۣ>�8�K�jއ`���'Q��'��!��O�e�ܣ@k$��@!��e�Z�٥&�O<�O�xaA3O4˓�?����yG抂�����* �����I�?���?i5�x��'�|ҁ߸3_ݲ��,e��z�+.
�	�:5��Ty��'Rr�'R��X�T��%N>2Ű�)�!)z��D
o��?J>A���?��'T�Zz-�Ո
�����Gh�(LC������O��d�Oz��� ��5)���C/�Dj؄�VC��7����?i���䓖?a��6�Y�ljN���-SLF]�'m �ue�`�.O@���O��d:��Bt�S�
-B�H�D��-!t�c�)Ҝh#��I՟�$��	՟첥x���'��l�wC���ؐ��%� �Ź��?�����O.�$>�	̟�CTa�� 9��M̍gX��S(XZ�͟��	�5���Ip�	�|Z�BV5I�֨�"��bq���d�՟P�')2 j��ʧ�?I��uS�/�bĚCEA*'��� D�[�>�ʓ���O���OiBI1���
m)� �"蔄j1���?��ilB�'�2�'�RO�I��f:@����D+5Ϛ��䜟/�(ʓ�?������'� l+�I%BU���D&�:"��q�'�U�D����p�	Uy�'��A�J��L;��ش]/0�:�&he��S��D3�i�O����Of	P����
��݋���.Mb����g�O����O��'��O-Ҝ���ǒ�*�C�j����px���䒶jD����I՟P�	�|�$Y���<r�m�Y���jS�̔'X��'�2�|��'���u��2��JJ�Xѥ�,1��"����d�O�D�Or�d�|��O���نC�PzH�vEN�_�
`����?��?yM>�����A��Z�H� ��A�vH��3�&!+w��<����?Q���'5���ԟ�) �C��@��1`(1b�/�ş��	ğ�?)d�!���� �U�g�Ѭ4Lh�q�߼;�����'hR�'��'B�'M2�'��'F:5�T$Л] e���V.w�U1q�|��'��.?��"<)��Qd��󶢄��} Ek�;� ��O9i&Vt80@_X����!�j�������u��U�4�L�]0q:d�Cŀʐ�z k�	Q��^�O>�w��l��?!���?����]�>�$��d؂+�vl×+<i^���?Y�M����e����2O�d8���H��ܹZ�Y�1��|��D��p�ld���i�، ��*],��NEO��e�3;�D�@B͑D���P2�U�(lS���5�L)��T�b�<Y����ss �A�B�fȶO�v)��j��\%mk�h�w�ژY�ؑ04���H�r���i��]9�"�gò����T'B�Lx��5���v�V����aÛy�!$�[�B% 1�Y*�9�	7mJ�DG98�U�Ҧ�$b��+��<XX�#s撎@5�嘑E�b�0"#g��!�@�6W�oZȟ m(��8������AC��"+2�����S3�r��1�R/�*����đsk�D�iZ7o�	KhܨYb_�dK�o�N��Cb�
M>TD���_P�,��d�L�y	��ӯT.��$$sE��'��)�ɴ>9ņ͌Z2b@�ƯM� ���Ac��l�<I��
����aJ).& -J 'i�'�R�~Z�ƞ��@�#H&Y;.�Ɐk?!��?�7nЋ|E���'��'��ۦ�S�'�*��qq/\�Wj8p�JЯE��S��+ ����g��^j�o	Fɪśd�F](�P��+�y}R�ӹOZh:B�.����4�,0�nއZ����#�ү@����'������?���w
�q�b�,�b���c�zU�'>�A`���nZ��鏽[22A��'�#=�Of�ɳS~�j���@z8 ���?�)�ǉ\��M����?q���D�Oz��u>�����9{���j\����ՉQ9
zj���!�!B�gx�\��ڼל`Ir���J^t2�\�m96�ht/��4o]�w��~x��pt/`�ya�9���&�� 570��Qܟ(D{��I�NLY����1>�đc �[�C��Q��h"L�8(-�ŋR���d�'��듓���W��Mm�՟0�I�U���M+?�~�k� �-w���2��S���$�O����O���l�O��O� ��X��P�`a�+s�`U�B���O�y��^8�Ȑp&
q����"YҎQ� G'X���T�N��O����'��C/�$
�KuhEK�)�@� b�n�傊�OL�$!�)�'�@l٧� !R EK�C��!��)�O>��޴�M��J�E��M+��*	�Ek1�ġJ���y�,�;ش�?�����'�?q�4}^)��Gv�����1'X�����'j��O�D�r�rs�F^���F�
M�O|��9��4C6�Î?$��.^}�!T�^k�lQ���MX<���ϋ�y&~���J��Plج�6=A�oV7|� ��E�w@�]J�U��˷`�O��oڏ�M[����'�rڴm�ti .@�"�xIg��^M���F�'�r�'Ra{���?<TL���ŅФ�	�Γ:�OD l�=�M{����u���Ҡ*��:��YW �3U�^��g؟@{Uȝ(�� ��(gB,m�d�3D�pJ��� 5R��w ��A0d�$s&�5*�eX�~��]�tȋ�l&v�,�b�� �C�IV`<@�)ǭS��|q�ɋ��B�QP��K�8X�i��D"�B䉤#b�N�̀�4b�)��B�	�(��)�`ħ_��a-��h�B�	)M߂ it��UK���OV�O�fB��-��,��Q�Sd�ʛ`BB�I�R����g�[x���w�N�h�(B�	�[�^�䁉�x�j�aEO.d�@B�I�~ihF�Wk�*�:&��RB�I����	�n�G��Ą�1H�TB�	�:������ �]^��f(�3<�*B�ɷB�TRb��QKd��LBdB��h��aҪV'���C͠#7 B�I�z�����0-��C��&n�^B�ɖ[t��%�l�Uȕ��#}b�B�I}n8��A(�O6��(�K����B�I�}�Z�wVQ�D� �\�<7�B䉸	=�/G	ތ��(DE�C�	�6`]�4�O�Lx �g!0�C�>�b�2B!ͥAA6̊��R� LC䉽[T��W��R�:�j��� m<C�	�E LRR�\
5���U�ObB�B�	���\�V��=��|k1�-D�� ����K� �����
��L0l`�c"O<�ꓛL�V�l˚� #T�:�"OɁ��ڞ2�pĻp\�\�N	"OP���}�"Lߨ	J 1��"Oε��%4�4h���v5Z��'̸��ubN)O�U��Z)���'��I�$��]1`J��ͮ>���
�'������)�0pȤ��Lp�p8�'�Z���i�4T8��sL�>>��9�'+��rHP�|"����
 �� 	�'��!��R�l_tU0��Ӵ3�E�	�',.i�A�j,�fȶhH�}

�'����"@ؗ3��l���?֊���'94s�������9�lƹv�\�'�*k�=0Z$���ǐi<|��'���+�%ۊ�*S�4�.� �']X	��*l�	��/�#}��5Y�'vP��Ӏ?����[-t����'�iF�ϝp&@��n�P}��'C���*0}�L��HOf�X@Y�'��$�ۺP]�}i�.A"j�c�'Y�$Cj��V�JyK��={��;�'l݈ѮԊb1�g���jiT��'�LM��c�
N�M2$���(�#�'��x����h��S-և�N�Z�'�,�����2Vqâ�"����
�'c U�VD [BtB���5 2��	�'��X2 �<x `�b��@=v�����';�\3���^>�X��À0����'B
́�b�`<�r3n�=dʺ	�'KD)��C`>0)@uE��d��Tq�'��P6��v@Pm�mҥd��[
�'�� �Y&{Ȯ�4J�		E�D�	�'3�e�G����؀��Rm��@	�'��%�Ĉ$Z�����`�2U�z a	�'�"��@Aҍ2ۜ���S�6�	�'�h0p�M�]H��A��1Rv�i	�'�\�F�F�+�Ar����l��#/D�T���� C�~���V? 1��-D��3R�<X��s���0q��ɇ�*D����)C�e� L��cU;E��tR5 <D����~%�C�!�i#��B�<D�xS��n��Œ�`�~���b�.�ɇ~���j��'p���%GjE@d'�y�V�p����N��2�\�w�M�.<�E;$���8�%�Oƙ[��ьx��q�q�>�a�5�sIv5�Q�P94�Hӷ�~����+;�1	���� ���Cr�<Q���!k������:�҈��K���&��<�6�󎍹�0�F�t��O��P[f��7�`�S��֬_t1Ob�C֍V,�p<�F� �D�Fi���VJ�&,�"`�op�ɖ
�b����*�ݕϘ'v��$�LT������9l \Sp�EVF��T�'*�H�
Ƞ3���d�4*��()�b$?�� �dF�Y����R?���+H,#rn��h��Y�#�J��䟘��e	���^tC��V�Sӎ "鉑	H\Ɋk�~%����(hE�I�-Iz4�[�F�5n��-@7&e||x`��C<o~L��^ q�`xr�Gǆz6�s�f'ʧ�����"/�`��ߒde|� H�Q},0�2m��8�		&W>	�]	��ts��O�J���L	(�(��4'��z�V���%�kA��hsY/Vb͸��0M�����7^t\�K�x� \P(��:i�'�Kt���	�V�&�!ڟ�6�ˁ|�p �hҞ�C `��YA8�kd��!y/�(�E�˳]�p����B�C�V����Eg��])�[��t���a���H�[�[�M
&i��}	�Hq�D`3ԫB�N�$� q% ���4E�2�����޽EN�v�j�$&3�RL(���ԡK�.	�q�v�S�&Ҳ�TH��v�L��@�����$Y?8d�ɱ��Gn�� �^�iE���s��|D��8���?-8���*@��!B��ޣ.��Zs�U�A�j�"� e�	
0�ڭ0�T�9���*A��= fߠ)���Ͽ��

>dT.(�C����04��Hn���#�E�2?.bHZ�탒m�.��O���?�5���2(�8�� d�����\P(B �b��� w|�O3.�b��"
o��#�B�]V,� �1	�02��A2�1�f`hRgB�(sC�_'g�">9��J��q��S�>*|qÔ�Y#.}�����I�+t�#��6O��9⢇M/n9�8�"�Ϩ8$b��y��a�ۏ&	���s��[.�94m'&�`�"&�<j�i��ێ ڦʒ[9r!�	��Д!Amɣ��-� ��!z���@ԌA�-�LAɀ��#������E���-��9�0ܟv���n����Q�;�"|	2�V>KB4[t�X�W8`6m�.E���AgH�b� ��j��r�m���]/y��`�O9d��S�B�_���cg�
z@2t����/-\j,�]��sw�Y
{B6|���O�z�e������ 'I~���Beu2����D��Z�։,�6PIǓ�8�D�]3D�����
Q�ɕ�5&,��	��̒``T3�h�juA����>aU!R���p��,ܖ����/xT\�"u��P�����;��ܲGŭU�2��'<�dӳK�\�'��L�&�ORz�)��%9D01���ߖH��ʏ� �֝�$�	%�A�TmVfB�H��U�,u���In�q.OT��t���q$*������(Y� Q?|�E[��	9i�������cLZ*.�R�� pz��i�h�_���,'
�ũ�#ڲ#�L4�$��(7�0�T�L�/=�%����0&����Ɏ�9��@���@�I�Nr.�A�e
�(<jq��`bA��Þ�M��O��6�� Q��&:��u��PF!�d�1fa�0���
)z.%If����IFXP�#��s�i>M�Si�2Zu�	"Әcq� (9��SBO�e9�C��!6�hRe,�W��$�%�ٿ
ۈ�O�,�u'��ي��$Ư���˲��Č��K��!�F��������`�����+)΢��K��PxR��q�a�֋��%�V�O �y���'u�1��ݿ ��pY�hT�y�A,p�W�ΐ�D�y�h/�y��2��4����P8��H��y�'�qId�Z!A�4t8h[������W
@����a;\O�1�tKY+{}h�B�ş�ȉ[g�'~N�
w�ݴo8�z�$_<=ڴ��@8Eǂ�!����<��X�1�]*6#�:lΨ�1��y�'����\0{(n0�D�ɏ�Rz$u�b/�!�f���
P�!���%KR���)��t���'j�9j2dD�.�,�Ҡi�<E��'��dƐ�sY��#�P!h�,��'�`"�hF�.8�֑g�L��yb �c�X���+ܘs��y��S&R���ϛ2�"��#J?�0>E�w_�3U�S(S]||�e�W�c2�z�Ň�cf&�#�'�����"̠lA`$L5*���a���8�6J�c��F!��?���i�C;`<ң�d��PA!d6D�8	([.2�z9*��X�/�p8������r���v��������d��/ ���U50�D� �CB�:�!�$ނa��������!2$���6���ȿ�&�1�ꚣAp��$@Wm�l���T"�}H�H�Ho�|�a�OR*�!P��:ר����1�r��D�3��̠S�Z�O�~�"~���0�7��3h(�@���eDzbl�@bԋ���4������Z۸�å �#q&�dsK�-���;�O�A��ͯk�&� �Bæ]��q��'�X|���4-g<9�I�Y�,,3#�ȁf���PY&J�y҉ݮl���j�y�^��%�H���'2b�qr��%r��mF�$�(t�`\�P(� ό�"&��&�y�� /F<�z�e�1��m�%H�A��0����(UZ�s��>�U�P���/d��Xs��M�9aPՅ�@%aD,�Mn�U(&@Z;���m�(&��՘w�9��{��
O�*�Y1J�9�ָq��ѕ��=)w@[��!(^���G�P�@"���Uڸ�5mR�dD!�d��9�d��U%B5;p���F�O
�Z���$�h��	�\]�ШDl�5z�K��A��!�ӞF�v(s�]�5�lP��ҒK�2�Q�33���'�6#}�'Rvb���2��:0o�
+�����'�e D6ܨQ��P�%Q�3��BB�uۗ��0>���N�Ai*�i��5A#�pb&��L�
Ɠ30���F�D��%�F1e�`�f%1)!��(���1c�I���*uˉ!/��ZL�(D'i���i�
DȬʣ��6lQb��5�O�M�E�ē֥�?��9"O�[P �b�12���m�� ��R#ڸ�T斲Q���Ex"J�?9�:X�q��;G�t��F��u���]�6��+E"O� zp#�� Z��](�-o���6A'�$���݇Q���S��yr��f����Ò:X&��ړAÆ�y��)�~X�r�ɒ}t"���yBMG�*{�	瀦@S�y��U�1��MjD
Ғ,`�3t�$�0>	P���8̀TJ�(�|���V�VA�U�T����Ρ�
�'q\*���K�R)��ߚKbV����+{	��H��
�k�|�?)���O i`����1-:]���?D��s� ��Vm�U�S.u��p����<��hp*T$Z#6햧����?�iR�Q��۵F4qW!�ۜ���e
eqh�H�
Y;:��$[W�hfg�f����d��/�r�+vNʃTr���Sf�|�CΎMPN����˽$������3|�V(�[��u�C�*D�X���	H@d�q��D��굉+�M^��q�D�$�(�z0��y���D(�&��"O��@2
J�H��$T~T�v"O�A`M��H��s��	����3"OPMO���H�qOD-a��t˓"O��sDˏ�ey`� �.��,6}�"O��!��+�<�bNB�l�����"O&�x�f���nyqs]((�6��D"O~���[6�D�iv+_�P�VE��"Ol�*�!�0٥��-R,���hژ�yd�/	�r��WJؓ��M��ybL�"1��"�!�Uq:������yrኗ1���h�"8�|D�����yR�N~l�l��0O�ʝv���y��(٤��r)֠<=bՒ����y��X��V-s��1{p��τ��y¨�}�p e�%"&�	� ����y2�B�~TRN[g^ )ӊQ5�yb�N�&8�P²�NQ_h���L���y"�H3DV�	On �A�S'�VB�ɶ#��-ȱ@$c�X�
&ή\�^B��.U�T��nd:�@De��B�	�{�X�
p+�d^�-8�L�0�C��*jP\�����s��!b���\pHC䉙QC�T1_�|Ǹ5qd�HP�|B�ɸ7qJu!�BU�1�u�]'&"B�I�t�Mi3H�8tUrh�6B�i���ȢD(��eH*ba�l"D��P@�C�0춴�"��z�d� h$D� 3qE�nò��'�,%�&M�C&%D�<�
Շ/�b�8�Dа`�4��� D�X���It��:�͎&I{:��6EA�>����Z+t��T��ɱ^ٰ��k�K����ޣk'�C�ɤ��#���pqH�:��C�	�"(�w�P5@}
1��),�C䉇�:�3So��;U	����<C�	<H��| &�(
UӪؙ\oC�(b��-3���;��f)BC�	9k�vU��D�(��˵���6�C�	�˼��qC�.0zzBő�2\&C䉂EU�(��Cj��)�f�o�B�I�c��E:Q���,��x����$�B�	�N�����	�2#r����ċ+�jC��	X�~JHѡ����W��<C剟/�\�1�	�b�f�����d�!��Ùe�8��H�q�e0��W6�!�D�!p!�EI�X6DE
%0�f)�!��t��`ꕁN�Щ� �x#!��۩{�0�d;�t�	��R�7�!��H-d�;q�ɼ0R����h�w�!��	Y�t�� �����R4���!��ʤ}�d<���'	�z�!��  ���$3m�*	4uД�"O�:2` �/�9��cҴS�B=�W"O �pĭB`���r�Ѱ����"O���+(�JTd�"��:U"O��Ѷ�ȹ`Or�	 l��o)`m� "O�\�'m_�4�DM�u����0��"Ox���_�=PȲB�	��s"O~��&��9'5:T�'xw�<(1"O��c�=[��̳�̢Il�5�"Ob�����68�eSd�4S6"OLܑ�M�5!�@R�f��"O�}�7�-���j�:=�a�"O�l��JZ�bEu�K�3�  "OL\�c�;R�@��סˆp���;�"Ox\hU��w�����g��\���%"O�hJ�GO�����E��dKa"O���� Q���̇0n��H@"OD��C6r����O�5a��|b�"OJ�) ��p�J�a�-P�f=��"O�\���Z:Hq���Ii��"O�('i��L����8@D҆"O�T�'�:�V��5*9J� dV"ON$�t K6�ѡ#	�Y�4,�"O4�p���JL��kN�S���2"Ox=Z�*ȡc��)J	7�u��"O4X��D�	��kp�H`.1�"O�`)��*Z�����+&鼙 $"O��Ԅ�
a6���G�C1qք���"O���3	��X��)(˅�V�(E"O$�&����#���y�F�	�"O��T�=��\�R�.e���e"O�9��J���]�`�J�9��H�"O�%��mt�f�(`e��4�5{g"O��Rf��J�  ��%�i��"O!W%)rm�M��M� =�XҶ�D�$5�x���1]w���ǭ�;=��I"l�\C��3Y�\Kw��lt|����X����շpO��d��i����nŒud�IcI��1�ax2��s#���=i3�m�ԅ{�]]��fcBj�<��茅]j����FW�H�9s�RL~�ڏ6����=E�$Ň{�"�nؽpw���߸"!�$]#3~�(C� Q���7F�{WqO��[�ƈ8� ��'Ⱦ"J(	�AߎV��醩)D�Ђ����cKW*3�|D�U�2D��" $:A杻%(�%���%D��c�$�u��*.Vz��� �"D�誥/��a�6�@w��`߀���*D������@x�Bf�:^Ff)�E#D��@A\!_E����H��Iv)7D�h��	ZO�"@[�J+!��
A6D�,K �	P�p!�tj6��5��G.D�����T��tx�t-C�z\�ʤ�6D�h��GO-A���&�®f�T�PwO7D��Z�NM�7}|t��%��J�<�O�,B%k�H�S�T)u`ԩi�,�bg�6d���>0h�>Q3��#{��03��->G�Z7IX*5�:�����Oz�9�Üu���Bs��p��=k��I�/}p��h, q5���) ���;p�4�`Ӑ���]N��[���CWl`��M�����I����1�o��� t�W��6���f ��/@��'��5�8/D��B��F�Xs����4�A�5��+�
A*��
(ZE6�ȓ6�L֌�0�ɤ�ڮ:��Ğ����@6-����RmY�Bצi�4P�ʢ�wݺ�'q��h�`�F�W6��)��İwP�u��s^@*�MA�u1M��Q�J%b` �2B4Bpu�V#������O�(!@+!�lt2џ02�y��۸v�����؉4�@Q��	�(OQ3��Èc������tn@S��%��i� J�YF)��n�����M�*2~�֪�%	��ܪ^t�&�'s�@K�
�%(��*��_�b���4'�Dm Y�T��B8~(�P,,�AI��h�(��O�"����0/yӴT+��� ��8Q�㕧�x�"O�`r�C�n'�-ڢĊ�g�����\�t&ֲ
,�+r����ap�K�Ŧ�X�I�%1�N� vIk�U��H�l�F�ʚ/4՘�<�O�i�7�j��H	�M_� �:'*�)��Ç͗�0xP��	��?�Ve <X|X�U8?��9!"{�~��`E�9�A��-ڀL<ғx ��7��r�H��4i 4eP,0��u/C�G�49���f��TKǰhw2�z�FӰ�}�eF�5�y�ˋ&>4
�Z ��A���ǀE��?�E��e �b�G���嚳Û~�
�X��6��
ÈU��y2���D� ����)0�a�f-Ӆ�yH��B�zjS(�.�y8 ��$A$)(���Ţ9థ��#B\M�@���?iU$�#N�zx;&���y�f��"���!�c�A�vt�`�ʎ��>�d�Ҿ\�f�(TEح��@%K�K��\�)nݻ��s����G���RI��{�8�D-;�Id:M�'��%���&�7'\">駌T�i;�� ��ű8���~��u %b�	�ʐH�1�Iڗ�W�-���4q��� �����չ.�F�{��V��p̓	X��T`L���TX�� @���ənEF�y��F�<ͧ�,}���6P�*I��0K,�Ї��@ ����k��XU��/y�yq�� R�x���'����O��z�@p��S�7��W�g��t��T��`�1��~bHܐ�(��Ƒ5�YW���BQlPP�J^PynM�6
D�EI
9�J��ul�!�(O�RN�nq�����@}00�I4x5���B�_(_� �[���=&�e�&]�]���b��.F�d��	��Ҵ��m	j6a}����%.�Q�ڼG�>E�h�2��DT5*s����}KT-�$hY�O<Tu��i�J�.�r�g������/�*�!�D���3&Q�1|��v(����!��M x�TYGϹ<�}��@2C���	z��6씈a�����L^�G�4B�"aZZѳ�@��v��z�ȝ�'��`�O졹q"�%�H@� D[K�'|h��Я|�҅� ݎQy���ד4��I�4}��rF�Y b���dkLP�X"�K�c�"B�Y؟��o�;]��\+�o��zD����1�}���qܕ"{c>ݳ�AZ���*]'���0D��)	 �Zԏ�����!�j�>y�Ă>4��<E���t#���@Gy*H���.�y«�6<K���@D8qq�F�4�yB�(u΅X��(!�YYш=�y"BXw�]�3�̚i��lr�i���ybFDOD��ΟY�6�1�$��0?��7*�X���G�,�"@�&-PF�U`�G�<iFA�=i"�["��"p�`1���C�'�8� 'L����X��G!� u"�G�1*e���"O��Q�!�|U°�Q92cd��02O�P��V'1O?-��K�4d�r��o�� $�>D��0w�\9u~l����T��8��??�L��;�ĵ��I-P�Qɷd�p�B]���8����DD�z�@��sIVM� ��:������8)�!���]�y��eJ<���pF���m�|C���88�"|2U���U�0đ��G"S���G�T�<	vaC���D�'������d�_T�<1B�5!�4�pI�f\�)b-�d�<���V$@�=���ԗ,rpH�{�<��
�e��l�"c:�Sd�y�<��AJ3v,zBjإ4-�$�U��r�<��lX���:9ۼˤ��D�<ir �f�റf͂�D�����B�<9`���z! 9-I��-�`(�<w�C�	�{X��F�ۑ;�deA��ڱ� B��2�س�B:R���C턧p�C�I�R�!���Q�NO�	(���%4b����ҡ~����<�â��[�Y��!��p��W�<Q��-��I����1yh8q��U��k��0�}���OR@f�m���Q&~Ѩ�e���y���
[��\�S�-`%1�i9�>	���r�f� jS�"�����Òфē/� � ���C,f��@�N�z��D9XT��S�? �M�Q���fT�% Ă��H� ���'\�@�{���F�����	Q	ܠ�#
��yr ь!�(�5��#M,��zq!�(�ygMS�8�2��q��%� �F��y"LQ.Q!���aU q�`'��yr�F�	,h%��Q�<eb�A��y�	�Bը�X�'��8N�H �@3�yr-�2R�2����H�|�����>A��.ƾ��ꖅo��������D�H�B�G[�!�AY]�숵%R�0����䔖P����U���*Jf䚒��I�o����C*sZܵ�J�!�$��}�V�� ��o^�s��J��6���1W��i��sӲ�2̘Mw�A�ң@6,A�5q�"O���T�ַ:����,���T����� �0E���' �YF� `�9ab�:Pa�I	�Ti�iY���7d�z����,��ić�<���aO�I���'C젚��:%����D"O������8���E(����	�"O����@**m��FO�i�P� "OB�uȋ1��(uD_�'r��s"O�@h�Y8��8��;cTVt��"O�,�h�F�0Y�AϹkRāS�"Oƀ���Bw ��w��|=���"O���w�J�d%#%�l!:հ�"OX���5hS�l��/�$"��#""O�k�I�|������^����0"O1�t���1CM(���6"OV ���S�X�!Bat�� ��"O䉩u�:J�����ܠ��}�F"Of���m�8����U�5�X�"O$��B�h�n�eω�?<��a"O�y)q	��aN���^�>4���"O�`f)��Y��QA!@C�t��"O�fؒ�)7� ���	A"O�lS���54�^�;�-,t]Lp �"O��0��< ��1��>f���G"O�����1z.�[�ץ^>�"ORKfG��;�@T�$-(6S�ai�"O�Jdk��")����"!UXp#�"O`y�@
X��E;C�! ����"O�!�o	�S��谁	S�2�lb$"O���c"iI�)�v�
�A&���"O��F���U�H�
iX�BW"O8�#Bϑ��8]�6[c���;a"O6L�c����B�,�=M� �6"O�ѳ&]6{�BM�@	<(̩"O�,�"@գg�8�SkZ�p����"O��A6�I05R�!��LI�����"O��z!j��.�tՏ4#�1"O�`���6`] �z@퀥x�ڹ��"Ob�Ѥ�?�����M6D�f��&"OBdBqLӜ��J�#١v�6���"O�����F�����L g�Θw"O�a�jXh�>��d˫����"O8U!M�^�hw$R1	K$,�1"O�`�2�X�|,\�سa��^\��P"O�=ڇg͹Z��] �>"J$���"O5P���+�j����.�e�T"O�t��ϐ�nŋ*����"O��sfхo���3�Y�;�X�3�"OJ`�%	��E>4�a��V���!�"O�*���2蜹A�LF'�DA(�"Od��ƇH�Ik`K��$_|�Ku"O�X��sz~T�U��'R���p"O� V5�u@�M,�i�@�B��]��"O���A�87�ܓF��_�����"O��Z���Kob�bת�f���U"OzXj���g�D�D�' ^�m9 "Oژ�4C�� c�5�"�'� �j�*O^dZ�lD�q_��sA�nN�}0�'F�# ��?}L�dR`El���'8��@��z�Y�&jD�W4����'|�=)�KB�)fV�㖭��Ob�tr�'�z����K�ς R��ED����1hę��A�f�C��87���ȓ8Q����x� \�����}�hX�����cJ�mN8IG�ⰹ����H���+#5$5��� %_����|D$�����/��(%�X6ڊ��ȓE\���D�H�K�`Pt;�8��% p��e[Zf���k�)�ȓ%��p��ŀ9H�1$�9%P����r��A�Ţ�^�HRFS6h
h|�ȓ}����@l�Y:|� U���{>Ԅ��4��I�O 	�T����_6��ȓ�NeH����r\6��gY�A��@��i�DH5GL�H�L����(!����>d��6��X�# ';��ȓ
LMzDa[*��D�ujEl(��ȓ.M�A������0���Z]�8�ȓh,��@���� ]ZR%b�����w�\��\�S���YPn�?�T|�ȓ�P�ӕh��k̊|����5m��ȓW�:q�(H>���J�_�DY���54(������:���C֎��|�=�U
(�T�0NB�h"���:�4#�M.>�0R7�ͮ+]��'|�k��׫A�z��p����%�ȓ<%��t�^+�,5QD(��Ꝇ�.b�0@��R���B^��
��ȓt�P9����4Fx��q(��:y�ȓ���bUf/p�� �a�n���� W�
Q0>]`e�ф�d���H�9%X��C��Z��نȓB>N���`K�H��H�1ˉ3CPԆ�[~�!4�.������OnU�ȓ>�P��$�1W�FS-N�z�(	�ȓ,V�̃�Iո��颴���M����Ov��"�� /\Z��ݫ3-�ȓ4,:��1#V�7`��H0��'��̱���^D��c�b��@8|���'F�u���v�0!*dBI,/�X�a�'y�m�D�Y��r���t*�x��'UY:w�˺J^�I�L"�(Q�'�H!���Ɍ��H:v*�4n���'����)��-�@g��r
�' �u��ȕ�xĀ���!=CX�r
�'�T��u���=^�!RN��(����'���J����e��#A���'q���'^�`O��kF�	*!��'�ܙ)�C��t��*������'��U#��ͤF]��e�D�d��'!`%�$��<�D���@�`;:$!	�'��X�E��I:�8��J\� ��'�BĺA��xb 1Q@��9
i,h2�'Q\���� �rd�w,�7�Z���'�����ΐe*����!�L��'�D��cn�0iŌ��n_P4���� �yD8`h@#���cvn�"g"OP��nߠP�$h���_mn�T
�"O*�� ���}%t)�#GT<�EX`"O̘2p�~_�A�s$$;��=�v�'^�̻ThL�hf�܁�ꇵN�e�d�<D�ģ򢁹?��Z�Β.W�����M;D�d��/1�J�ꍔe����Հ7D�Rb匆
����
"?l�@5I6D��P�)c�p�2�I�I!<����0D�hJ�+�`v��uoɋStX�JG+3D�T�P���P*ؼ��jEv��D[A 'D���àIV�ҡ˄,'���3$D�\2d�/2D,�0�f�1A�#D���bc��3��x���J-4N2��<D�t�b���Zy��@ǳGq��-5D��ǩ�U�B�Ô� �����Ů2D�|83fY�_�<E[4&�vZL�[P*+D���c̞�z�`��Q8]�2���C)D��J�J, ��x$ASt\-���*D���f��`�@*Q/b���h�@)D��*��( V���L�`�M	�c:D�D1PJޔ^�2�`���E% TQn7D�lrV̙�(Nu���߽`͠lb`�5D���gɸ9d��J�R��h���2D���qNުz� �h���~��ҭ.D��re�0�ŀ�P~Pѫ�.D��el�	Z�@�!��M�6�4�c�:D�� �� ,X�;���==��$h;D�P��[%��!���Lc�L�1=D���G��}Ϫe�*W�!�QO9D����=��
��.6h��ba<D�,���B�!��<3t�!0�̘���7D�`ȵ�F�	n�{��1Y��D�vA;D��:�I�'8@�U��'�j����Ǡ7D���'�^k�
� ឹC�5��5D�db��N=<"P����2h���4D�����6 FX����i�j��'�2D��N�"-���v���!j�;D�8lE�Uۨ��+ܯi؈j�%D���'��!kf"��r�FĹ�F$D�d��>gΰ�,�8;�F�j�#D���xIsp��!fN�P���X�~n!���9~������[N��c��_9!�M 7��(׃XK�)۷(ݦ#>!�Wd�BEM"@��а��;$!򄘴S'2i�
�s���׬R=z!�TL����A�ʮ�rCl��v�!�Ϯl�=Gȋ(T��j �5!�䊏p9�A��.K��@�I"L^�~i!�d�;
�L���+E>b�d|��1O!�D����5�־s�R����,)!�בs�4ኡK�K�@!�"H�%!��/'�Y�KI=$��a�V#I	!�ę
*nd��,D
���%ݰ-a!�$x�AsV4Q����G�l!��H�6���*$nU�{� 0�a>x>!�D�h��8��������`ӥA4!��,�(P��I/"���W�-B'!�]�yt�d��I�Qt�"!��>a)�9�����B!�d۱jW����;��q�6B�!�^�.rD��a-�h��iVRv!��[�9�x�F�׸x�lia")���!�3|R�-3٢dK�g�!xw!�� ��r�� �&������
��`��"O"��ƃ�#S�(��I_ވ��"O��7E[ ��1�I7m3����"O�koM�:O@0�.�k����"O�mC1`V�V�N���B�z�萴"O�E��JX+�~t���� ��1��"O  �"�Φc��:T�P���}��"OBkt��E�����#8���b�"O�� ��.:|.�6zq��R�!�DCl���sF.�#=��Ag�!�ē�'r^�٦#��7�m����j�!�ę����#/��R�.���/�!���Fv��0�'[Ů��M>|!!�d�>w{���: ]b�@���K�!�DZw��m gc�[M�ɳ!hƟp�!�O;=h��Ԡ�
TR���7fI�r�!� 1r�ؐ�L4>�}���[hi!��]�P�S%R�Dy� !�U�!�dG4��4Je��H@Ea_��!�䕤5��Q[�f_:�QA���!�D	�q��5p��ټ@�/P�q�!�䎔�8Вo90�4m�Sď0�!��$%��<��e¹r�
�o{!�dT�Ya�UP@�̟k��<Q�Z�?!�$����Y(��-�V8��.]g�!��Ա%'�$��L�%���'̓�
�!���1��"�C�2_���i���.?�!�$O� ���)�$G7?�l���/�>D�����	J
� ­��S�D)���O5�yR�\*jx���	�s�z='l߹�y��D<��
�\#�<�v���y2�N�y<v!x!HY����`�$�yR$�/0��T�wb��G�R���$K��yBG�+KV;�GF�V+��P�&]��yB J�8������� �� � G��y�H����$h�
@F%Z�/���y�'G�r�f����x��	b��Ӛ�y��G�~g���D�%�ؑ����yR��%x���U.�� &�e��h���yBJ!G�� � f%���R���y��Hd����z ��˂'�
�y&Ri�"�!�*��"EG	��yb�Ӻ�*5�ܒ�����7�y�FF��(�� �*cyj
��'�y"+��j,�Hb�;�x���Ҍ�y2 D/��(dW|��(0��yBi҈k$
iz`�y$�(7'��ybg�H�,K�oԋt��y� Z��y2 Q"p�t�SeI��m��1a"�yr�ߖ���F�Ph� � 	��yz�#� q8�:���.~��w�L�R��	��
��Jw����ȓh��8�J?X��%�%"�J�J��ȓS�)�'���0��x��	0D��j�@Ea�Uvr!�5�\�O�b��ȓV�� �BκW���0��O��zX��<��q�C�	�Fs�r�&�s>U��t�(��I�Μ�B��5�ч�re����J�:�Qjb��H�z���"Ƽ�\&�ެ���&A�����@�"�"�_�w��M����@����6NBA"#͍<Ml�x���$=����Qx����$r��(ģ�M$��h�p����֬f6����-V�D��S�? ��CrOϼS^�ܳ���I�h��E"O��Pw��R�$x�o��C�t4�"O ��/C�.m"]�d��/^q�p�"OX�ъ��S��D:�<}xe"O��Q!�:[~��8�پ�H��"O��f%�5��!�B.ߥ��Qz�"Ohp��t��`	�-ա<N�:b"O~�3�N
�<g,u�j�!�T�Xr"O�I���\�h��P��D�V��UJ"O����k$2�H��)�9S�<���"OZ�8�M�5�
���H �ZD��"OѲ����7����w�j��"O̕����
 z�H�ڑ�dT�P"OJ�R�bO�
�6���C�pP�"O��C�q���ȵ,f�L)h"O�%��K�[V�`�+�//sl�h�"O.��v��2=���@��R�qJ�"O�P��Eѐ_*�����7��(�"O�,Q��S�&���C�Bň��D"O�y��L�q^z��P���|���"OT��5C@�N�V�8���i&��"Ox@s,G�M7z�����[2��"OZ�"���&IEB���B�!B�"O�`6��U�h�)C�SL��"O`�@��I;�$,�����
2�A"O�x�U��;5��X�ϙ>&d���"O�a�*?aɒǡ�)��"Of�`n��7m�Ⱥ���yeF��'"Od)[!��1aѺ�ha�R=pPP�k�"OL��P�n5 =C�oF8rc���"O�����Q:�̓��G-k�$1�"O:,��J@,Bh�u��l�7@���"O����˒-*f1��kU�s%n���"O�l�"*����tؗ�C��6�"O"4��l����Gaܶ 1�"OVP�E���2,�uFR7/�|a"O�٢嗭m9��&q��i�p"O�L�S���8�H8s�cL���`y�"O�����$dmd��s�F� ��)b�"O"}pwI��T�٣/^-*���3w"O��C�C�r3���'�Y�O��Aj�"O�,r3b��:�d��Nm�ph
�"Oh��4�ۅ3����$<���Ex�D��V+!�Th���� ��("?D�S(^o��
4��*�ٳ��;T�ؐ�l;@�H�j��W�r��7"O�iB�W������
cX�r�"OniFD�L���6-�&DB��*�"O�LJ�*�2&!s���f;D"O����\�Cu����:9v8� "O�����M�k��@�hY��e�!"O^���E0`H�)��~��R"O�x(`���s�:�.������"O�Mq� �弡q�,!Z��v"O�8q$��c[ĉ���R��4��"O�q�A-օ_V��i��&�~��w"O�����x�T���GO�_��l	a"O�,�PgI�19�c��ˤ�
�G"O<�0��'V�H�d�G?�$��"O���t���n��䎬�t���"OV�cvc��#�̼C�F�2����"O����G�3��� Z�V��"O�Q�a(е/��P�Ĭ� G���R"O�1�Cj��(8����J�d|�t�"O� ҁ�Ц	,(��`��ߴ1`6s%"O>���
�,ܢx�Éʀ �$��p"O�u(W��9�� ZBЏ:��9k`"O䁋��8�����m+@q�@"Op�3⧔ztt�)C�@n���"O��J`g��p�x������q�4m�"OV��խόQx@�'w��(�"OD�#�>&J�9����p�v�P"O����>�~�x�f��T�U��"O�!��#n�č�R���rP���"O�QtF�3 E�7GdP�2"O<��5B�+,eI��:H�C"O �au]�be$Q:�቙��9c"Ol���k>3?���C`Q�T�ʝ`7"Oء�2l*X4��t��'���sF"O1�Յlk�(� dЍa��1��"O@��6�_�1�D�А@X���(�"OP��m��lR5�E���J�"Oth�FbC*�p��r��:��4"O�
Z�|�X$.�(����G���y�c�,{gf�S�8\g�\P��y����f;������'�p5Q�EF��y��+�t��ɕ��&qh��8�yR ;Xk����#I�?���b���y�@��ɤ����:T�e鱯��yR��f8y�G1H�q�f:�y"`׼]^��"��H\�l���y��7 OHY��j�Ey�u��@:�y2����h��^�A�(h�s�̂�yb"S�V�[P�H:P>,{t�*�y��ҋ=��Q�m&l
4�Y��
�y�bW��
Ez􎚙hHp]����yRf�8��(��a؟*�Z=C��Q��y"O�s'�����Ҡ��J)�y�*[[�h���@�U�R@�� �yRG¿r�B����T�g�L�	��[�y��~�����cם�¸���$�y�@� ��ͻ384�:V���y��QN�
x� ��08=��P��yҬ:m�^�R�W�:1v�����/�yRǔ�k�*�y$��?5pF�1R���yB�;��x��� b0�剰K��yBOƜ�u�g��,ъ�Ȅ�y�.�|�Pq�0���7���yB���yR�Vd2!Е ��y;b��0�yre �p x�\�{��P�����yrc�1_�c�k?]FMk6	��yB'�x�4�+�V%�Y���^5�yr�Q%,PQ�(�XT=�⋬�y�[O�<��t,	���� #��1�y���Bo6��$��64�hB"i��y���44���4��%�t9��C�y*2+�#�&�?��͈�n��y��� Ϩ��"e�9t��p �?�yR�+X�FT1�ѶW��8����y�kY�-F�+���T.&�����y�KV+��yC�ꟴE�Ҍ1�!���y��P#�TT��*Ćk��}������yB�_�`lHh��A�a������y�K_V��Ӯ���aa'		<�yR.��nAT�r�@ Rp�1j^ �y�E�%d�f���c�&����.�y2ĉSF ��f�Ը1L�S `���y��?����6�V1]_N�`1�y
� \ ���V3Z5���3iB�������x��'H.�P�o��\�X,�SB�I (��'d�c�ʈ)ْ�2B s�t�ON��D�2j|����̒$,��A"�R�^��f�>!J�"~n�3K\|u+�ǫ=��y�b�h�.C�I�0��-����^�X$�t]�%�4C��a(�X���ԔG�d�sf�~�C�	&��X�����KFL���C�	�o�vX�Љ��mU2�
�	ݻ�C��,K�B�4�H$o��̡v($l̢C��=��!��]�M�$� ��;+=&B�ɩ� $oQ�;X�P�)�*H�C�I�z��5pWk)2�$��l�)��C䉅GP�SVEʁ?�8z!JH�TF|C�	�Y��YJ� Ei�q ���/�xC�I+���)5R�:�Ʃ��˕�Hh`C��m���󌆭NΜ)Ѣ-&��C�	&L�"Շ`��M�t��6
DC�ɭmZ��ʵ���P�c�Ƈw��B�	���(�"�~:�=��B�I�<�> ���ӄG�Fh�t�@�Q�C䉀eF&9�=[:>d"�_FB�?%}PL�'G8>�I�Sn߃�B�	�J�c�	"�iڗ����C�I�7�*��h�>-�d0S/Y�C䉍j�}xR*
�r�p+W�քS-�C�I(;��D9ec��#)6"C
�F��B䉔>2Ҵ
0NGJ� ��qb4p��B䉖�p��ٿ1�2�X�&��=�B�ɗuj �ڠf�+Z�)p6I�5O�B�ɟ~h�)���Lʦ��M�,%�dC��0p��i�Mߎ!����fѯ+��B䉂#�P�BR(qZ�������y���^�`�0d�UOv(���I���y�$	+;bf�s�h�5@����l@��y��3'��{�-ߪ?�=*�c���y�@\ ]�Vh
�L4�P�� F�y���%UY��ɚU�}	jJ��y2�3��y��#T�ʭy��"�y�_��,�;�5Q��!�0����y2�: t8鑣ȝ �!`c'ۚ�y��U�k6�us� � |)� Rr���y2�S$?�<\C�u�J1��%�y�B*^��]z��5k��Aaūݨ�y��]1!�cƅ�V��@q�J;�y�S� ������"K��9H0 S�yb�P�U1��e� ��N��ja�C��&T��tH��  v���@ݷ��B�I��N�҆��1Ae�
��ޏi�C�	�s7���;�
�h� ]�dC�	�k����dQ�ab�a�P���C�*G�<��G�Y�u.|��G��D0�C�5������(KDz�s���!!�B�I#R��0�OF�vz&��%r�B�	弹S�A)�V)�뙗�vB�	��lx�S�ܖo�iO��P�lB䉘	ӆ��5j��Z��1���	"B��')��%��Z$p
�ѢP�ZC��^=��ȝ�~��� �� ��B�	��HK��.:X�u���%��B��
kUF�Q��NA�}!���&�B�ɣ3P��q�)Z����U��>r��C�	*[�vyid�2���r�	�/��B�	�2��̑weݝe�|3M!c�:B�)� �u���$s��[��F/X0�Q"OT���l^�.5L�5a$U*�	0"O�iU��N�(�`E ��8C"O4��q�M;InM��O�i�$�4"Of����)
�H1(� ݚ�"O�{7�ֲri*y20N��h1p1"O����`.��eiD'E@Ȉ�"OB飖��8 C>�Kv*$-��Q�"O<!��,z2���ȝ�jq&�	�"O�!�6U	�����O�i6d�(A"O��bC�؆N��kanϚ2���	�"O]C��V0K妕��M��\�"(�a"O�Ha�d<2Qk7L�7y�f�h�"O����!(D�9���%��a:S"O�͡�(ƨ]+2DcPjܳ5!��J"O�0X�@��@�v�J�,*�"O�C�B>
3�L@Lܒv�*��"O^�z��]�������'��t� "O�$�(�,)������lv��F"O�ę���UK����=g,�:1"OR1�n�),ϢS ��.A�X-�e"O�]��M��H��-�å%l�Ԭӆ"O|�(ևM�k��$`�D�0%����0"O��B@O�'��`�#Տg����"Oȸi� Ӎg`v�����r)!�"OVI�b��-_���"A� #�h�[�"O޸¤K� ��a �*IbP��s"O��{PNڥ�4%[t �Jx�r�"O.����q~|M �:3|X�"OU�����8����5t��i�"O������tm�a�aBAsn�+�"O��"q
4~�(��L,)jƘ��"O��#�� /3Z������P��Ag"O��x�E�<Kq��+�Oܗ�>qq"O�D�"~���Ie�((���"O|�"��X9J�z�,�����"OX5�c��*pM�T��z�\�"O��@��M�8(�Q��~���x�"ONl$h��@D��x�i.'��% "O�Q��9q�!2p�T�;���#�"OXu9��ga\�n���2���|�!��2.3~���.ȴd�60�U�W�A�!���Y\0C�=_�@��FÐ�t!��	)Պ���GX�-��|�����!�DL�_�2�"7�ɳ.�V�B�ן$�!�ދ��y$J7D���O	�!�D[5#B$����݋��i�0� ~!�DC6�*lS�L��FsT(��Sz!�d�\1(pj���A����
�!�dׇ�v��צ��q>0��ߦ-�!�K�D4�("��o|X��#ʮ :!���>��V3{�Rm�pd��I1!�� �f��r��/o���T〾!�䈓i�Dy{$.W�& ���&!�Ė�h�fPB%%Ԯo�@C���2[�!��M�+D�x���]�L�����Q�M�!���<e�Y(2gۆ"y�����^�!�$�0�.��*�4�����֠	�!���;&b�I\�CZ��QT��!����G�&q ,I�1H�3/�!���EG�-�g��B��� �-g�!�H�����m��CnB̈t	#�!�d�2cb-�'�*XO@���A�7!�$#���˂��"@�(f��E!�� ���G;.�x�K(Q�$z<��"O�͛`��i�ܩ��W"U"���"O 4�K�'$!���d��"�"OR��@E:-1p��/��;0"O&8i6�:��s�NR�[���&"Ol�hQφXi�y�� �81�� #5"O�P`0[� �aF�(�$��"O8)�q��-
�BuXa'N�3��-R�"O���'�U�yɀE�g��=Z�F���"O�Z��P�gIHYaeQ*O�D�G"OrXQDF�+d��##&ۥm6���R"O�1I��zV� ���L�V]��"O֨�I����$bRD��H�,�a1"Ob��ei��X��`��H�3Nz�a"OL�`��Vi1�]�MM:!��"O��xd��1"l��{�KK趐�b"Oz�����3��5�'ɒ3	��]z�"O����cS L<�!	 )��-��)q�"O�t+dgʽ_�	�r��jM�=J�"O2!� ?'��7�C)QZ8��q"O��J�e¸(��ey�΁�+z�݃&"O$�b�o�?�.偗n��%p@���"OP��pE�A��C�T+;^��a�"OXifci�L�B�Ԉ ���X�"O��w)��l^�⨍�G�n�'"O�m,�|�P�@�������Z'"O��ې�J�����
~ݦ�04"O�`rc)J�+=T4��/�	�
��"OJ��b�-&�ƅ ĝAJ��!�"O��ȇJ�30"�qJf���-�-�"ON!rà(�>EX��8��B`"O,  �"�LHsD�+���c"O,a"M�d��y�%d���"O���6e-h7��N]� ���"O�u�ؤUQ4���ק4N�s<D� �F���F�Pc9|�k�N:D��)ŅZUZ1a���0Qt탅�8D�, �H�F�J�Y�eM��(����8D�0�(��Py�a��N�6��c)D��@�Ǝ?�0�`�ڼAb����%D�n�B�^x��O.H0��b� �R�<��O
T��X�7,HT[Ň�Q�<�r�D��`1��ptj�� K�<1�kۨ
9d#E`�"8P�ڣ!�q�<��H�Kx�Ls@�o��|R�H:T���c��4r~�rץ͡I�,��4(5T�<��Ë;��1��X�nA�"O�A�!A[-��(2�̜�}@U"O]��E���^���!gŽ�ybIˣ@�^1��K�~�x��F�����Of��DE�����E�D촰�����S3!�V� �fԑ�OI�_��"�#^�!���b���5��~��y!̀C�!���+�R8�#�Q�DT�R�ԏ�!�H�\�x�"۩(邹�Īբa�!�DF{?�A���=ծ`;'���O�!򄟼-X�!�R Ԧt�!b�M�>�!�/.��%�F��j7�_�a#1O�������ȃ3�إ�e ��I:Ew!�d[�$��:1f	slP��q!��H?*#�X Ab+��0��Q�']!�$H�&"�T�fd�$�2��W���lP!��t	���y��QJ�iB�W!��'f3D���*N�)N|a¨��c�!�� d�I3��]�p�x�����ء��<��4�xh
�i�.AB2�"�z�q�����I-|�F���"�+��u`�nL�jB�ɩo\\�)v@7I�B�C�K E�@C�	�Y��9�m@�),в"H9<��B�0qb1K��9�"��UҴ;ԘB�	�!h��J��:R�(88R�s�B�ɮ�Z0���B����M�����?-Ol�=A��E��8T�bG��ig �|x͓��?��kQ�X#(u��lW@�����O�<�g퓉VT�'D�2��K7
	L�<��+P1b�z��P��LAB�n�<!��L"8 �\�� ���8!�g�p�<�Al��/���i �@�5q�U�<ac��g&L\[$@2I׼�9P�i�'\�y�¬X�Vg
$�>��':Wʡ�D4E`Dp�M����Y�g|!�$�!��`�)ڵR�5��A�jp!�d?A��I�AgB0#��9�b��~a~rU��s&��;z��ta ��SKN���Cf������S������ M�M�,�b��!�d��e���P F�	Β(�[��!��==���w�ȸ7�@0.�Po!��lsڠS�=���8��eQ!��Ur��9�j��GoD��JDpH!���?	�h�gC��C@�Y��l^�:!��A�*`'!9�J�Jgl&!��O��9���Ŝ!�r�-<!�䆡'�" �!�Y�F��Ա�G/[�!�d�������EDW�>͓A� lv��[��� �0��%�H��&�Y�&�0U�q"O2���瓤-��)1i!_�B�{�"OR����/QL$���\�2C�Ec�"O*�N]�i���T�1��ڄ������(Hl2զ�.K��كN�NdC��\l�D+��y�P��@	U�x�n�����=õ�ߕ"�Vɩ1a^�I�0ԓ����o�S�O��v(, �=�&n�yjI��'����ݴ*�J]��K��>��
�'�l��/�;<����E*	���+
�'�V��G�K���yS׌~�X�(
�'=��@&�ky� ����p\|e�	�'��}�Q�/)�B �j����)��<��[�0̂��jU����J̓�hO1��5Cg��3bt�$���0^*|pJw"O�E�%�	>�����+�WpD�"OJ�[G� '����ɹ1%�H:�"O���l�-~ID+�J��	P��"OđY��V�eF�]��O;>�p1�p"On�Y3�5/v�K�HX e�|���+��ԟ"|�'Ќ���KT*8'�<�cҘ
8��	�'Ɉ��թ��4�0�s01l���'��H�'�W���[�'�*2�� ��'���R��~�P�z2�C#2���'��pT�ÄJ��2q.��`�(�'H)��ւ2ð� ��P�l���'��i�*oaf↬z��eh���y2o��Nh��*v<`q凇��0=�� Ґ�P�R2 ��Q2$����yR�x��[#�_���9ʓO:�y���T�h�P�qi����y2��$��M�E�߸Ӵ5�ɐ��yr�)�qJ@b� %2�~l�u�"*(���hO?]鑯G bǀ$p��4�&��w�4D�� ����@R)}�0U�q�4�� ��"O|!bU��`��TJ'U����0"O�����
6B�9)՗_���b�"O��q��qX��v�Ř���"OHI��V�U���b0NI�Fݲ���<�K>E��'����&-P�-[x��i�:n�p���O��$1�)�'[Ȍ)j�M��+�^)��H�6����=[\D�T��)AD4��cJT0B�%��= �{�gJ:!ʸ�����/ep���0��X�,V�TF�Y��D]5Z9����@����s�l�qG�.��Y�ȓY�h�H�*��b�Xp���1u&\��ȓ\Ҹ�#�e�"S.�J�Ē<V`݅�/��0*ƿ4ݲE;C��N�^�͓��?I��3]��	���*.5*A�FnR`�<�T��jH���d&}��Yj4��Z�<�feāͼ��iǦc�!*S��U�<��<��գ!o��>1�����NG�<�n���p���ıZ�-�d�A�<��$�C�H5bͅ0��4�s��z�<��Fċ>6К�ۢ��B�eOO<i��
H��*1+F��z�m*G �H��?��Zd��2g����Ǯ$2�R4�ȓ��m��
eϤܓ6�Eq�(��i�l\�oI5(~I�B�>T�*M��T�J ��P]s@���FA�	��������$b�3G�>.�qDx2�'��e�S�h� �����?&�=�sO�ٙ��d��9Y�M88\�$�"O���'GP�-Q��C�i�61"�"O��
��3bY�1��6x�<���"O�Ԫ���t.�0PW�ߠw5Yh"O5xb�*y�r0��C��y7��P�"O6}y̑�z��1	5��($��y��� |O��K�@�T�Ա�bI#.�{5"O~<0��Ӿ,p\Pҁ�!i�>IX�"O*T��ÛvR�Y�Aa�x�8Щ"O��J��[�i^�C@�sP����"Of*0-��f0�T����=0N���"Ov�*b��F���pbYG�
�s�"O L��	��Z�/�GN|��"O�(8�/�1A�2 [�N b���"O�8��HĬA��^�q�>��O��dR��:=�#�׼1�j$ I��!�ܬl/�%�t)��MS
z3,��W�!�Pr�vE1��O�l�@
�D�!�$��p�.�{j�-j: �R���7!���O�D���)PI@��(l�!�����9G	�0�����;%�!�D)#=
�ZRʋ�knL��@�h�a|�Y���Ɇ.	K0�(~6�ĠǤ�hn�B䉎8M�,q�������!B�\�B�	;P�N�녆O0t.��:����4Z�B�#	��Հ#M�s't̛!�3fc��G{��d�/gH�`pM��g~�[�EZ��yR�љ)TJ���$бY�&���2�ya�� ���W�~�@	�O��y�'��	KF`�r�]5p�T�i��.�y2O]�'tl+(�oZ�PH�A��y��2�"��D�'d���k%��&�0>YO>�5l܄!����/8,���}�<y�#�;L�J�B ܕJ~��2N�x�<�囱IP����k�&<��t�o�<�ݞN���'��lP�;��h�<� �d9�BVS�V�(�aG�f�F�hu"OAh������qP��F�$�"Od%���N�y�����fϼ7��Yx��'?�'��cHZH ���CCj��9�yb�'�y�,�m���P���?�����6�yG�B�H�`E����R���yҬ�&t��#�g45��!�%җØ'��{"ꐫq+���.��9��g�R0�Py���"7���d�0�L���,QE�<a'd�;ȸ��@ېX唘����J��D{�g§Z�@� E>Bp���,�Oz��$��<��h�B�E�W �	!�Ĕ}�0ԋ� ��	p�QTʎr�!��ͼp2�Q
6��[g��9�K�2��d=�O�T�6+gIhg �0R��Iũۘ�yb��ynXz����X#aG��y�g�k���13c�>��P ��	�y�9M��I	�g��bR�CFS��yb��u��,�ɶ4��@���y��ܿA�#����+*����S��yNG���m�"���C��ڣ���?�ODx���4��]��	���Y�@"O̭Adߘc��Ó(
�O�^Ѷ"OHi��)K��RA*g^R@�X�"O� ������҆�C�?8�[�"Ot= -E6c ��Q5f�_θ�f"O���æT"�M�q$׸3��Qf"O� 
���� /��`f#؎|L}"�"ONa��͂� �`��G�61�:�A6"O>�*s����&�7τ�"O�	��i��a�H�yY�e���20"O��s"�[�$�����$ǰMC�"Op� �dC���k�d��"O��ؤ/S�BX��D�8[�I�"O���(T���ܝ>��< t"O�̠���#t�y�L`"OF���KT/w����Mޢa"��"O��Ӏ�[� � kb.S J���"O�Tr���(	lqze,�%X�(��1"O�E�RK
 w��y(���_��q*w"Ot]�a��zq$Bu�qO2��"O���cu�|�V�pM�I�"OD���ЙV�Ё�����!C"O~�!�ʚ.ը2G���u�S"O$CBhȣk]�ɺSo����h�"O`X��
$A�)PL	2Go� BA"O ��eU͒,"�,W<X�%
d"O��C�n!ma*�0�T��P]*4"O¹h�.ՆH��( !��Zc�E�R"O^�Z0��(�d��d_+(��j�"O�ċ �A���W풜@�E��"Or�QU+:Ժ���+J�*M��y�"O� 3��*,B\��פ_�@�@"O4u�w�Ɛb��Q��xӒ"Of%i2/@��yx�A��N�
ģ�"O��@gm]s yXA"�� �
�>OB�=E���q=��`�"�b��4���y��7`Ή��
I�|2f�G^��y�o�t��Co������I�y�&
�[��0�T�e��0���B=�yR%�P�1p��m���Z� ��y"ō�STlT �j�&k"5�����y�*�	Uղ�K�M��l`v�`��� �ў"~�:M��#��B�	̽goĉ��S�? (�jD��$od����b�I�ޡ�d"O(`��X�|�� ���ȥ {�Ūt�����)B�Jl\d��u�(��&��9!�Y!�xl��%D3n���Z�d�7�!��?H5�d �B���s�d�v�!�$�rw����n�	^:�Y{�%����%�S�O��ErfE�F���'ۮ����	�'3��0�֓! ���t,�(t�x	�'�B٣���8s m���n���Ѝy��)擊~������[V�a�	EPC�ɑ��ŉ�T�����ֺ)%�B�I�Ra��!�L��-�B��J!�C���s�Oؘ��i�Ҭܗ_(H���%6D��Tm=6�t�@���K��0#F.D��Pl� Bq���X
'��$�#�*D��P,=���9���S����bJ-��hO�S.?�!5�N�5�r�V�
�E)�B�I1?"�@�� �N���	�9#�B䉕
�L��7�Q)W.�h��B��d�.Q)B�^�I����#ɏ;DB�I&7@�q��i�;u�8i���)u�RC�	�7E�
��K:&�`�qo���B��0DΔ��퐺=��t�lw��C�	�p�����Ah���B�	eNT����s�0�
�
k�B�ɘ2f.����.A.=��!��Q�C��^^�U�#��!֕����{�C�I3A �͋>���E�$n�VC�	�_�<]J��L	�l��Ì�n��C�	"2\�pq3 Bc����1��'G�vC��p$:q���j ��)*;DC䉐���� $D�)�zMY�MT|�zB�	9tlBä��dh�+�e޻J�~B��%c�~E���NJ�d)Z�đ;,vB�	�Bp�c֍�:0�J!��!$*B�I�j�"�haa�vzP}��N��	B�I%]�
u+��۟
��D�CYVB�	r�FL�aɃ?6�����	ߖ7�@B䉞t�H�1��W��� 6fݢE�zB��?�8Z���U@f�K�,kV�C�I)�2	��#�R�k3�ڋ=e�C�	!Ƅ��	́Z��(YCA��\�C��(|�)7J�}d�\���4Vj2C�a�HK�NyԤ(�Cw�w�	Y�O�����,<�=hv�]�$k��	�'����j?4�e�*Ðe�']�|9rN��Y�T�;� �$G����'l�1y0Ʌ~�A�2O��g�4H��'��Q�s�գ;����c_]�t��'�,� *�)ZӠ]��C U�*
�'6��a�j�&�Hy�"�ʲ��y[�'p~�
��5"�#�LԺ-����'��"����mH l�V1�>P�'U��ks�8�*�@��J���'�&�7��7L�^d�4ƃ~]:�����/�S��\�8vX�%�T#>�N�����yB	!��	�#"Ѷ2@�ݓ��0�y��٪-y�)ɥ�=,(�� U�1�y�aH3&�Lp��/DXH�dn��y�E�-%Cb�@��N� �������y����)�4�a!G�;(�R\�sdT�y�I������(4��	��yKLs��ZS�ƚ)(y��E��y�]�:�
��˖2o&hH����y
� R��M	%rYȢf�.MA���2"O� ��.K��Ru�E2L+�I��"O�	���֋U�
- ��p��d"O�s��0a01�SW�-�H�[#"O
9�f-�0�<�����-�@��V"O�*�-WwI� �c-Q/>�JeX�"OŰ�Β7`Ё���>U�@Uw"O}����@ml�K�$b��5A@�'��'�XA�A�e>����)R�VH��i�'l�@0�o��;}~�(�D%B�HL��'z�����'3$tA�f�*P�$Yz
�'��}����9���2S�Q�U�`�	�'�\d�a)�(J,hɑ��r�%�	�'�"E�r��j$��I����9"���'��U+���,~�l2�[q:V���?I*O�eh��U�<v�	0�wo�$�"O�T����8�zوqKԝMx,�p"Oֹ����m���`���xb4b�"OH�YgOK���2�H���~咖"O�x��Z�4��
�Q���"O�H�Y4S許�fȿa$8"O��V4@�q�� u�4���'��O�r���*5Fȅ��'/J�Ds&"O����ʯu�F����¹<�n��6"O�<y���n��ċ�׋�^z�"O�d�$�Q D���3y�ʵ:�"O�Y۵�_/a�h��0�ތn�@H�"O�:��������j��c��#*O�]@ӉÕ0���a�`O�huա�'���% .^"쩙�G14�l�H�'��H�,7 ��Ur���B�4��'�nˑ�!�`�p��C�p���:
�'��xh��>Lp��U��*o5Zp�	�'I��c�n�y���� O�_f��',���X*	�UXC*�
����'a�i��hܴi�K�_=�a0P�U|��&�xZ��L����6˔�R� ��6D��C7KL}Y#��"��S�8D�dr_��qHp)Ã��l��`Z�"O�]!�hٳg*\`2�Q N����"OZA§ Z�`lɚ���$�@Ey"Ojy����I��I�e�_�V�T���"O
�' F�M}��	�a�'�z�kA�'���O-�\s�V�B�%��(N5�B��2 �
��"6�T���T5]ľB�I�i,��2bԏM��@y�iFC_�B�I189�D�MȐ)�L��G�ȬB�	����en�.S@Ǆ�,\�C�>3�h���V5'䌕 Nv]�C�	:V*Q24�
?o~X5 @�S\z��:�ę�_�~H���P�|�&h��̀J!򤟧c)�5qva39Ʊ�b�T Y/!�/;�x�6!P2"`<2���a:!����`i�Ck ��b9��!"!������`s�Xp_��i�"OڱJu.��8S|j�_U��xY�"Ot�ʷ�U �h����$36�0�G�'�	:Ws��¢@�LQ��!T��'(�B�	6w ���V�I�t9�7�ï}ZFC�ɟR&��EF��q������C�P�C�IDD�]Wa�1]�A�&&�+<ZB�	EV�aP���{hQ��d��&YB�I�M�j���Q p]	�����B��!h�Z=�V�W�*�X-�b ��h�B����� �uY����w�R�[�&ٳ<���"OR����!7M8�:6��^.b%��"O�A6jM 1�C��dyf�a�"O|t [u�إ"�OH*^�H�)s��A����'�I�z���bV�mԆmȕFϘo�C�IL�媁�KZv�%,��.��C�	�>��JW��W
��Z�&�4ZRC�=R�D�	�h^�+��kU�)S:C�	�IG��g�,P
�9p�H�:B�	  x�q@��	Vw�YJ��%q,B�I0}x|X��]1"ݎ	[���i��C�I�&��AR���:�˔}�Pe�ȓ(�^@����J�J���0��ȓ3@\U��n��*�C�
Z��\��A{^�3��Q���Z��ڄ
�����'��`��N�S�6
�����|��'���Ȓ�\�;��80G�!t����'H<{�$O/E� =s���8l���:	�'���zƋC4!�� �*1�&�C�'��	)0�s�X2�π�w�vtQ�'9�Lc%K�*fXX&+�s %��'{�׏�?>��	�
࡛'���+!q�x�⡋�~�]n�;�y�	�7U�6%��.X�?R�#T�޿�y��
X�j�C�2H�h���yr�M��%�Ĉ5pR���1΅�yR��g3�����Чm� |�Ѥ�%�yr�]2��,iQc�e�~K�( ��yB���~�"�+�G+h� l!��M��O:��AoӤ1BV��� ·�/j�!�d�.5�R�Q���y����qޮ"&!�Ď�p�͉A���FB��X�w|!��?�ء4f
i� ir�	^{�!�#��qa�iS˼PE+�"T!�$�I�Ȩ!���D�4��� ~�!��+P���Ǎ»'���B)��z	1O���DJ&)� ��uC���=A���!��X�lP�"_�/f��!��)!�1O���$�sQTrSd̔^�Б�C5A!�[�^�`�+\�d�ڄ�9U!�	�6�����Q�ap��==e!�$`{rq��Dʸ~⮕ pL�HY!�KN�JDp�	��/��c3�W	Q1O����kQ�D��'ɳ<0��F�@�;5���O��"|���7$��#�8a�h$y1�&}��-�ȓ�\��a��K�5��[�]�Px�'� ���@ع{�5��
I;��(�'� ��r�A u���6��&5�HY��'!B��ݘtk�E�])=2(��'K,ݘ�%f("�F��3_d���'�$��F������t`�
,�L��Od�=E��D�Wt� ��<q:��O���yb��'v>�jc�]�^
1��ݸH�"�x�'��m#rc�	I�nd��F+E��L[�'y��QtJU���+��I+@9��B�'�PeΗ�d��$yw��:����'/b�8�+�N|�TQ�ٸ6�^mK�'Q�֩χ[A8)Q��B@�;�'�҈^ �@$z��UC��9w#ȭ�Od�Ob�D?��_!|�̸�&�wp
�h�̑�2�!�Ī����a��1^�U H!����4�+6j��Y�\Q��!96!�DM�/'�:S�G#BX��k��=5!�DC�HUJ�I�� <`�AV*	��!�� v�;��دJ�c"� `��t1"O��0"��ID���A��� ��hx�'��'gR�ch����W�ɖ]�<
�'L�l�dفc��Փ�j^]˜��'
��Y�D�>5i�σ�\%�+�'Ú!���X>�Ufj�2,YH-��'F��+)�"�x�N!���J�'�@�"�!I��T��Z�M"ܳ�'I�PP��z�h��DMWV�:��!��:t*�"��Ih�cՄ�3j����*OZ�O?�I2]�!@��
�?���G�ܮu�DB�4uK�tC� W��8��J\�JezB�ɉY'��x6`�����zG�.G�JB�I9q�p�{e�5,Ll�WX4(�>B��%`�@�WI�g[X#B�Ԡ{k�C��as��O� E� ��� ��䓛hO�	��#�*�#vh�]������'-�Qj�)/�(�8���Q�̐��'�ڠ��%��~Fh�灝ub 8�'���(j�>?F,Z�`�ztI�'\^�)��Tv�9Ӄ� ��
�'�pԋW \�"&V$�G�t �Mюy�)��_�����G�5��z���q�xc�Ї�;T`� �	zGV|�q�d���-�i"���
��s��m�W�\�ܵ�ȓpR(�aD��9;4(1.b\���#���eJ��P����مȓad"2F��V�\�j�@�zE��P�V�8q�����"�v8�ȓG����#	B�%6��b�,��V��y���iy"��]�!5� P�6-2��N7�y"IE�p
��B��<O~Т��U�y2��DhJF�E88�@a��A7�y҈��d
nt��j�=ǀ�R�D��ў"~�E�&]{�J�,d�EEw��5���ny�κ^�Т*��b�B�3��	4�yROK�\�N)����"(���*��y�	+Z����n�Bb91����'%��'!$\C�A��P��T+�!����'�p�H���H�eJ$-��6�ry#�'����őxX��[���2,�t��O��=E�t��y�VaXbH�}FVt"R�M�y�鄬vΠ(��1K��&�y��˗J��|J`m\A��%i��y��5���E-69���)ݕ=��	Fx���)M�>��`���	�Z��0��.D�0�NW�a����m��;s���+D���2	*f>��j��տ2'��
�i���Ik�S�OjF�`B���$Z��ϧS����	ӓ��'~�A��)C�2��8�+�a�±#�'�%\����`��	��'hRn�u�&���6R�e�eÎ��D �OryT+�]V�1H�6-^��a	�'%\\b�Q<98L�CD�.:���	�'ot� T�B:D�h(	_Xob���'����7�#v4,���x�p���O
�=E���ȧ.O��r��H� xd	Y&����'6�{�]\Ft����.�jH�U#M�0>yL>��+:�˄��hX~x�[>
B�I�!�\�)^QԾT�1*�#o2"C�I��U�f	Q��|����..C�ɠ1ET=��<[6�D1�GC�n��B�I\�4�ӳH���N9�EF.g�*�	w����P�������B	Sd� }�)��5���<E���� <��g�9	�ZXр嚠3p�܀�"OXT`���xw�Ի�D�$M:X�"O�-�CA$(�A��U
a�1��"Ot���QͶx�3I@[[�$�"OV}X ��WPT��);If�"O�ոd#
�B�x��U �лD�:�S��y�Π*����tiR�Ɛ{1 �0=i����
�m1�, ��{�ǐX��'��Id�'��		�0	�hz:�IBS��y�i�S��;t�F1}��䡅���y�$�rdF�Cn{è J�$A%�yZi):t�E�P*,X��i��Q��zC�3|n��@
�%Y����@
T�fC�ɧ{]\Ppv��!��0R#�Ԙ7C�C�I)���K�^Ly�nSL�#<��m�J(	��֎�dE�$�p�ȓo�L�i�&�M��r��*}F�ȓ��ْ1@B-B�x0�7.�&Kc�e�ȓ!�������U�n�i�f��Cr��r�	�v��!P�Qh��D�����0���*_�6��o	>7��M4�7�?��P	r�Q;?���+�"�Aꃣ�dU���I�|A��|˶	��K���6�HaA�rc���>,A sI�9��M����w��T�ȓm+xh�t,2���SR��fX�d��j��`TFM�\`f9V"[�U�:l�ȓ��<B�f�P<��8v��,t�U�ȓM���E��=J��8�a�"V����ȓI2A"�	!`�1��X�P�ȓh��0DBס1�LTqC�KU�p��9�h��b�� +¬Rң�WRN��ȓRԠ���![jDd:���-(�2���N@	�Bϣ'3�%�����TȆȓY��L)`c�,x"r0�4�U���ȇȓ?q����BA�]������jQ(х�(�@�L�6;[*�����Uǲ�ȓW���T�*-���h�%ۼA��pFd�,O=�Bb�V{�H��ȓr���poѕsq��&p~��	D�Ip�@e��+�6�Ztj��(2RB�#E40�p�J�/ 6�S��;fn����O�ʓndz���a�!�����J�J�����s���C|�h��&� w�`��" D�L���<i(U�a�:*U$q�+D�����G7���򠗓e�$����.D�x-C�% ��7��|\��#�+D��"��F.y�893�*��f��I�&�)D���@� �R��@�H+�����H*�O�˓J�KM��ub�ȸe-Q�~�~Մ�]mPU5K�,.'�|h��M�,>D��ȓxVLIH׃�A�`e�$�4"JP�ȓ{L\t�2�W!+	<%�@�''F��ȓz�U�� &4,�s�I�+!�\��ȓr���*�kI���b�K�*Z5�I��j���S���|DJ4*d�V-4�`a���?����*A@X�֫ @�v��eE!��'<�y�O]����A1!��"h�E��d��y�e_�L���iM6��c$�ټ�y��ĳn|�L� ��"?	��P�#��y"�ZFL�,�U�B$=Ԝ��#�\��y��9J8�oՀ7�"Qc�(��yHͦy�ܸDB�*$u��zE��<�y�mS�TU�T0�Kݨp�­��/�y
� �0 fل����X�#�"Odh�Iw�!�P��<�]��"O=�Ckoa����`N6Pr���@"O<@*#@��-Q�pr���(8�#�"O�Acr��\2i�BE��d���4"O�Uy����'�u��c�}��"O*]9�O�=�N��1��9¨�@"O�`�Q��	��So�C��@"O�,��̚XS:%KGoY^���a"O8�K߳G<a���*����E"OJ��:���xR����e�t�D��y�	NYm��2$̀��l��ĥ��y�闯������;s�%�C`<�y"�K��qp���*-������1�yc�/F����c��'�D�ɂ��y��~�̀#�L�= ���S��U�yb��P��%�0�ͩmo���d֕�yb
�7rn`��0)��d�y�CXfm�TJ�({����5�y�`�%0c���d���y�lexw/���y�QF�\��1��n�L!b��?�y>E>�"�S�j:����T��yr���iO�a9φJ�z页Н�y�/wn;s�KG����4$�ybg�;� �а�n��q�5���yBbq�E�L>#��H��BD	���	�'fL�emӎ.h�m�1�2|�����'e$�rE�B�邐��Ċ#
.�%��'��S�+��
��H�2�;r�ڝ�'�d�a�nčH�$��D�u~���
�'��+���bĄ����0r\�)�	�';���vY�h%�v�1k��=��'�y�g�؉;:��G���+jB�y�'�B����Y���	�M	yujaZ�'f��P��7)�����pZNУ
�'�nq·,�$�8( Q�� f�&<j	�'�R����Ȼt2\Ip�ՊN�f�	�'���k���}?���7j�HD2-�	�'3� ��'��Fl vEb�	�'�	˳��/�f����G�zL�1�'h*����^������n
m��'=$�0I.O�lj��ւ1�(��'0���
�/e(�l��I��%F��[�'L��C�EYX��E�)eN���'O����#)0���\��L�'��	i�a��qpHR0-���t���'��Q3-J��M�v*��\��
�'�<E�d�jk��aK1;�m!
�'g,=� �� _N�N��K7���	�'آ8���O=����Aux�Q#	�'�H��� ~�b5�"���m�����'M�Tq���1iq�h˅�[ T��B
�'&�pZ�l��x�fP� _
Ȍe3
�'��x1�HH�5�>AX$�	�B���')�ijC̈@S�B4% �"���'�8$;gZs���SC�aWڼ�
�'��lJv�?,���R��U���
	�'a�����Z�O�H,�a���y��Pך� .ELI*Q��%�y��Ϸ[zFX��H?��H�Ɏ�y2vGL$H�@,68�I�>�y�c�=cd�<�"��=�pD���y�þ2��ɱ�<��-�)���y��-2U�Z �>�P�ub߈�y
� ���i	6'C�	�IR�^��p�"Oڱ�&�%O���a4�&u�5�"O���	BP'��C k�M��"O�H� �_(F�MK�f� 9�A"OX��gL�FD�#��U���"Oҁ У0Cr��h&�9T��h�"O28��bL�a� �C���i}��Z"Ofm�W��]��r�a+^o���"O�H�HΧA�4Pѓ�F�y�"O��'��,�`x�f��`��%{g"O>�(GnI@�@�[��'W@��)�"O�y	Ɗ̩$�V)d��c3���"O�20�l������`����"O&���.|hfU�g�'jᖽ�#"O��p��)G��'˖	s����P"O�%���?�4��1�8�T�P�"O�Iv#� r�ш�mY8Rr�ڕ"O¬��(�L3ܼdoK��ha4��?�If*o:�h�GOf���e� �1��
��i�ǋߎ�z��ȓI����bY7�|x`,��-�(�ȓ �Qy���{dĠ�)��^�x��ȓ|�b��ռ'��d�0���wX\���
3��	G��6��7��g�v|��~�X�p'	;P��a�U�E6"zl���iidp@s�MAۤ�[��˄NdC�	�+�:�bq��/3@LQ�Ãu�B��[쎼���ΚY�����W.\B�	%#�R�b C'2f�Eʞ/74B�	�W�U��(�]IY�	�"j��B䉧P��jV��L�9$-�.J>nB�ɴm&윓�@U uϜ��(�g�VB䉜]�`@��&Q7`ݚ�bW`��$�pB�	�F�.��0&�7E�|���PC�	�		�|jw(�Z�xՍN(x\C�ɮ5�$��aD�x�� �%�}��B�ɍGK� h�M/|Q̈!��<A�fB�I�\��QT�
<Pv�̴[�8B��))RjI�-E<nw>Ա��xp*B䉅PR���`ڛN�����%�JC䉩htD\��<v;�H���?�\B䉴<%h�X�B�� ��఑I�}9$B�	�+z޴i�g�ZЫi�y
B��y�X]"4֠f����o��j��C�	��M�� �+}��æ�;;�C�I�@�n�cS�h��*�`��C��@��b�%>{�b͋&���Hy��d�7U���G�G��2��ڳ7�!��<M e����'x�mC��R�2�!�ƢO�R��'�5W܅[�#��3�!�dŐ1��AU�*RP����$�!�DH�e���FK|P�a��
�!�� �4��� 5� }�
�0G!ێ.�!���� �����=Jo$m�P��	�!�NQ�(4G�XXp��O���!��i����J�VD&5��M�
*�!��/N���90�216�p�WM__!��C+N��]�ӣK�-�T�u��H�!򄐖1(rm+��S�ejh+��)w�!���V���:%"X,"�c��+` !�E�`y���&C]@�i4��0�!�D�)y�� ФMP*{+�)QnO�#�!�qix�N�\�5���1�!򤙥,*b�s��T�	3�Ҫu�!�� h���G�#Q�!� @��Cq0�KC"O�X!�세$sL9[g.�:Dj�0j"O�cѪ���,���;G�@1 "OFe�A�T54�u����%0@�3A"O��+^�r��"G��7\	�Ջ�"Ox��0JR =5�G:�ʠ�"O(��A�C��D�`Du"O  �ĭ� V��9d�ǋ}�te"O����
\�0d�v�0n�k3!��n���a�c��
<�� �9-!�dʨ��-3!��.T0-Q6�×6�!��W�N殭��hB�q;r��e#Y�#k!�Dszt�CH�PվU�S�ɤ9]!�Z�9ܝA�H��a�&Y1�B0A!����ȃ�ˉb(`�eH�rI!�$A�d�VH��g��+gNd�3(�!)!�1NEX�a�Ԇ3X�P�Q�H�}1!��)?:p�Ç++6`�y��&��&!�R65Ĩ ��(s+�)rQ�0"!�䒾*��<�D�R�h��m�!�DJ)	d:���Y�R�;�+,(�!��89t �����E�Rq �W�h�!����U� �W�<��$��a܁B�!�䗆]4�t T�S�T�h��>&!�d��r��	��^�P}�S(^!�!�$^�^wD�0B��m�-p�G՗�!���Ԙ��#*��V�:���	v7!��Y�p����ė~�~|�s�C� !�$��Ur�a���g�t�pt�.�!�$�
�D�*��1���ƃ�	 !�DL��V|���G��(k2%:K!�Ī;�t�A�I�Sw�3bD��p!��Ū��Pw
�&~mD`a��n!�$#c��8;��.fLmbDRm!�I�3f��s`�h��ቍ7W�!�$N�5�Q�F�ɑ!`��[f�ME!�$¡Q��i�Ԣ�-�<-r�l0)�!�d̿0��|����2C�JF��!�D��}���aMOHIX�J0,V�y�!�DC>N�l��霦.��Ӑ��E!�䘮O�8K�J͘=�D��"c�"
.!�Dc�H#���84�|�8% B;!����LY[�lΎIhL���&W!�K�*�������Pa���GoF!�-.���HW2N��D�*դ}1!�D"M���o��/l\M D�#S�!��љp|�
``u���֏ä�!���-gP�LKsiH� ���raՌ[i!��B2	�<��kN)�m� �6u!��<\��*�4Vv&):���%q!��M	g�@���U�&sV��p�_/9�!��yV(u��� Ydf;��9�!�$�� ���ȓ%pT��4�0�!� 5�h�Id�<B5�䊐p�!�T�H$PƍF/J$ڍP)�e�!�D�dO6�S'H�F$`Xؕ�Ga�!�߷d�Ѫ%�(6n�
Ԍ�nG!�D���m�w�ۓ&Sl�H�ş4)!�D��Kq���G��/4��*�a�!���:)J#C�e����ï��VF!��̫�L5B @�>WA�M��mټg-!��=~h
����X*\�(2$�!�.�Hq{�Ma�~��׬a�!�dG�`[�$S�	��JA�'�Q��!�� ���D� =P��4�Q	�\�R\��"O�U�3,C���3�H	�4x{�"O�D�K�^��Q��f_�>�dPr�"ORԨ51,���co۩+z��"O���*�S&��gN/~�y�"O�p�0�]#'	�1�Q��,t�l���"Ol�b�N4��mC��UPg"O��zu�TDń����O<h��"O�i�R*�H<�(��ρ&���"O2 1E���J5	qV�ŷq��`��"O���mK?qK���i
�X�"O�Y��Ǯ^�\��n5%�LĲ�"O � A�͚-��U�%@<qH��"O�ᛑM��9��C�E5I���2�"Oެ�Q@�'O�\�h#d��*�ְ(�"O��i�H�FYR��#�,Q�i��"Oɓf��8�>��,^=[ް�&"O.�aE�x`�5#kO�OoB1��"O֕�2Ɉ�?�P4ix��@��2D��A.ʣI
�)8PLC��JX`!+1D� �&�c�Cta �>�b�S��<D��s!�R�X'�1Ht�߅�b#�;D�D)��&=l����Y�k�`�:��Y��ħ?Ǿ@��_#�V1悝~$�]��l�Tdy2�<b�HGl���~<Ey��'�^I�6�ي##ީ��υ�e�Hy�'�D�2���M�\9!塌�[�m�
�'���Q��Ы��Xg�+�'<p�z%aƽႤ 	�>_�2�	�'�QI�nȻo�\��E�L	]��ۈy��LS���O�(%y�T�F����%j�	l��'ȶ�(�X�,�B�i��;�f���d#,Oz��dKG:p�����OS����a"O\͊Q!V)Bら�S�N�����"O��cݼl��X��$ƵZ�Ju�"O��&D]<0�Va���Tx����"O�U��c�,u�5���C�9�Bi��"O��y"�Z7V���B�pY"�qp"O&�bt�{ٞ����[$U�"O
�t�ėd|� T��!%"-�"Oh��h.�L��E��8���nx��pC��IZ�[d@Ə�0}Z4�4D�0!C�\<���3�`B�vt̜@ D�<�֜�~0цa��x�cw$,D�(��c�q�♈7�޸ R�0u�-D��#��.[��s���>$�BE�a++D����U�⸒$倆3�:��B�+D���CZA8q��[Q�D�w#+D�sfN�
z�C�eV�Q�R�2!L<D��� $��+���q�T*�����:D���©�37R�a�m)?{ 0b��7D�\2g��yS0����O1 �8�{a4D����7 �Dl��(F�T�R'�4D�th��(����R��*�3D��x��ZK��ؒ��1o���t�<D�\(u��Z@|( !���"���8�;D��xR�L(� �c
ך騁$9D�Xz���71����CM�<���!F<D���Z�i-	�fV�M�X���9D�蓒�F>v�Z�K��ԱZ_$SQ�"D���#�E}	�Q�� 	�1$�?D�H�ug-Sn9QA퉑2�|�g>D��en�.(�a8�D!F��8:U�;D��C�
ʭ)} -��^�Ɯ��M=D�� �Q����'�<�V!׺T��Y�"O�}Qrk	1O��i'�ϯ{�ͺ�"O��#�S�r!ʔq�	ܿA���h�"O�T�T�PQ黇�O >���Jt"O�U�� غ�V�3bK�����"O<�#��H��:�@�KҀ�L��u"OX�M�ȡ�-�)����"O���4�ъK7���f/�|��*s"O��X?O���f�M
D��h�<�wJ�'��a�qͼ:Ԏ#�y�OԦ8}�Ց  S�TOii�&ٸ�y��?2��E�0����C}kM�	�'��8���"
�E��DX-ubL�	�'f\8�B,"�����"Ƌc��X	�'f.�zr��"U&:�aQ��_׊�9	�' �80L�+.k�(�-�$!��QR	�'ꔨ�2�ˑC;~A��+�.S J	�'��̘ыև-AZ�ۗ@G� ��:�'��ѣk2|@  9�H��.���'�8�P�L,s� ��fmK4�l��ʓ&�%���M�/$�F�?,L��ȓ�PaKm�t�)�͔�$x ��pD����M+}�!�rOǯVh�ȓW\��qn�Vv�G���~Q����c�'rp��.�-�<���J�P��.�9	�@��Q�ƾ~����9���PC�5P�Ν�T��!�^��ȓz~<)�Ə M�.0�$�T�:�fą������9FxjrO�p�",�ȓn���1�V�+�r!㎮T��7�T�X���7��1�ˋ*}�p�ȓ#9��#��ٗ��Z.�������
����Eqt&�
g�R0�ȓ5�t)!�Q�(A&_�X���ȓ=�
��n�� 4̰�t�Eb<  ��S�� L(� Q����P�)�ȓ�9�Պ[�:8�G��?,!:8��i'`��gP��
Yzk[�[`��TS*�p�.�N�^2�H؄
��h���P��u�$q�|8!#��>:���ȓP��E���]�%n�-�� �;"�d��r��0��K�5�,�$��p�R��ȓjIR��"_��x��8>�jE��q�<�A�Fل_v8�� e��fhq���2aub�{
�M����Z$��ȓqszE1�J�~+���a�Z�$u��2��=1�ď��}�R���(�����6!�5xT���h
���ȓB��H��9��)���D�1��b��c��<�.�z���pf�Ʉȓq�^��I�(Mx��4c٨|�~��,<&�����/K��Kə%�6���gF���C	�>%"A�G֒�¨�ȓx_����GҾgVf�����:���ȓzlA��A�3-'y�!��=GB�9��dL*E��1l�#�g7cW�M�ȓNMް2PH�PBH�C�j�9�Ćȓ!��r�d��F��is�$��\X����l���,ۨU��-+����/�f$��J�x3% �$s�J�#G�\T��D�F0�F�5	����֋Z!u�0���b���"�g�,j��1z�[6k��q��1�,�CbL�f�J\`�W�y��A�+���5a� ��j������S�? �L��K%z@�Uf_���T"O��sC�� h��S��0p>����"O2*�+�Vp�Š�"�m�Z�u"O�Y&�:��p�T��w2N��`"Of� �+'P�h1��vv�"�"OF�qm�;"5H��A�834�qG"O�	��/��U�ЙSV�܁/t��"O*������<	��Z��A;g2"ű5"Ol(�Gmλh�d��,>D�Ae"O���GƱG�8qV	���"OV9���c �a�$+ɖq	�z�"O����l>����<[��4��"Oa&R�&#����^�7�<9E"O&�26�ƑT���"�B)�"Ob�S�Mg�eR�`�3j�:��v"O`��bF�?��y�OC�o��G"O������d5��W�	~b�"O�x闠�2�����G�Go~eх"O~�zE�S�+oZ����U� ��"O� �R�4N��p���sC�Tqr"O"4�#�n2�� G�Я~0d�ȷ"O�8�����*"z<�c���h4�D�W"O `��%���ʸ95ڮ|��m:4"O��BY�\��u[r�
a�j�S�"O��sV���s<ZI�T�G�`�F���"O���Q	�W�<@@bBHZ��$"O@��&/��5=@I�� "�Z���"O���R��7*FF�ZwB�y��4��"O]AV'B7�&��f�/N$P!�7"O᠀��'�h)K��Qn1�&"O�5�g+�!C���B%�=�9��"O�ث�&�������cмP��E"O��'g�
sB�h��N|��
"O�R� �n��-��^Z,Mc�"O�xX�޲rJ��P§�efq�"O��Y"���i����&�C3��"�"O:����!�^(;s��1v�1 "O�}�c�\�j^e)�	��P��u"O����F	�}2�Y�cB��9���x'"O��7��Qc��S�a��x
�"Oꄳ6% MT���"c���
""O�	À�='f����6�2"O�$1��6רm����:R�$�U"O>����Ͻ_�X�Ұ��.6��%���x>Q���ƚ���k�LQ?p��yЊ8D���E@�6��B�Z2SZ��M4lOl➨3���4`a��	�>,6u��1D�P ($�t kp�Vi@��1u(%�	N��ħK��qѦM%(��*��=20��4b|�s'\�G\֨g���A��+��T2!��?h�d�Q�_2Y2X�ȓ��U{Se߷-W���^.\r�C�	S?�� [(;4�Q��Y!=�C�I�-{���Ͽw�*�
��tC䉳;� ��� Yre��F˗"_b�<���)�i�9C�|C��	+N�Q�p�K�A!�D
�ur�p0��3e`2�R�kJ{�ў̇�I�J��С�O"ʌ����*��?����<4�xa�s�G<�jFOG�)$!�d@�?�x=S%&R!& ���w�   �Ol㟴�=����v�`���8!^D���a�h�<�v($8���*ŬԲ�5��IEe�<��a3#v�qI�@/vj�D" ��L���hO�]0�x �����v�s��S�? VP+�&�=0�<9�OQ�3����2�xB�)��$�
��ěf�Eh��ށF�bB��*����6(r���)y���ȓ3�1Te��BHஃ�(�6���4�r1��A�
c��
��P�#4D��K�L	�gbB�1�#��]5G5D�l6.B�&LP���ep�5ۖi3D�8j�p��i��C�{b`B7
=�Ot�ɜ^RЀ�CC-j.B�KQ6��C��<)΁�T(M�fnȁč�?�C�I?C$$�ID<���L�B��2F5��ہFT�6%2�8�(ƧU)��'�ў�?�F��^4�ەm˙vҠa��*�hO?��G�L���JТY�^�T�P�nJqO���$N�bkքJw�K�##�S��;�Ol0��\�v���QC�8b�0�"O�����E�vT�\[��ú(� �U"O�������ن]���+��d �<����b��舴�ӽA��Tk�'�_�<�r(غv�4Á'<@��p��*�_�<�燾?���2�h!u�U��A@\�<�/9���V��Z�*���Z~H<� �=\�, ˦B4%t.DC�2�!�D�\�|a���'g�x,��e[K�!�d�����0fJ�8�e��`�!�A4�.A3�J�G֌����O�!�Y }�@�
uL��'E�h�SBː�!���M-\����0)��8��ڗ(�!�ӗ<�Z�Z���H������#D���Q�ZF�=9�3(�P=8Q#0OfJB�I�JN��e��%s����enC�	i�FU�OΈ%�bn�6ŤC�I�R�^�9��_�-Hf�)�iՠ����޴�M�L>�-OQ>5;7��
=~�l{dဓ)�*	�ve#D��QW坾2�愫�Děs�`�k�`.D���C�R<PJ~h�Dρ8z��a0፸��x��T�Q|l�1�j��aǔ�3 ay�Þp�Z$T�Vl�e,��� �]����D2c*:5�� $;���>	�{"�	�� ����w�$X�Ȁ�H[!C�!򤗉I�m7E�i�ڬ�t�_X�1O.�=�|��R
5�N�C$��3��INYQ?1
���p�t,"�TՈ&���]hf��Of����4��O��Z�/�-蝁��2240��d"O�������r"3�ǚ $J���/LOD�sSYE�2x���az�(�"��a>yq��F�fh@��#{ l���8�I. ]az�`îam��(�?�N����M��?�M���O���f�H�@իDZ	����$���IA<�0�ȹ�.�H�F�""�����x�<�T
_�b�����$&�V 3g�s�<��fC�e��򢧅�_� ���V�<�R� ��L�VeW7��y�.V�<12	1H��ªтB�ٺU��x�<����o���'���I�4�0�CN�<��#�9�h�'�0.M�8�F�a�<q!G�
��Y�W-�j�j6MFe�<�'I��n� ��	�=�LТ0��b8��Dz� �!,�F��6!�Cah�a�բ?�B�#}�(�C��՚xA
���"�oO*B�	��@ik�HD1H� a�cJ�!,�>">q���	&#��L��"\@y�x#����=!�$��{:��FI͵
��qxP��=!�DEG��{�&`��{�I�v�!�� &a�j�<	0t��"�H�20Q�"O�=�a��
<�H�rk
�D�H�"O���ϒ�t�0�q*��aD5�"O6��rCK��<Y �I�EC�0�"O��`�@J�@���g��b&jX�'�'�`QϓT�0��N�*شQ!����b�ZU��t)Zv)�-���ۀ�A�?I8)���E?	v�@�|��PL1e
��⭛B�<�3���2D���x�[�i�'�Q?yY3`�A�(5*DG��"�2D� ��DW'�(X[gA�+�z���,D����
$��Ԋ*BJၬ+�娟� ��e�>E�H�&���|�f�5D���"�˘��#'+
_ɖ`
��/D�0�`JC
L�Ը��-���j| "��>!�V<N(�@�L;3b�SB���v�ȓ|�l�dk�`(L1��#S�!t����l�e3�"L�]k �Bp!f�ȓ�@x@
�'ߎi{Gū/BּExR�xr�2&}�� ��N�'g�a8mԓN�B�I�j1��y�m�=�Q8eѶ4zf�J���'͉��s��$��-B6D�����W������Op�D9���':^U��h0 q���>?�`��IZ�D"e��tEz�e�[WJ�Q��#/D�|!�hѽ]$�10�E�hi�ɓ@�MN~R�'6!���8O�:��4V-l��'�fx�Z4+��ek���~�ܼӏyr�'��q P
� ?dh#��v���}��'��$��S��PZ#,�8p<������3�!��-w�f�)�� *����L� G�L��Iq�'f��bL��!���B�zt��K�'�Iq�.�5�2���ƗxL(p�'����%	�� ���K�K�#!����'�F���j�=4��jp����\��'F��r%K*�����i�_���'��޹P�pp6��m���6�\��y�T?~�!��.b��z O�y2�M�a��b�+uX��\��y" H.w
-A0��$PL��f�֝���.�O�SA�R�x�Xb�cY�w��	x��'G�)̓cW�\�4�)�N�8��ԧ����;Z I���$o�Ѣ��=a0���!挠��A'� X"vNS�:��ȓn�\�7'�=T���"��Ҽ5���ȓnvRɒ��ܚX�D!�Fě$.#V��ȓM#>I�lԃ;y<q:�)�m�B��ȓkU�"b�{d�Ā��ՠ �D��^+܁�)M/J#6L %G�P�~��ȓR8ȭ��%&�fP�ѥ�(�|��?ό�	E�.2EAv��[���ȓ{@����`Ɖ7L��!+T Nm���x�����$� $�pёSa?���ȓsy�%Aq"�25,A��H�h�$���E�Z�UE�A���f�F�,}h��ȓ�Dj�Ǆ'G�l�4��e�e��7��Dj�J 9���C�#ՙ@�B ����o^�$%���ʖ)6�Յ�{#T�g�A2������?&n���<\�7�� D�9ghp�ȓ}�`-��)�⤊�$��t^p�ȓ}A��;�Զp�j�"��ߊ��ȓc�����ԑj�2 � ��qO\��ȓE V"�):t�d����@'n�ȝ��8�hBP��;�"I����%,��,��S�? �5��M�*q�9��6G���(�"O^-1�`Jʔ PV�3Q�Z�x�"O��PS�O���wIُfi4 �'"O$�IW	-Q��Xӈ�.OD�8"OLXfO5Ey�X8Gn�b���"O��2�J��ʤEa'N(9��t��"Ot a��ԯ��U��� 1�^ X"OhK�.W�R�v���Jr��TQ�"O0}�q�����)B�H��\s�"OJp��(J�@犅�4�2��t"O�1ЇE�	����򉖯>� �`"Od겦�T'D�q�Ի l,d��"O��+#ӶJ�T��RF+[n�F"O��zPECm�Y %E*=�<m�"O|�;���W��fe#� m1�"O�*��]	7&1
�CK.0�֌�q��+5�Ʃ��� w1�����
LRI3�nW���QV皒sL!�)N����&��r��1%  ?�!�B>_�}R�)�1_l� �a+ږk)!��/@�(d0N[���$Q� �!�D�a!�p��P,wH�<����
�!��Y����+�M��oC�i�VX9<�!�䝛{�vuKP$"d6��3�bˑw�!�$�q����E�:a)n9a�B�'�!��$�Z�X��/v"N QGB�4f�!�ė�b��Y�jA�E�1����!�d�F���d�L5�� S1 \(	�!�$Y�n���F'@����ϐ��!�䔵!�5B3K�'>�|�;�O�>�!�dܕn�D��f�S�T��y��!~1!���NA䏛3�rM�r�)�!��ç�z,�R�0��k���0s!�D��/�v<�j�4���rgU�td!�����Q� �<Y\ Q"Wr�!�$�+$�Q���R/N��)����!��1S�;D�,.�k�-B�(�!�$+�t��K�>�@�Z�J�"r�!�D�u/2�P��ͨ��X; �A�!�D
S��]�$�-4��i�WGD'Ki!�dG f�8,�D^�9�X3vT8>T!�D��8��(�J�1��H0�/"k!�KZ]�I���Zg�`��FY�Y!��,�I�d+��,��!OC�K!�$FJH��S��C��|�50!+!�$��p�pX`��
�N�H�ЗHċ^�!��,�>}P�	�z0�1��x�!�Ė;��{�R(Lh�S�g�^�!��P�P$�]It�޾Rś�F/.!��6<$�I9vJ@�R��d��'$;!�$5D	(Y�5'&~`tk���!�ބw<TzD*���z�$��W!��$ցKWN��$�����B"�!�ц?��I��J�{��ѓ�`TX�!���=k�x�����V$ ]`�O�N�!��1&���	%ðq���U��!�DV�]�&Xcu*��`!�,L+.9!�$- k�C���h�q�� ��*�!�dѹM�x�1O$3݈xnT�F!�G�����[ �0��M!�$<-�j�����/�t6��0FB�I!����c�YB�	�%
1~"B�:z� �"���(_���ՀY��B䉇J�f}9��ؼWD��F��:uʎC�I�:l`�!�M6y6�a���_�jC�)� JlI�`��葁k�1��m��"OLء�WN@Y%�
�X�t��"OB����t�HR�
�����`"O�uzQdX�)�j|c�K1+�ڌ�"O��k��s
�x��ބ7�B ��"O~���+�F�9bј~�J�S�"O"�H��H:����
��M���"O�Q;��-]9�]ڵɌ�
v:�%"O<��E	�9Oj�lÁ	T�B���"O6	[���l�h����3��@�"O��S�!��3$g@��s"O�\���R�,?�<A�H&6JJIH"O�����ĸv=���`0�O��S�!h���R��
f��H�fE�v�<�7gʋVQ��cwG�SW,�W�]r�<�u�_(|�-�q�	�����$�7�yb��)nf�;��φ��!cG�_(�yR�Z�`�N�;��J)�8�h�+�ybn�Uc�D�UD�Y��&c��'X��6CNL8�ĠB�yÜU�˅.)��!��,�O>��qKD"gr$h��D�F�^�[ӣ� �9Bf���?�c�L5�Q``�"��D�C��V�'"t�)1$LAd��R��X�~�a�bm�>�j`���N�$0!�D�eZ����f�>�����3UB�լ�C�LӘk�n1s@�S���[tBg�I�0N�T�Ԛ�I��G��x���-m�jyg���� � I�7� ���w����H�r�\R+�1O��$��a �E �]7����Ú�S�:& ?lO|P�2J�"_�ĳ�l��l+#�D�1�������_ǈX�lA6�~�WW���*f�Bc���⁘J���ɝ�?��G@�d�9���ȕT�@wj;ғR���о�<-"�CҐ(�$��O���d 3�1B6�px�P�LX$Ð!Z�2�4L��ʇ&-���t�E2Q>!#�&�W�$��eȯi�R�	p+."m�`X%���{Z��	�8�2Ҷ�^�@'�"��AB��w�{��"�ԫM��E�ÌC�I��G(*B4B��t�^9�,���Z��b�-rj�⃹�� y0��f�*yJ5�@���|�d
U�6��?�lZ'K��!��g�,q*��A�8.9��ۣI����$L�j��T��A�(
��t��o�'����0-Uow"pr�B�-A��9�/ùd@|�#Nb ��R�h�b���!̉*,f��A�E3X���L�q֬�"��J�EAT�k��D�ņ�49���"Ո�=�(O��3�T�n��|�%	6<����l�Y8�>�����!	0��5��KBaI�Ҿx�NiJ2@[�F���� �����C�*�F�#W$ ���$Ǆ�: ����pB��� X?K~Z���+�D�3Ĉ���t��~�]q�H�&��%�l�7�kю�Ag�o��%R��|��L�FM�~��l9�ɹ/�a8�M
���Y�'�;S{f�ˡ�نsٛFC�:�(�1�j�N2��J���q��ɏ�R{`����Y+�=��\G�x���쌌Rp0 �ҡX�#��0$WX�'����1��$X,8{���Qr��g�	�
CjA��� �. "EGIqV���`d�RH��0,��?ݬ;$�.�e��k�
� �ܜ�(�a�%B�&�B�E͍%Α�$i�΋w��C��Qj1ɂfFc�� ��ޥKP&u*���} j�""��D�I��& -���'"�+ ��$a��$IR$����9��I�?M�F��I*JXy�0?J͈'������((n BfGH�t��@'-L��L���B� a�	�jb�@�Fыq����#�~�
42q�1Xd� ��@�9��ǈ���2��?#<a&�W=L�:����X�"E��]d~��TN��LQ�����q�;_�<����C�j�,Ok�]�9�p���q��푣�Rw��}����v�ֱ�S	_���m�(�F��y2��s�����&k�8�2���%얕*/O��KQ�e���K.O�)a$�0��qt�=R d���ɟ!'��B�<,���W
�T��A��I�\�Ӱ/%� a�E_(	����!Q��+���z�0(+w��"!���%܃*J������Pp�-�XI���%��DI�L�rN����AFH��F<8Z����F
1a���eV�yb����\,�����*n�fe��"@/¼��=,^e�e�C�  |��'u՘C"��\��ƒ��ݺ|xAA�-O]��u�p*�(E�B�	k��ʤ��1U3���&�ۤ ���-�1m����|�A��5H�$˓��<y$��8D�԰��ɂ.K4���b�����R����mB"w��&�싃��s�Ԇ�	�]�Z�G/�-�` � ��C�I�\�^L��O�|�401�X<8�,ă�!V$+���2}P�����}�f5k���Z0!���v=���:�Z=�G�Ƌ/,!�2�`5�s?ok<��AEW�E2!�O�I�^�Zdk�  Z>u�0Øm!�� �����~
ΰXt���茩�Q��CP�E��h���&Z��q�D��KphЃ�f�$Ŵ��$B�_� ��	�8~�Z�j�&[4:\T���M�P�؀z�'�8�;Dl�eV���m�mGx��¶nim�H�s���rP���	Һ�Q0��?^����"O�Yys������%E?0ʼq2wϟ�4�:��N+nXV�S��yR����*笂�iz  eg��y��>*�a�vmE�k�tH�dE�y�b�7m�N��/�VO�y�`Ȏޞ�i�F�h�|xB����0>q�#��s�ެ*���]1	���8{`�Re�[�c��-��'v����$@	�d)T�����j��ռ@G�l��� J��?%���C���ä�1i�081d:D��(@g�Ujq2��2 ��`�)�� r�����%+�)�����dηz��y�G�\�PŠ��]y	!��%+��|ie�G�R}����Z�DIW(DI��U�I���^?.�}�QNM�?�dY2-K�LB�|r$�5.p8���K�!B��+VADD� y㷎K1i��y$��cF�"~ΓG���@5B��#��k�� F��0Ez��I�s�B�
��8D�<<@��۳6�q�g��P�
��CVx�)KC�9�Ob�æg����͂�*lZ�z �'q:%r����^
����10����U����>�8C�ɁY7��Y� !X����o6c����Dv�P#�Ӯ1��+Ŋ�=W6�܃����z8<B�#��8��Q#S��[a�º
�5`ɋ0%�=�O�G��O���UdބF!�Cw���"OfP��I�(� �r7@��lMY2�i�8U@%'W�`��p��GW�1�$u���U�<��D�%m�Q�*�&�?'�T�Y��D�%kRY�xj���c�<��H9�lh�d�����1�BPY�oa��@�!
P�}*��;}��1�瀔�
�,0�&Q\�<�c!�&/' #�A\r|�1/\?�t����	��H��	�
L$���L�W�M��Y9%�JC�6S� 8B�c�;x��cC8<��$#f>ܨ��a*�O.�ƭ�=w�,��p%�Vu���'pZx���m?)�iE�IOP�	gG�F"�ha$K�<�P��+![����a���'�K}2&�4>
\%3�'��@9F�
�Bc��5�� a����r���S�&�!R��P4*&	���6� �r��.D��R�΂�+ �A���%2�j�P�*��Y�&]�vQ
����tn�(W#�P��O��K҄����y�M�\.�@Js@��c�JLQ�B�Jڼ؉EB��14`�Z�"~�^p�paA��	vZ@!�-4�����
N��b���=<[��
R��128|�gڶ��s��&o&	3���hr�VR:@�
��X�����.��2��z lpӆÏ7j�>�zcBU1)�=*7��wh<!�S�c�F��f	$��!�#z�'�zx߆�0˲�����G,���V���Az+���!���W��iԃB�4��S@�]%��]A5J�C7<�ysj�<E��'5��
w���W�9�ĠK�F����'^D��/(X��MG
FG�0�'�X���b՛:�x�pd�'-8d���Z+t�RLR�")1w��<���9��
��ٲrH��"؃?����Kʔ*{4C�ɯI��]@Ú�C�&���
 :�#=a��W�k�����)[�a�b���5`����rD�
qF!�d�-p>�m�Vn�1z�	�6�vN!�F�'�Y(�gڸJ�NHY�BH)y%!�D��3Z�Ys�f�j����у!��_f�PU�&���G�Y��͇ʓ|!`Ep����@ �A��zDD�ȓw����t�9g�]+�$��OT�ȓx�H=�T��)�lx���W�m����)�lW�U�1�$1��JےNe�<�ȓ�,qv!��6`൉�o
�z줄ȓd� I� "��M�(�-W����S�? �DF�@f�̩CD�"z�L���"O��Jq�����������"OTU��`����C��\��"Or�����1nF�tsEI�!���"O¡i'c�;Ĥ QR��%%x��@�"O�)�Qk�!;V�Ժ' , r�})�"O詫�˥A8|�$O�g��m[�"O��X���[����3.��5"ONՃX�J�E[��M�@eL���"Ovy�$QJ��8�
��h<���""O�	���4#��A�7R�J}��"O�}��m�0X͙Pf4j���"F"O���bB<f�4�SOU�"B&I�s"O��6�ӏX{��4/	1M4��x�"O����6�����*pR!"Oڈ���Ǩ_�zp�u"�by�yB�"OD��']�a֠�lE\�fi�Ux5"O$(Q���]���8  "i8!�w"OJp���"}�D�Qu�ր< ��A"O�$(�aE�%X����.ѫQ'|�i2"OXAb�iƕ �L�ۦl_�
�z�"O���عM��
��1���"O>�QS�D�"�ib�]�j�d)�S"O�A#qeT��!�_|P�`"O�)R+̕*�\e��M�F�jI�v"Oi6ԇxB�0�C�Ȳ�+5"O�=*�@ؽhEH�y�(J����'"O"��P	�4D�D�����O����"O���(N��l����%o���"O��`f�6�\%0��)�D��"O�L�%h��R�>��P��&�U�"Ol �/9~�꒣�����S@"O`��
�$C*I#b�h0 �"O����</���h�ě�V�d	�"O�3$I	�Vz)�C˨{hU#`"O�Myf�̉l��݃eoB7zgX@ �"O<�N�Y:���6��X�'��\��ˇ	6t�8G�4.N�u��'�9ɒ�D�]�b���,ԁ,���`	�'���)� �]a�mZ@l�^U��C�';RY`�K� TL"��&G�����'1��G��x5�Xʐ/_+ْH��'Zr����.z����$R�'@qrLRf'�tW�L$��D��'��{Ҏ_�Vȹ�DңD#*�
�'S�l�M;*����&"�<r`-A
�'F����.�<uV��#A!�G����'Ex,�)فD�ZM��D7X���'��!��#��L �`��/��5@�'������8�p���'���
�'��Y)3�I`��1�2L��ؔ!
�'Ѩ�E� �L�qJ��0����'�-qC��h��ue��l�.��'h*��©˲r�p�*Vl��b���'Ґ�p���aK�X�f�#uc�ň�'��m�������:�a��>�a�'N��gN�"W�l �I��C�m
�'i��S�O �T8��X��,R��1�'?���R)v����%#��t2�'	>U��ȗ�iG��"��K%A�`�K	�'%��P�v�,�R7�Y(ne�0�'��Q��,��e�6KZ�[F�u��'�8��$`٩Se�Qp#&RV�ĺ�'v���d�p([U�,DL�1���� `��T C
M�-)�I�#؜�"O`�0ױ6P�Q�B�� i�@���"O���W���.4\%B�Ȓ;^3���C"OZx�T�[j�^H��lѠ,�}�@"O�@��Q�.�p�tl�

�ܚR"O�����sOd���,�4햔rU"OB}C ��3�Z�o��X,jE��.D�Ъ���(PR���K�1Se��B��2D���B�ߴ<�bX	@a̵'����'.D���/�|$��3tF͈}lʳ$/D��	*A�X�*X�6��d�t)!b D�H����N�mN��ZB)�ӡ�D��k�@���Ij�Z�ɖ�!�D=d��`��|m���,	�!��1����N�Aif���o!�dN�6����T�̭�6gĶ7\!�G���6/� 
����d�[=mM!�D�1&M����Ã4a���c�N6!�䓂i�-Q��3GP�X9F�"	O!�ĝb��q{bB�T����`�h(!�D �l֌92 ��%]V���@O (z!�ĊF���)�J_�L�p�Ɋdo!�ʕr��
Gi@�^$h3��W.fI!��PU���[��[�Ԍx�L7!��'v|��ҳ���w��I��ʐ:!��>3"9��oҹ(u��T+ښ!�䍝2̄�3s�@e���$IM�0!�� �p����k��Ȋ��#!�D��x��E+��t���ƌ�1O�|���F�p<�Q�! Ӟ)3�O�5t��6N{����Y  �f)�S�X�v$�Xj��*,���*�/�R<ɖ#�*jw�9��\�rP�b�H&�')d9pL��RE��/��20���
�9�m���!?�L �I	�e��
O�M�D�Ҝt��q��X�
&�숡��
!&�agI]�zy��:=j�% �Kt�Qr���^~q��O/8� �z�l�cQ<��$�fytݑe@V���I?3ȍkU�ϟKqPX��mP,m���a�U��d�E�?�����~��G/��lB�a�I�I� �³�C�
H���a%'օyҧ�)׆y ��a �:���)t�_-t�y��D�sn�ã	J�A��������=�c,ږۢ��	S�n��!`�.ѭ?æ�'�8� ��!\�u�r Z7,}��R8��	¥�w�6�kC>-��
K�k,=��'�<�;f�N)
�:qs1h̙S�yv��.XJ��� K���Ҵ	���e ���e$���0y�J�ቪf�A{�cZ-H�<�VY9v���0; ��r��DIv��� 9(�����:Qm����;j.d�kP?]ʴ�CХP�+�����R?�z��$��5
<xs5cA�a<}ʔCS�>&��� �@�Ҥ�
�1�����DwX�0�恧?�<�B�K�66U�	���N�H�2l�CJ�(P��@#3eP���ʦ�Z�k�8A[e��2�R�C�m�I�x�H�d����u��%�-O�VI��DL�։���wqr�)�흺�89�f�=�l���a2~��3KN3O�������E�>#B-Kj:e�D
�
k��pd�C1#и�X�FS�N�����ޟ��G7���I���ԡ����!�~A�a/�cҚ#>� !8�t*a�V��~2�ن���c5lJ�f�V��n//}Bb�*U=TĦhz&in�R����O�2��� �M
J��!e�u�:��v+s����|���;��5� ���ʉ��'63�"�[T�0I1�E��Ņȓ�|0xC#،=�ʕ ��l6V��'�l���n�-˘t��R��]y�^���,�wy��cL������	�(y����0?������8��ۻP�Α�f�/�ʼ�0�Δɺ˓r�
�K�C>8VJ�?q�͜��T��E�;Q k^�'/��CP��i���'����N �}�օ"7��A���#a ;0�`����h���Y���C��͉/<t���/��Z���zE�5�'��hx4N^�<��N~r2n�<{�f�06��!�~e�7dH�<I���Qb<MbDf�G����A}}�)R"1-N,¥�|�O*@0����OyR�
$���8t�˸e�J�ㆆ�yr�I�G��)Yc�ݰH�p�Xc�/��H�x�p3k��0<�6-�d�re�ҡ�v��Bs<�m��e��H���1-�e���z8Kf)(�� �����S�^v>�� >M�8��"O�km�;)w`�8@��;��SR"O��a��ß@�:|�ԏ_ y*��2U"ObD�'��&<���Ί�Z�*(	�"O.�a��Ҧ
���,�(��J&Z�P�p/Нe��A���#+� �f��;Z��-�rH�V�J���J!K5P��H�4D�e�t�ˤhd�H�V�D��"�'���*D��[�ܥ0�d.)lF�ҋ�M�Q|%�%hH��5��D��J<�:&<{��R/% ���'u��Jů��VM3�CU��)�pG[�P�.�qQjT5!:�)��<�(?
�rR@a� �ЧG�<q�h	����s�Ս��1o�<�I�<1�B��!���<٤�Aո�4N��,E1�*�w��(i��R�]���*.8D��B�%���i��G���ƓD�D�I�q*H�Q/�]FMDx�k��!4�p�ȋ&��L�B'��&U^4����>G�2�Z�"O"�"'�9�����,X������o*q��E���LȆ�S��yb�M�;��Y�%�Ö_�����Ć��y���*����@#ւ#�3 +_��y�(Y93l1 �@1��y��6,�L�;F��i'����M���p>��NK�W'Lx`�-��}�&�p1o�Z1N�#Bo� 8� \�/��qO?�	;GU �(�k<�~(�0L9< "=i ��+b���	I&#��`dX CpT�АE4}�"O�dE� �'�@�GFp�.���N�TD^��ۓ~�ؑ��jH*<�2�d�=u�LH�C��)|�<���KڱU!��/�.���4x�=xp�_?�O��B�;�h�������:�>�Z׀�-���Q�ʛ
f!�<);����k��g���s�	����r�J�R�'"}�'�n�#$��+���tj�!@�����'0�$��AF�f:2izDK�N��rߴE�6�('�ƤN�l����6W�.,`�	U�:�XЁp(�| a{rG�
?�2��џ�bp�ďZ�H�cB�+oG��25+"D���6�E�!B��C��
 ca�TbV�!��$��};0OZ���>�9�)(Ԙ#���.:^i�1�<D�hг��L<Z	�� ]�~m�# �>|�u���`�d�\����9� m3@阢~Nh�����!�D�;�<���� �h��� `��S:3}J�P�'�+oJ�)��A�$�98�ٳ
�$���ﾟ �`��*BY@cN�$ǜmR��*D��ʏ�a,����3D!;�C�>i1����h�)ד�:���'}��<�Q��<t����	�3�B�qG�O!h	*�ɛP�4��w�p��C7"O�\{'���>o�� d$���m�0ተl걁���bx���Z�d)j����@ƈĚ�aEb�t�<1T�G�����k�Z�p��$j5B�|�+
y�z��-O?牐䰫�hȺd�P��E�(��C�2��7	ʣ��x5g�*�h�ɟr��Z��Rt�ԅ�	�f2-i��� w"���Ɛk�^��$!>�`s��1� �9ՀOs}�P5��R�0h+gH2D���wL	�;H��F۔'��9�7�I�e��!�o� |�
�M'1(t�
��A� ��f�<��BI�^��� !�����uO_Z/���5L�@�)O?�ɍ:btʒm��6ʜ��"�<�C�I�+;��.K�X�*��bj����	�;�(��M��-�b��	�#�����!Rp���.�7&���$��BQԌ��d;<�񩥋�*M�&�VѴFq�$�
�'�zK��.\pG&�+	dj����pL 5�m2�'}�blc�o��Z.�b���|i����6�K�ہ5���*���)F���ȓ${��RH<=dD��ާ<�&����*�[S�T��:E�OxQ�̈́ȓ�4�����#�H�k�#L�<�ȓ(?J!�(���\j'H�eQ�0�ȓX�����e
��1Y�x�a�[�<� J��� �D����$%l;��A"O�а�,�_���B�Ï�[ =�S"ORċ	/H�ޔ�� �^%�	��"O�p9ՠ|7x�H�	*5�@"O����X
?��ɢL�4��)�"Oz���,U�'��`���&#�F�yD"Oޡ���J/�Azc�&���"O6�b�"�
A�<����?�,"O0A���eF����)(/�C�"O� ��R`@~\�iQ$2�TPb"ON���-Q4Ff���/Ԝx2&��"OT1�1�1 pq�τ�i�
��"O0b�lU�)��gD��l�!"O�=ŏ��h��ãJ�A���"O�a�E��>r�H�,�5���v"OxD�"
�6'�T���Q�<Z�"O4��c�E6N�@�hS�"R�eS�"O�|��`�C)"���\-h��j�"O���Q��	y$x�5�J!(e 9Q"O�P34�������o�B!T!��"O�Qi�@�$^|��7�� "O�X�ʙ��h���I�p�2"O �C�g�"p&2�xb�Z�~	N=)�"O�QAK	jR���KQ$n�H����B���P��*�
��${"d��v���r�n͍q!��[�鐖F�;�>�:��իe!�d԰[n��G%�� �܌�	&P!���9tw�(S�o	� �}Pτ�{O!�D�th2�*�����D���Y�a !��)Ld�`�dL�x�))�>Y!�'&R):�(XY���cI�_�!�
Z�r��D%N����"�GB�����JT�4IQ��O�� `$݉�1��H�:l�A��E��
R��O4��lZ�< �b��AE�0p�	FP��+��Oz���Q��G_��T�Y�{	��᧟1�Z��8O��%�װi;a�d���A�tW�7i�h$0b�@$X�p�	!�$�eh�5Y01$�-a<a��JF�Zl-��ګ|P��'�%]�ld��E֣t���7�x��M�ç%�>�2��?����̞W��z�i�,�M�'ᐽ%����bJ���$�N��p��aҝ5�@0�	
ud�I8���Sg&� DS��}J��1?q�P��/>ॣUNğo"l���E�x����^jMh#(�#�v�A�)9D��$օ4��~�mߌo��pˋ�!����Um���y2"Z5�ֽˠf��F���0�B��y2�����t)�d��E�H��#�y2�@�Ԁ-0#��1�x!wh-�y��\ъ��s�&�k6�ˎ�y����g&��WHUqT��베\2�y"�)oc�ۇ�e�pM*�����y���,>ת�
 l�r�j�y��[��yR%pna�B�rZ�iSgݺ�y�%����⋞ >1��+ �y�h��t�8�"~��s��y���=� Xz� r�~��p�
�y2�<��-Æ㏀c� %yQ@�:�y2�.'�xH8&�A \FLT� n�y�"O:8�B��t���R]*��%�[��yr��6%b2(L���sI�yB� 0�@��CKˠ��Q�I.�yb�Wr��QV���AΜ�Zf�N>�y���7c9V(��f�?���R�%�y"LмA�ұp�( �M�T��&�y��d�x% �6Q
������y������17���X~�P��F<�y��Wt�1
���z8�@�"V�y�a���Ib��O-m�i�5߻�y
� b5����//(�Tx�A]
|����"O���wc���ɑ��̔���p`"O@�3��f�|K�����x��"O\��3��0D�zd��p؀�B"O�@8'��i��Á��U ,cw"O�9�d"��Κ6����7"OΩ3Bl��.���������̀�"O��2���$p"D�6�.hc�幒"O�9K?����6oZS Ũ"Or��g������N�~k�L�"Ob�+�ʪ>��7OR�i��#�"OL}�Ì5v�Y�n�g|R�r�"O���`���$I@cM�W���"OjH���8��&��%=J�h��"O̋�R��8����J`�5+E"O��IƖ.)|��y����:U"O����\�f�|�j�"��e��8�"O()J�ǝG��I�qb��|��pu"O�Y"!�% P��FAD�]�ґ0C"O���C&:;v�����1�@�7"O���ϟ:��{goIxE:���"O��ʱC�
Mj��4.A���A�"O���jC!��e"�
<�Фu"O�� �E��.��`�5�.m8�<�$"O��!b04��{��L�X�!B�"O \A���9&R��P,$l�Ra�p"O>�A�ޜf������ 'T��)�5"O�q��U�D7��;�)�;e�l�:�"O~%��ѻR���y�	�9x"%A�"O��Q�CI��>Q�EȐ�&d"���"O�,�g/�/_���$[�qG8��"O��x`aǈ`�b}�ଐ�IS��X�"O����H�+�`�H�+H�c@�e�t"O`ಁ��?�6�
rMW��<�S0"OD���	b��#K�k����"O��Y��V�mҭˁ'	B�V���"O�P�&�QP�¢%C?F��e��"O8i9W`�-�l�7K�H��k@"O��`�� h ��)ܑ9&�8�"O�[�¨9����6)� |���"O�,:�MԨct���sg��\<��"O�YC�ҙN_�Dq��9T�y�V"O̬!t�p!3G�=���{��6j1!�$6�x(+�&��l�fpI�Bi!��Z!0t� �,=���!+0!򤍭4��B���A��k�
�1#!�Ԥl�V<i�N��f�Pq p"!�oS�г�!s�@����!�$ޅP���b��a�D����*�!�$̞����Pt �����B��"O ��Ю��dvƕP$��7�aj2"OV�ۡ!T���i",^�8�P�"O���$�*e(�雧=��@�q"O�PD��;�tH`W���$��e#"OvX�n��]�V���P�`$S�"O6�z�@�B��{� B�BZ�dJ4"O^�˂��<t�&�;��ȩuK	q"OИ�F#�^��wE�_�!�W"Ofђ0���� `�ù$�~��&"Of\�4�^=6�
���LF-BvP�W"Ov ��/]�8�+�(,�3�"OT4륂�c�@�)��5N�D"O��R�Nݲ>tX�4B��Sd�X�"O���a_9QYn�`��j F�Xq"O� ��*�@1^�q�1�ڡҲt��"Ot�aWÐ�u�YV�)�8E�"Ox��'ҟ5�!�Uk�<�.�h$"O��P�ա6��X;Ѩ�whD	b"Oj�I�&+P��H��J7#ZJ�"�"O8=�WM!"!����fVPM�)"S"O>]�G����`�$2=~�#4"OĈ23C� ��I3"Ï�3&�;"OLI�A
�?2��"���!E�-�f"O&@��O�8���Z�E6OЭ��"O��j��X�sp@{FDK-���"O0�6�S#M��]5!Ҳd�2@y�"O���&�ƞi���� �7�� с"O�4U-9q�u�ꖃ3�|�"Ot��K�JM
�@!��(L
hI�"O<��F �EBF�B�'@����1"O�t���Đ1W�$2��h{�$�f"O�u��S�\}@�� ��Ug��6"O���c�� � c#O�]N�� "Ou��T�A����1��l:2�`"O�h�e K�]tHDZ�,��	&0!��"O�E����2ZD�z��ɖ)$� ;D"O�鐇�õIQ�T
X�-�)��"O
��c[�+�Y�*[8 �P��"OD]sO�sŮtR�һ<� ��"O�L�`���_�	��c���d$k2"OĐ)@I+Y�i�)�$�"D�"O]��B�wt,��]bb��g"O�:�i��Q���S�Y[R�B"O�U����8i�:�%��L���"O܉ʶ�I���OƝnUx�Q�-=D��(dDۃLACdH�7f���v�9D�lp"l
�>��Ci�<&T�a�*D�T*�"P�O���	B���W����4&D���A�95��<Pe��!��
O(D�بg	6	a���L�a��݂�
*D��z�^\}������o�(�sd##D��+m�@��0Rۼ�>���+?D�(�G'��$�,Yj�ƕ�-�(�r�m;D� RD�o�|�w��NM�s��yr���s��qs�A���ӣT��y��A�OzRu�YjFhG
�n�FŅ�-��(S�{bu�b[���ȓb5(�RtDH�y%pYCr	X9Vc:����~9s��Ec��Q�dcл^|-��bz,�q���P+&i��5������l�jr�r1��U��P��P�@MY6`�ǲ��=8o`	��3zH�Eˋ${��c�,k�1��cW�m�Q�1���4ټ�#��c�<��Ȅ
�}��.a��x�D\�<��b��EᒌK.5��E� ��a�<�A�E�oʫ�N!��"�_�<��)�$!��¤�&
�,�%��Y�<�4"�0q�P��-�^�í_J�<��ɛ�H�V|��i��C*�P�F�B�<�Q��,4:*�-�$B�����y�<i%'�M��;��M;$�fTP��Fq�<���D�(���-��`�j�{
�o�<� e	@�P��y(�,��͞'�yI/p��!iw�ƞ �`����y�:w�b�b%ѾB�J �����y� V�|��\(�%��<x�(�%�yrF��euH�ᅭD�/�Dh�a���y
� �br�Z9\��
e��'��"O8���d�gfʩ`1�� M�N���"O����oD13��Y�%��%�h��"O� h֦�8-��E�ʃT��$"O 5��@Ԧ;avL; *�s�z6�/D��{��V�s	����杪/��#p-#D�h����LA �I�j�M�!"� D��q���}o��hڠrΊ��`?D� ?nJ�AmX�-txl1�>D���1-�5n�J$	�W�n��U*v@?D��HjB-X��Bc�eT�#D�"D�PavJQ�*8bR�Pu�q0`N D��S��'%��q�C���6(h7';D���s���M�J�c����fZic�E>D���ǂ��H��	�/��Ӊ:D�\�a�Y9\������i��bm%D�0dC&$d�MC��[�s�&e��?D��GFU 4Vvt�@%DT@�X�h3D��2��-o��c`�ȓ-� qH�0D�h(U���_fR����
T3�@�g�/D���I�/Z�![�BƆJw� i�E.D��A�K�\��{ǀ�-U�8	c*D�8I�i�#�4�;�ֲY�z<QcJ)D��[Dk�Q�r��"��tDL�b�%D��s�M�"E ��Q�� G0q��!D�|X�홋PZ�@��O{�ȹIe$D�40�W]�@����δ!ń ��� D�����>�ڨ�b_*Y�dܱ#�3D����Y��$-A"X'y�BE2D������*�L�B4c�	e�k�d/D�<C��R
��u��L���K�.D��Rro�{(��p���c��hb��.D� �5S�3��;�(�9�L��g!,D�D(�㞾i��4`�%#!0�)�d*D� �ũX���Kc�~U�����"D�DhP��	��eX�@J,Q��9�� D���� �:n���X�-� ]8�PӉ+D��G!�$G�h�P�MFSw����%D���a�	�H`F͂�!T�<��A>D�`C�@��k��@Al�x�%"D��9��( ���qV,�0�8��#!D�@H�l^�&�2�c
�/6��A�<D��G��eYY�b_/3qȨS�9D��x'��(h���{7	�)fc�	�d=D��������$
cD�v���F�<D�숤e� ��h�GX�}�B�	:D� )�80 F<�%iA�!x��=D��^�#���66�[ǈ�,#>zC䉆Yu��r�kլ6�M��#E�pC�I#���s"C�7��*����.C�	Q�†�N89�X �W�B�	�5��z#�[V��u!�II/L�B�	0=��;R ��Q��ͣfH�2����"#�&Z�\�)�S���ڦQ��@�&D:x����-j\��n�Xm��'���d�g�	#xPr���e^�9h�!ؕ��&d�Ѝ�ۄ<=(Y���ܙn���ku,_9O7�jiλB4h��+f4���@C�b�%j�'%��l��Č3�H���$.9��Y�{��X�F!Y$Ib����:lO&d9�"��jI<hSD&lj"�[җ>�'�F@iӶ�Ă��e�O����i'(����Y^��*�@͌))���'��1�-�Mc��?�����|�ܴD^�����mil�K���*nT�I���Y�a���4��}��� ]�Ό��@�2�MC �Z�?��+�5�ʭ���љKGx��f`B�hn��T���OܒOV�$�O�O�)*F�	�W��]`B�[1@�m��a�eH<!��M7x���3�D�>�����	Byr�|��c�X�d�<'�T?t�� Ȩ��ƓS�%I,��>h���ڟ(�IV�i>��	�6�� ���j��A
A"Q@�+8YN�0P�l.lO��{čF.VQ@��[�wސ횱�����$�H�/��� ��2-���5ړVw8���䟐i�lJ0^��pbP��Dp,�Њ:>Q� �	fy�'��f�O����K�Z�P�SGD�R�ɻ	�'J�����B�#�kV0��dk4y	m�Ҧ��������4=��Ub6�i�[�,�OA��
Ѫ]��l��� �Q8"���'�r�'��CB�|b�'��O�pESeT�e�4�c�̕0�%��}��1vi�����e
Q>aDD>��]�6mE}?�9�M?�	w����O@����a��E�UB��btX�aS�Q���v�d�O��=�]�wr�xJ��D8�r�̇������Ħ��A}Rd�C0����$n`&`xAΤ>ET��d�^��m�IIyʟ:���O �d~�<�PDC]�.���,�5��8C��P�۟� Q��|b���h�|IʒAU'r�FD*V%=v�	l�'x8�,�wh���J��Y�L!���<�X��vmh��	��?���G�	&S���O��O'c�p��e�2���o(
x��H2>��=�O�<ڒ��*q������D�������)۴��O����ip�t�t�Ӥd�>�s)[�<��'��(�Ӿ���O��=�4��6"[�����O<?,�`Bk9E�%��/�u؟��Aظj����"���S�fӺ���F-�`�R:\O �s�\7[-�	%�Ƈ*�,I r�iu
�C���?Ya�x��'ur�x��D�^܀���5���(��	fX�h � �eAL�"bD_a,���� `6-9�DE��S�	Ɵ���RD �  �