MPQ    ��    h�  h                                                                                 �;I=2^
�nc���nS~���R<K�їn���R��8�Yڧ۝��s��y�X�?� Z��O��nBU�Se2�lB��j!�m	+�]�[p��U�k$I��]w��_�a�A�C����wlbc��0�V"��g$�z�?���ӑ�L�2��d@�;/%�e�`Ywr�c_���{F*��{��J��Z��_����V�<O�i���Ӝ3��@ֲ�i���Tx���W���M�u��C֩�b��q�w]��B�vܒtӆW���gz�JAS�C8�u�7~���ۙ��.͖����.�X�$Bot��<r0,X����4�ϾN���>A�����I��R�5Ѳ"�0p�u;[^�UL��h�0�+�;����V����9���;n�./�u�F"L�JJJ(Sb��\����Rsˊ��4ɀ/|yX�[�Z	�������U���6Gפ��z���6��_��c.0}�l����a�FT��y�M��p)�$J`�"(�:�>|�9zo�x�K4�\����X��0���2a���n�)�h�]�?��˿����h��۴97m�y�	�D��;�"e�0��Qd&m�
���g�/
�ԩ�T��G��#h�r3��0;&�FG�
�ە��\&Y�h�E��V��~��R@�*��oA%�fލ:�7Nt�O���)z��E�T��+���?ʺ��kN,v��#����J��L͘t�B�(:��,�y1ܰ�@)ռ��%�V�<@�����?���a��H�W��;�L����WT�`��7����W�������_�Ka0��3"�s��f���z󺘃�m��A	�y�Ҁ���$.����}	�c#B]������v���$��ʦ�o��Ow9�g�_�-5�wb����Y�|5'�3�o���w��+��P'E
[��oߨ�2֩n*Hn�q�w6 ;X��|�tf֔��<۵�u��~�֘�ƽ�͹��\��oZ���r/�ƴכ�����9Y�>se����h���j�7�2�E����w�F��C��y���<�oT�b>�E�|j���^�GV�$��E���x�4O�2Ϙ�JZ��]C��y[�٧��hd�@��B�5�ő#`�\OE��x�r�x��K��d�G4#b���T����O��.��a�:}u���
8�"��3d�W?��3G������@�������H͒�4i	��x����E@����P����&�'V�f ,�+��HL�E9[��U�����F2����L<�a/�RY��zZ�Ƹ�M[��c��?�e�%��A��3P� ��	��f�;�(�d�{��j�Q`�$x\I4��.i��W-Q�A�=�]����
k�xj鄎�&EV2����ȌF�����}�H��U(W
�� �>/u� ��XsةF��DY�q�4R�۶RC�鐶˫��-ْޗ��U����C�IŊ����
���{Rՠ�����sUct���# �~���~�f��a�K=�>�v?�R��14c��~��7���L_%l�Q�j63
����rc�����&E���U��x��z7�-�+��P���w�V� ��'>�,�|#���UVNB��%�O�{Q|f�,����Z��k�Dt��B��EZ1�(�͏#�Rk������x7{�P�;�R�`���ܡ��d���.i*)�3ш�f���W`@&Ml1d��輜,7>�k�q��8�hiNA� �2�2f�t�$�g�ʏCFA���rmP!y�(���*����{��y�7�j�UV���z�`�yjӛ��/3�\�_��<��ؔ��12R�I\��e����V�mǿ
��L���?3v�3j���(� �w��>��Q2`C�b�H9Iv	��8��{� �S7��z*So%Bl�,��}w`!#pD=��������ޝ�C�$zi���r���B3b @2�Q���F���	��)Xg`8$[R�Dk'N�-OD�����T�z3㮝�.��ʍD/����s+���nN�D��
ɢet���0�O;��6�9�1�f2��9}���^��e�>b�=����H��&�f��[BO{��Z܆ȸL�r}mp�W�-���������#|��}z��ŒA.��-����ǣ�-��`�G�Ј����m�=�6�ٻ0���P�fT^�� \���U3�e��D&^��Ӝ �����ov�Q㩧�"ŹDkT��R}'_j�p~�6Ɵpb{�R�ʗ���*NH` m�b漓�b������ D>h�M��A�i����rg"��66�2t�i�	�>N�b����X�{`i,�xz*;SB_���wx�Se���sS`D�K8u<�:�v��Z��?΀����)�����p����0y\?j��y L4Ӭ�b��&q�-Y}"�uE���F����Y�\�D�O��3+1��zآ8f���Ͳ�3��w�!a��Op �)���J��HUR����$��E�$کl|�><���=1t)�M{'�����\k�0�4��I'��\�Rlt9����6�a�͋�r99��QHw��R�^�F א����g�lU������pT,���pA�	sxd%����$��L�G�'Z�C0t��[�*������������Cuu�zAl� *��N�6�h��`(xkg=R�q��qė�=�,�������y���ҹj������G���S��@�/&��3�"�.��������lcM��馅_�JC5vCXgW����C4�(��;n�E���������l��N�ռB]d��b���z�\����݋g��*Pڈ�:�=fp���r�%%�������sowN�	���
����	�wI��F?���&LܖX^,�ȭ�ܿ<K{�:L�9Rx�<އ��tc������p�`pH˶J�	��&��V���&��k�܍%�.�P��DO�C��Ľ\� �2;6�!i�dT�����yn*C�wlbj�_���;��!�n�AHً� �`�"E!���RHq�I���h�&���? X������'A���,�'4e㯌���|�5A��]��3�!�����UD�K�7��M���b��� 3�b�;���t���
*I��bXH�ւ�Kn�A0�'��������ί3�CU%dIW
�/��{�5� �� ���˺��N�I�q���C:t����Ռ���aҬ��.��!�0g����4�Fa+�DCF{����XmQ�:!d�(�q<����۾�Jbo��R�N����eQ��v���@�i�5�Ö�x���#��}�0��X�]i����1��H�R�H����,S�3����|~�R��X������$ɉQ��ߥ�t�j�r�j���2�I��j���߿���pP�*ˊ�4�]5�k��O����^�$��6t�ϩp+��Z����Vh`��?�C�\n{�h���V�*L �RJ�r9b� ����_�s>1s0P�89;��,X���Z��]�C����q��6B��-I쐡��w�_8��.�$l
�J��	�FO�9y�M�+��$e�"��:�#7|�D�o��K/g��m<Xl�S0��2���I�6�����i �P��,��h{����l]7�)�o,DD��� +�Qv?gm]QF�х����/��gTK��G�N�#cEfr��0��aP�
<:��PYYPJhKdy�Q�/~3]@]oz��c��A�h�Fz�t�n���)�>�E�<��F�!Һ���}�,�������JEw�%�-� �G��E1	s@�4���xiVB��G������_�Ŷ#b�3�-LW���u<>�(���L�Ґq���J������"|��!�Q���r[mr��	ݎmEs���.Y���8�[c>���'�S��P��Q�$0�F���٪���"���H{��򏬚��xܔ���֫.R��ʠ��eА�w���E�Y�ys�ͷ�n%]Hx[��2v�;sE���f����w�(��r~�I�!�U�td \���Z"�r
�Y�L�P�I���{ҙ}ݐm�h��,j�>`��a�^��Fё4ޞ%�4���4eo��>��E|�l���ZmV�e���,����04jf22J�J5"_�����4[����p��h��@��qB�c���\�^�������p����x>m���G��_�WT�u��J.��a'�}0�7S
�_I"h��d&�W���3B�4�O��@�T9�I�#*��mw�iD�Ax��W�@xԎڝPP���A� ��
�A�L,4f��g��9��U��J�Y���:x���<�,q/+�k���Z6TT��h𢳳�ӣ� T�A2�TPA���ZfC��(j(���>7��4�,��_?�\�g�)��M{�-�X��		���4Z�>�@��!t2%��d�ȧW��Z��}�s(��(�0)����>��2 �+s��~�����ܬ/�4�~8�M������Ҕ�Yb��0���X���@��!P
^9�6���0�U>9q�%�� �e~��٠�صg�KXgY�~u}v.������y"[��z���l��]j�ަ���ĭ�طM龓!6��ߠIxɭ�z��-�qL�+���k �V�ٞ�/c���t�#�����Np��`(�eff����A2���D�X�BZ�1��c ��N�k�I��!�x�7�P�Rj8��N��9E�4�y.dGBƎ�ň!���9X�W��E&(��d�N��7�>�Sq�٭�#<`\�Ly�o2A	�t!��g7��CA��0�P��O(�**9��Vg|yOu �(�P�����`cbӶ��/���:�<4�b�`��-�I�	�e�c��0�����
�,�L�m�?�3W��4jG��(Ά� 8��򬫵T�Qm��`�P��C�vdz�8�r�;ѹ���U�3�1l���x!�!~Y�=_���A�`p�4�$�c�A��n�BfG� ����l2���+�䬗)�l�8���?�aN�l���x��<d����x '�'۔Dʙj��~7�La�	���wZ��!3������V���0��,n��<���y���-��MHe�	'�c���ЎC%w&Z'��X��[]�A�%k��.�ĭ�?�o�(K��#�c� �|� �zh�d�O<�h�?�j���d�	а��Z����y��=����w
�>fO���A���)3�i�]�6^�`��;'+�Sh�v������t<�T�ӬR���j��*�N����{��U��F���Њ`;Gbaځu/��4A���p�>c.��oTt�$�x�[_g��A6Oet�ܘ̤��N��B��i�6��,�(|*��B:#�< w���S`���1�=`��x8���:Qu��_(c�zW���O�����p��s�K��?��T��Log����&l:IYؐEu ��ַ�0^��}�\2��Oes�+,uzxq�8!L��)VI��R�a�R�p��������H�λ �w5�l枿�$_i|^����<1��M�U���������wU�40��'�� �sRǎ�K��Q�i�HL�M޼9�OH�7.���~^LL� ������\�w��q?��[�T�-��k��	��c%�%ش�������"9�6	���8;��w�*|��|����t��P�>uP��|X; �p��5�6�.$��#k�p���g�L@L�x�],8�V��p��Ԙ���������?ݢ����C�9קx?���%}�����d�3�4�`�AM[�T�������v>�h��Э�COb�T�En���6������ǹ����w �d9�b��z����Y���x拫���&�����p��rx��%n��O1�e8N����p\ߨG�D$h�wď0F�'��_��1�I^'����� �i;7<f�:ǉRS��wR�Q�kc�زR�pBJLH5�J�����?��n6�?P�&���7�w��i�� �NO<��C{\�`m���S6��Gi��c��7�S�* Hl���_2�T;�u��1yH�) �B�"�F�ի'�qC@b�xQ��!,�
�X��}���'�1C�r�4�^�K��w��A@��]eD[��٨�n�M�'@D�Ѿ7n��'bH ��V�`�����I�fX� �}�xn݌�0EԶ��ef�CC*Ί�W~��d�z�*��o�5oBt����Nh���˥����~F:�\��O����E?�'���	��!W�;0����a�F������{��ӟ����c�S<�7����Yt����i걚6�x�����>�=�v�þY1^�Aй����"�g!�]DW���b$Sɕ�M����&���|S�C�k߭~��N�Q6�.ZT��KY���W�)Ht�e2r&���G\̄�^�������g�+��E�􂯅5�Djъ����^���喸�C�+ɽj���VC�єG���z�nv���+ڣ��BL��J��b�O2�������s���]�����X��tZ�t�C�0���jB6=WΈ�~�\U��	_�gc.�f�lE��ė1�FJ�yz"���V$�:"6_:�S�|(po~gK*eN�: X'&�0�DK2W�-�${����ug?������h6�<�꿧7c����WDKS��X%&�AQ�:Hm�F����%����T��G8"*#^�er� �0��	|y�
�T*��IY��h�Y�L�~�nG@쮳xa���C(`Y��t!��	�)0��ERDl�a���5o�ꔯ�,�M�Y����.J��C���H�g�uٕ�!�1R�x@_�m���V����׋,ʠ��2������n"�L��7�����;��є���MT§7DZ�D����ݟI"_�b���@�������mM��	(��3��|[0.�$v��f�cYN��<׎�٣̌��$�������TT���Մc�y�m4C�����?�ϲBޫ)���%J:�~:����EE�����32�h�]n ���/���Պ;����rQf�����E���U�~嶖�|�B�/O�\�=Z��-r���M5�뮭�}�Z�����(R�h��j��0;���<����ZF�'@��z����L�oJ	�>_;U|�R�Ԕ�V��e����o`4�iS2�EJJX͌��,�[����U�hںS@�oB-�������3��6�����(�ux�����G*�:��T}��y9.�U�a�}��<"�
��L"C�da�Wu)3={5����@��������HY�i��x3^N�;У�_1XP	��\3��k��,T\t�~@:	��9�PUUkX���J�<c0�}$w<�_�/�gV��Z�PV���#P�5GΥ�6lAm5�P����]f��9(%훱�c����\q��&\�1�$Q��~	-�v0�sX$��9����� �|���2�/�����w��L�}v� c"(�w���8>�u G��s�Z��&�������4�0�H�,�F��A���(Œ�L�Av�:��ގ���a
w���g,�Ͽ�}e�Ug�`B F�g~�m�4{��p��KsD<����v���=(��� �th����� tl���j,�/�^I_�� ·�FۓG;�u3���M9x�`�z-)�-�W��fs���rV{�Yʰ�;�#���N� ˌ�˴䱘�f�Z�����L�CD��B��Z�mߜ��F�Y��k����|9�x�XP�R�/�w5j�t�����._����i��R��T��W��&p�d����i>�["qS�B��.�wA�-�2F�t\��g�i�C<�����P�T>(&AC*�%�1O�y�X��r�Kr�P�`k
���,/)�����<o�`��8�(RI�gex�P�K�T�c�|
�jGL"g�?STP�Rj�Ew(��� S�Xmf��<�Q��`y��>Sv�X�8hu�V��I ��02��#�l,���s�!�b�=��(���]���r�$�}��D!�{AB�{F ���؇���<����r)Α�8Z�3�:8N6�s��f����pގ�S�O�b�De��ǩ�����ă����[R��t���ő��l���'d4��؄��Ą���e��[���C��>��&�����[x�����~ģ�����V��#�$�~Ĕ�uw$|�n�z��/���iԣ:����ۻ��@��	"���=m��1�)�3�JfJ@.�;�0�u��3�j��s�^���v�o��!�v���]���/TT��(Rs��j��欉;��*r{����M�g��s�`VAZb�Pt�o���, �>^����6�߻G�@g{�6���tpn�?�vN��ɁD�ڝ�*,��e*®B]��w�fwO#S[�,��ħ`�*8���:̓��:��� ��- �z�$�aZ�pQR��f�=?`u�/*�L�,����&g�Y3�u�(��H��+���\m�9O C+'}�z�*28�0�a��-t�a�p6�U�8�� ��H���T_��@�yYE$P4z|������1*(�M�PA��jP�Rv��R�4k��'��$���R"ɩ�l�l:��,��(ΐ9Y��HG����~�^��B M����9��m����QrTb���fN	)y�%g�I��f�����~�q
��ya�ֳ]*y7��7ҩ��r��yfu+�
�dY `k��;U6V7��k�k����g��'��Գv,��q��B+�/�h�Hu�/�������,�~�&�B�г�M��S�qt>�N\G�ۑ�M6�������"v9i�h6�Cj��ϼ�n�_y�q�.L�H��߹>S��2�xdT�ybz9zk̓�����<����>�1���p�g5r�\%I����` Щz�N}{���D4��6?��w?^nF�.�7����9�^"!�U�$�R<��:B��R.eh����앚c�v䲭RXp�S�HP-�J�P�c�5� ��ڦ+&�-*��@����k���O���h�(\�δU��6���itm�?H�+5Nd*�i(l�T�_��n;�5E�$��HO�x �D�";��Ն4q~Ю��m����a�XN,�� �X'7�g��E4��p���r�A�.] �������r�Dxb7�����Mb�W� ��B�qF��j�ޭ�֋I��XTٜ�x��n8�10 ��������eUj��>d�N�%:�ʇ|5*��72~��$�ڦ�<������ �:*K�
�8�ʄҢ����c!�t�0��ܮF�`��{�r��N�s��D�䞎I< ������� q�<����Dz���L����y�n�eù<=����t���g���	�]O*�'Vk�#��HM��O�{�0S�s%���~�x��4�����ĉ�?b��U�ztـ�r�Gs�t�̿�b����'K�O+���@Ā`���*O�5b=���U�F��^�"����y�E�-+���V�ꔂ7��y��nq\��нw��L6�J��bg������Xs�YO���`��XQ�Zz-���k0`��FK68�=��1����_.]�.�vl�/��2y!FEK�yռ蕡z�$���"�v�:b�|c��o�0�K%k���#X�(0��u2����u��Y���V�Ұ��h�/�3�7޶7l�D����a!)Q,V�m�>��"8���e<�T�t�G��#Y�rDg�0l����T
2�f�Z�Y��h���G�[~��@ӈǳ"���S:��i�^-t�����)�W�ElG�|�Ұq��ok,'�D�H����UJ����P��c�v��ɕ��1��@�Sھ�~�V�����H�G�9�U�h��>g����L��+�� �X�O�٬����7������bk����"����/��8|t�	�}m(�	S�{T�wO`.���E�ct�������B�ǁ$f��LC�`���a��~�����%��o�
��M�=�$F���b�9/.�p.��vE��� ���kn�p.$�ȨUF;���fg2z��*J�F��~���׻O��Y>\��ZMLr�H������Ƀx���O����h�=�j��Ҙ��7�Ȕ?�F��'�T�]�����o�D>:��|Y��/֠V�G5�VM��D4��|2@̗J�ˌ���[�]J�&!{h��h@�}�B��j�������+�-ڏ{�����x��t�*��G�Y6aTQ�� ��.�7a�>G}�=&=��
x�"7xd���W��38(��8�@O�����o��#[Yi��{x�B��6H���2P�k�w���x���u,������?�9l(�UY����ⷫ��X|�<2��/a"��4Z�ΫX��س���䥶9UA���PwK���6f��N(������|ё��	���[\�����-����ú�;�қ��t�G�2!2�},���E���<�P�Q}Q�^��4((ޭ��N�>@�� Us)� �t��ս��"$�4#Z�C��Cg��F�CC�OWy����u�+�u���
���Ȭ"���ь����U�"��( �@"~���u��+�K�A�t��v�m~�x��4�ʎoΗ�H�f�}q2l �ej����9�q�#�����x��Ѓ�����x�3�z�_�-�]>ɡ4ء�Vv�0��9��]""#�v;|y�Nӱ��֗��L��f�!���^ӵa6DŊ�B�bZ���٧A���Kk�M���
�xhP��R`G�R<���7�j(.Z���Df?��ڥ�o66W�'�&�!^d<	��m�g>߃�q����A��}�o�2��,t��:gmieC7�	��	&PR�p(A��* 
v�Wy�[��;�>F0����d`ٓp��X/�8R��U~<��Ҕ�e#��Im:ge3�E�f���m
b�IL]��?�a�U�j��(D�� n���?Q��ENQ�"`���962vW�8#旫q�i�D���d S�l�0�nի!4��=�5d�C���V�X��Ѭ$+��wƬ�v�<Bи >\آ�&ڷ�x���])	�8���5��N�K6uiy���{����.j��[?D )e������y��(�բ֢�OW� �����"zeC���?[������d?em� 7���9�l&@�ε�[�x����Yz'�#q�A�������e�0|�az^+'���F�޶�Ǡ�J��2��q� �I��$s��o�A=H�F�lf��<�fE� ��$k�0cI30�J�S;�^����+����v�a��1Y��vT
-R��Xj]6��ĭ��Ao�{�z�ʨ���[6|`q[=bWub+)���qB�ǯu>YT��%9���	[�E�g�#�6Ǟ�tG#�����N�L-��󫝬�!,�7*���B�τ�iAw�CSV鯢��`ue_8�m�:G���$]�������u�b����pAm�k�?��.
��L����3Fr&b�4Y�͠uv����&��%k\��IO��N+""z.J8�5#B�?2����a>�p����[��H��E�6��+e��T�$�)�|������1�W�MHk��v��+��-��4���'T����R}#��>��p��>-��޴9��GH��$��DN^7Q ���,���۾��>�8h�T���a��	�)�%"}?�-*�}#�����+W����>*�������n�F[�u���+ �����bc6�
��=�k�����2���%��Cb,n��4���pЌJyÊ5N���n�����kڳ�
3j��,\�i;�VT�M���W7���v4�?h�k�#�cC�֭�J�_ne>��T��C0��l�������ldob�b�[#zF4ɼ�hi���k��$�ڙ�=�n�p��rn��%$�����C�D��Nxd��&M	����Z^w�L�F�즄r2�g�^�c��?���X<�}B:��R	�є�:����c��,���p�}PHk��J�f�>��;ms�u�&�w��ɼ�_���6(�O2R�C��\@u$��v�6� i�!���~�b��h�*��l��_hE!;�A��HH
�� �f�"��>�a1�q��/����b"����X	�B��g'�rX���K4�O����m�A�C�]�������d�7��dDA>z7Q��pb��X dc���)`��߭��I?�)X��B�s�&n��80��£���9F_�@-�Yd"�� �%>5�%Y�R�b�DJځ��w��B�w렢a:��z�śd�)n2������
!�f[08I����Fr�u�U{����dצ���ًS<�`���#e�[���֪����,>̲d]������:uô??��/�c����]�]�f��bi����CVY�S�64IS��D�af�~^;F��R�d���]�ɚW��1t��Hr��Oa����;A3�Ћ��ɨ��t�{�@��8�5=Vr� A���i!^�Q��G�� �2+��b��V�KӔ�v����nlV>��,޽2�LQ{�J�bB#�Ha��D��s���I��{\X08&Z��f�1���6�BC�63W��>���*���_�r.��fl������VF@��y0w�\��$��Q"�:=|�&�oU�K ����X�')0�t�2M��ڐ��TϦ���e�ç�=��h�Ǧ� �T7Y��Ga_D�5՜�G���Q���m��3�"���P�@�wT� �Gn)�#Tzr��0'-0�+p
�M�5�Y
�fh�"�B/�~Dq�@�Eĳ= "+Y���c� `tWt����b)��Eȳ&ԗ5��+���Js?,b����m��rJV��#�~�-�0f��;1��@����1kVS�x<��bԚ�Ѓ춴b��,L(����qM�x
����C;?�]�`�T������P"U7�R���SgZ��� m�	��� �rc�.j+s�iDRc��o��Ob�wK��fD$���+�ٻ�o�S�\��^߂c�T�x�*�E� ���������i��C3�0֒�MEvR�[���n\��8��c�;Ī��h&�fB�o�(0���Y~��2�|ͥ�\&"iZ�r��3��%�!���s�LҪ\Ɛ��h��j|�x��d�1S��/�)F³�ޯ���e��Xo@�k>��|V���îV�� �����K4�ϭ2�r�J�#Z�IHbZ�[�ɸ���hPH"@��B���s�D�3ؠȝ�v��ުxo�
�E	6G U���T��笻�.�9�a8�l}a��X�M
�"���d��W�<,33���`��@
�L��"�A���|0i�?7xiG�1��@-P��NÒ��1�҆R,�-������9���U�f@��H2�2�3��<m&�/�����*ZG�g�����cA�+�祑\�A�qPWx���fT��(�3ٛ�����aƽ׀{%\�6��o^�;-=����D��z�}�v�h	�U3J���26�d����JJ��U},��@'(�d����
>�� �WsDZ���񞰌�]Ί4���>w��/�*�^�ђʁ���W�X�ߵw󻎑Y
-�p�g��΢s0U�G���dC |�~�ÿ����8�K�^Z��V�v�=-���^��l�jT����_�8bTl��j"����^��b����+�]�A%�x'�z#��-z�����<ھVq�#�@�װ)L#U��hN��P�����_uf���R%ѵ���D�SpB�{ZoEΜ�����k��!�2�Fx#.�P7L�R�~s-c���뻰r.U^vƟ�|�R�����+W��&��7dw��?�>��q	P͍Ttn�"��2��t�Źg��C2ͯ�A|�P��(\*�"���~�y S��g�A?�0[`��:�xk/����(�<��16�I��e�~��es�Y�i
=F�L���?������jX�(�BJ ���c9浪n�Qg�`�S��4uMvuu68��~���-?���湵[��lbG�i�'!���=��
�^E��\o�P�$f�h��q��BwD+ �~ؽ��2[x�u�X)D<i8��u�0+�N��0������f	�	?1����D��vƽ_��]`%:�ȤC��Q9�*ו�;h��x���r����������
 �eH*r��ym
�4��&k(U��s[�ŷ��_�4P;�^/ܧI�O��4;���ĵ|0kSz�|J��q��S��;�;��ɪ���R��?�X���=#&�٧��i�kf@�n��Ņ��/�3K6���"�^g�������$��v}E����ť��T%a�Ri1oj8����j ����{�r4�ͧ�+`���b��TVȱ�9��b�>TPր[��Uw��j�g�6�v�t���u N��l��@ݝg�|,"��*ɺB�BN��G�w�NnSQB/�B��`0�8�hp:�0���Q��+��c!Op�����p�O��Q�?V��廚L �{���2&]�Y�nu1<9'�E�ۈf��\�-O6ǲ+�z��A8RZ>���qJ��mayplIb�"5���HAQ�Q�����/�0$�>�|/q��B�1��M���3oE�H}��W4��'����^R؝|���2�M
��)9��AH}�dƿ*�^]ܿ �5�����Y6�����s�DT���\E�	��b%�X��H}ɲ�тʳj�l~��!�̋:*/q������\:u��Z-ݱ ��Ҟ�6B��L/�k�!z�]���sJ�)�",	Z���F5��,�����e���͢f����M��x\������w��c���:��6&M���z����pv/8×���;CC�����nn@�2�����φ|�A���Rը��d�7)bp��z!�N�
쟯Ivr��b������)Ikp�r�sa%��d� ]���LNsmV�u^�xѦu	Vw5[F�ʾ���!���^��쭚v<�:86jR�V�(�χ"͠c����c/�ps�xH��J	���6��vШ��&��X�Hs����Q��O�A��T\{/n��xn6�5�i*�r��������*�]lN��_�k;�ي���H�v� �M"1w|�<f�q�P�IxS�-L�)X��
�6�>'-C����4Q����h#gAQ� ]��*�(�l�߲��h�D|$7켟�}�bY8C �3��,��`m�g".Iz��X�� �n�n�.�0v�>�#�����;���/�(d��s�b�x5��q�mď¿��\����݅Q�dy:� ����t�D2HҘ&ȅ��!y�0Ӣ�Ҩ+F��0b�{���D�Ʀ����q<V%��{��C����X����?�5���l�դ�ïb�o����|��QJ��:]՞�����$9��>	�������S4L����~9����
䖛������tlt�r��l�*�;�5b'�ֱ������\�Ȁ�##� B5���;���|E�^���������+�J�|7�V�/���՛��Pngp�<�˽�p3Ll��J�0�b�����p��D_s�?¤��֊XK?KZp�,ck���� ��_%6.[ΙF����8'�&_$��.w��l��hhDF;!Ky�Q���$�q�"�W:�<|ٱJo��uK�+�KËXX؍0=�2ȉd��ʁ�e�F m�Ԛ���/hg��;y�7�Ý"G;D��-�)#��Q��mI� �=>���>�T7��G	]�#O!�r�S50�~iʹ�
(�ýHYEmh��=��~�"G@I"��Xt�"���|M
Æt�}����B)A�tE�
Բ�2Ҧ��%$,�U*���zwJ��KtP��>�⏽��sx[1��@0�۾��V���3���}	��K\<����l�L�I���-���Yŋ��/f��^��8�C��R����z�"p�a�7'�nrH��k�m���	ɳ�5�m�.����$c�c��X�	j�R4��=j $�h��*�����Ƅ�?~���ϚSw܀Oσ�����6R��x�K��w�EQU��"'�9~�n��l���;�a՗��xf�u�cU��|[�~�v&��Z��`�\AċZ��rvR���L맼�)�n�_��>�Ys�h08�j����1��l����dUF����
;;� HUzo��>�$|��A�eѴVکȉ��4�2�269WJ��x���	��[�UC���h�@��B�j�N"��J�8�c�/qY��9�x*�d�`B�G�����T�R��V.�[qa��q}7�s#1
n=�"�Dd��WF��3.���0@���	4��پi0�xl��,���p�GP<��í�����s_,�ׄO��$9"��U���.R⭜!���<���/��&��Z�Ƀ����4��a֥l�wA�bP�������f��(Vw��k�r�=Ƙ��K$�\P"����HE-�����z���a�Q'�F���n��p*2�z]�Px��ܟ�F
}\� �(^���"~>��| x��s_օ�j�7��{ܘ�N4Y\�9\V�W��r�˔y�#�E�+������-O�P�	���?
���"��� V����U��i�E� �~��GE�uء��Kě��j7@v�-,��;j!�e�D��O���r�l6�j��R���ę�7���:ↄ����"x5:�z�,�-U�p�����Vl	3ΰ�O#1S9r�ZN�s��L����?f������}�gD�<AB���ZJ�}�O���*��k��纍�x�j2PR �RV�w�G�%4��ۚ.P������Jk����W�L�&��!d�C輣+>�3qd��ȱe�n2��{t�lg���C- ��7Pȍ�(w�.*[|����y;�l�q�<��a�`OEi�"�f/�=���< <�����I#��e�r�����ԏr
��L�U?$v��]Rj��(��p �R��R����fQY�4`J?��/Ԥvгy8��)��:��s�����6l��2�d	 !�>�=K?��y1"�L���m$����),�l��B�؝ ������pڭU�Pd)��8+�z�+�cNG��
�4�3��N���3��\�D68@Ƹ����J����^lq�̣(�ww�v��={��\���ص����w����e#u��<��/�R&�h��D-�[�ޫ���F�ę�Qw�;�я����|KmzT��T���e�̀��'�q���/�Z�`�e��=�q��Ԁ�z�f;f�L����3f�C�I*�^B|ܜ'�����vx�!�n�(�`[=T@��R�jZ|�:H��wX{��a�^�w���`���bM���:� "���n/>O���۝��N��g��P6}nPt����{N䈈�U�n�"�;,=)�*|��B��<�(FSw �SL����-�`�V8��b:=�,�˟��f����Q�k=3�rD�p�~��W�?�q>���L[���i]+&X�YD��u���B��AM"\��O��n+�?z�8��Y��5�	ž a�;0p���=�1H� ͻlIF!��
�$t%|�M�ӲQ1;]M� ��N!�������(C4�!'�5���R38�7�轊[�4�F��]�9
8�HB|ƺ0�^��� ~�ܓ)B�x�|�]�����[T3��W+	:�b%�T��c���s��ʎ�"�9�J�H��'S*�)��h��*-��<~�u�N�hI� 1Z��46g���A{k�j���뼖�o?�d�,��Ӯ�x��@�(�y�3�����+�K�A���/Ц��U����
���䘟Y��L95M�k�����Q
|v* �_�Й�FC����@E*n�W�"e�c'�wr��O��c7!d�,-b�l\z�c$�E�*��Q���x�O�u���p�WrdW�%�Lf�;'�z{�Nn�&�ܽ3�3%%�Ԟw��pF��f���ܝ{4^�=�fƭU�}<��!:���R����c�·�xc�Sr��͡p.1eH��EJ�pu������ ��j&�k���<���|C�l �O(Q��~�\�	��&�g6���i��:�O^�1`���*�*l���_�>N;�5�5�H��@ .�"�f���q/À�oZ�2�rs�X��QF�'�3��s�I4��	��VucٙA��]Q��C�(�Z��]JD�*7������b�ح ښ���O�����BxWI��=X%#��i3EnI�%01�^�>��/�D����j��dPIZ��
�5[�NĈ��:&�7�#��x���F�:;"{�;i�_����uY)!C�K0n���U�F(i��9{3��׿�B���|�O�<�	[���5�w�m|��Ě"в��*&:�p�Sê���c�Х�٨�D�S�]]������8��;�9DX��S0�;�Wm�~!��=�K�0����P�V�x+t*�r���?��p��qB��Ƴu�`5������-��kX5��:�v	��AU^����^��v�+5B{����V�3�3UE�JU*nb������L�ӗJ
�b�JԤ�Uחz�s�q��.w����Xff�Z��~>�/���x��6)�S��	�H��B�*_��s.R��l1�y��F6��y�K2���r$�n�"
��:�R�|]
o�+K=�����X�V0#%f2Cu��&����l����h"_!�VL"7O�b�L�D7������ Q=hm���X���3r���Try�G���#J�rU�0��f�]
����RY�D�hR�K�83Q~��@j�s�:�ޯ�'E��t����D�)��\E>�����!9�� �,�B�Ŧ����rJ��/)�ന��
k��N��1>��@��p���V	Kr�W5��^���TX�j�G�Zo�L^����q��� �JM��9��C>FQ���_��G"˅���&���>�z��m�R�	��Lv �h�. ���ߡ�c��i��❎-=?�x��$7����I�q����^��@e�Y��.+�ܻ<q��m�� ��/�j��f�]���E,����\����fn��?��ٔ�;�8��^{�f�����HA~�����7�:*\\�VZ���rQ�9��WMn�i/�`���ishK�jr:������e'YF���e:����7�o6��>˦�|�+� ��VՊ��g��u�G4�(2��J|o'��
��kE[��7Ch�U�@8h�B�-�)����M����l�Ͷ�7�x�Ղ�{��G.����T���sf.ᝮa�bW}��:�g|
��"��-dMgW��3)���@�+-�x�Fʹ ikZ�x���'p���΂P�SV�����w��,@=���>���99}�GUA�8�23:�(E
��C�<�l�/2r�{�Z���B���)$��!U��G�AYn�PHB���6�f
n�(�՛Ff��,&�s����t\��L��e��-�q��߰��pxr�,���������?	2�(��d�.�=���h}�YO߈(�щ���M>Q�? 3�szrd����f��ӂ4�6�4����-*���x���6W�whx�&#��됸����
�
�����;�H�i{�U���LE ���~����$9�\d�K�����7�va={�)�l�9�`���Y�rݮ��lQ">j���tI�Թ�T���˴��43��|#xPm�z��-0/b�R8��rKkVge^��ke����#Lq��yNd��������Bf�6��8v�DFZBx�,Z%�����*�ŧ]k��	��>'x�ǘPm�R�M��ǡ`P��;e�.K��U���1T��s�W��&o�d�$�>�>л�q�>؍�9��{�ࣜ2�yktHVTg>(�C(S0���P���(�U*��1ݝ.=yv%ڈ�7*	���h`
���=�J/Ô��.<[��gOQ��I~�fed�<��[��O~�
�L�_?�&��jS�(u`; ���Y���` �Q�OV`�J�*S8v+}8T���v�5rT֜��ѠIl���_S4!Eȓ=�̔}g�����e�6$�&�H �g�B-� oޫ��b�(p�+~)�ff8�F�&˪N��>�i��O���\����H��N�D���Ƴ�y�U����yy�GT��6����I�؝V�|!T6�p���0�β �e�ߐ���h	�**�&!�����r[�����!��[�ԄyS�G<��1��a��|f�z��c��ԏ�s�qfƣ�W��Y��z5��u>���1=��=����H�f6 ��h[�a)B3�^\��Q�^���b�
�ZH�vs�;������T[_jR_�?j�y�uE���{��*ʹh��>�`�i�b�M>�ݱ[*v��~ >J���6 4�˲-&�g��6X�t��̫�N�V���;`���^,Xy*�OwB����cd�w���SGT"���Q`�P8�\:�Mn���奘��Gf�Ů�'�p=Ͳ��}�?L[���L�,��\&S�XY��Ju�ϔ]��$6\Y�qOl�+��z?P�8��t֠�P5řo�a�9p�LOlwNH����0N�d�� ]$<Ɇ|eJ���B]1���My{&�i���>���^4WQ�'%�U�L�R������GL��N���9E�2H�lƵVx^�� 9�Dſ�󐯾8����j�T�!�Rm	���%Sp9�~�L��f�i�t]O���C����*�di�#��E�O·��u��k��� ̒���6����r�k	�>�Sx���ԟ�,?7O��ʯ�/~�4F;�����t5�c�jrd׮�ǳ��D?��]�Θ����[�M�ݰ�����^v%�yFl�T�nC������n���]��"7�r%�������d�A�bf%�z�+J��R	����>ڪ����np7��r�Z%����v����Ni���7&���'���w+��Fa构#^�8|�^�ԑ��?��)<�M:.I�R��.�����X��c�2o��:p�H�qJ�To���.����FA�&����%5���S�̚O���ԝ@\�޴���6��mi���
�Y"�~�w�*e�Jlĩ_9��;�u݊�.qH;�  I�p"'����/MqjQ���#Ԗ�ݒX:Ch�l�E'#D��N�@4Ǧ�Rٳ^��A��]H��^R���I8�dD�Pz7"x����b�� �f5�ݒ�V�(��I��%X�{��d��n��0�E#�Ya���y������d�y�V6!t5k�ģ��µV����(v��H�:�cK���A�z�Ҏ��PР!~��0	�֮�"7F��U�1�{No��:|J�\�C�<�m�͋��lo(�G���,��6T��c�e�;�d�å�%&l�`�z�����x]�nk�c�Z���4E�jEh�g��SKt�� y~�C��xmT5v���$ɫ��A�ntE-'r������̫T<���w�x%��;^��`���5�`'ѱ�
�\C^��8�X͆�1$�+P��r@aV�Wn�n�����[n]Q��F�c�L�/J���b����1�Gs�-�Z��L
�X��-Zf	]?өWE2��_6$���O<�[6]��_s�.-�YllpĞ�GF1w�yAf ��Q$$��"���:�"�|O(o&;�Kö�.tXΙ�0>-12����k����`�|;d�Vu�N�Zh��$�q?�7�P4�r�Dry��_E�^Q�m����sڞ���ѿ�T�eJG?$l#E��r���0X�('s
�Q��]Y�;�h���3�~U��@�;���O�q>ފ�����t(�����w)�EE�J���kҜ�k�ۈ,PH`['���	JgC,�[>��2D�8D�)R�1y��@f���

Vd�������n�Am@�E3��� L�>m��Ɏ^=;�լe�z��Z�������x��Ĭ�"&N7�������<���Sm�Н	?O���c_9.{��� c���	���f�̳��$҂ɦЈs�̫���H��a���J��	�-���gϹ.�����x¸%B����=�m�sE3���9�o�Un{��5=Ȕ�];0��U�f�����~��T�~̖=�Cy����k\wh�Z�"�r,ܾ�t���j�d��һ[��~�hf�oj������d�� 
5F��_�����i3R�uo�r!>��4|�XԛL�VЋL����0
4Yr2,&GJWEf����3$�[�ͬ���+h�'@S�BBul�^�������gg.��5x�e��G��v�%5T=�c��.��GaI}�����/
d�"��Jd��W|��3$~�q�&@;��HDpy�͏�i��x:
�"h֎&��P�6���y�e�c�	,{Ʉ�$��9���U�O��MX������<@�/�L��	6ZXD��z��D4��hx�"�ZA�L�P�����wfe�(�^��8A��h��NQ���\����
oo8-n�=���Һ�!�������&F��.$2G���Ƌ��I^#�<�}�C����(��ئ�vy>��� �'�s�.��`$�A�����4��>�/F�����`��a�;��RB!�a8�߆M��!�
>Z�ȘM~�VZ���PGU`v�e� M>~�����<�*JK�ud�`X�v<m�d���&d�[�b��z��i�ll�Vj�����O������|I�<^�rX�xk��z�y-��ɍyQ��eVb��Qg��I��#g��h��N?�A���z}f�}��c8K��g�D1o�B� �Z yM��Dv�`�k�Շ�C�gxTD�P�(�RL����6��� ���.F�ư�4��9A��r=Wx��&J)&d(�t��O>�c�q������e�[�v2cV�t��og٧>C#�
�R�HP>��(�*�*,��x��y�������2h8��`�v��XX/����\a�<�8$����I�ge�A��^�ʌ�
��LI%�?Zח��ji��(0� �^(�孵;�?Q��+`�v��%�v��@8M̫��*���w��P1l3���Z��!�q1=��V̯��B�;�@��$�Z���b�B�a� *>y�]�ڣ����)�+8a�M�!ˍN���aT,�j���9 ��}���Dl��Ʈ`��n�k�v���-��$l��+���s�����\
�+�߰K��{?e�j�#�J��%�)&|I��$�[�đ����ő��vS����
s�E����^|��zJ1��>��������_��NT��/ð5ײ��H�[��=�i0�X�4�:7�f1ʂ�j�V]3�"ݏ?�x^��p�������vn�ҩ$#��֪Tv�Rڈ�j�����b�����{~��sx�G�`�[bC+5�����R��3��>E �֑�瘆�QA�Vg!63�&t30��F��N�DT�鱝�-�,s�*r�7B\�j���5wV��SB��S�<`a4^82_:3�큛��.]�4�a%t�(+3p�;���.?�d�v�Lр:����&N4�Y��Xub�hx�fy���\�?�O;�+��z��j8��I��+���t�?a*�6p=���qÆ��kHr e��7�O���:$w>�| g����1�TxM4z܄�ڹAh�Ҫ4��~'�.���R�̤����$�*o#�o]f9�.)HN4ư�>^n�L ��W�_�%�n\ξ�~�$�Ti�M�	�*�%�?��6�i���D�{��l���۽��*@����s�`I@�2!�urP�ށ} g���>�6u��}�?k$]��$��nǙ��`\,��"��<������"'�����!l���I3�4�Iұ��>��0�;������B��M}o��C�����Zv �>�MW���C�>�6@�n�O2���S��m�X�M���d�v�b���z����5<�����܍�w.�Z�pRȡrZ~T%�R�����а�NdH�撮^��,���Hw�FYF<$g�^W��Ӝ�^	㇑MY��z<��:�^Ru�X�ً���c�1��tj�p�d�H�RJzY����5�'�ި�7�&��Q�Y/ȀK�G�Oп�ܞ\,�\=�6���i;3˅Ž(=%y_*@�{l��l_Է�;}�I��iH��$ d/�"��=����q��;����N2�(h�X��ˇ@u'�t�)�4���{�Y��AbY�]Ǩ�y�Y�P���D-�b7����`�bjy PR�������`Y���ZI+&�X[���_+�n��0����tZ��%��άY�:�d�����G�W5�lTľ��0�2��r�c|����j�:������Е>��	���+g!�o0�o���F�aaI�{i~�׵nަ7N����D<'3��Cw���4�Ĝ�=�t���PM��q��hà�~�5��_�:���It`]fD�N�����/���R/�"W�SfDӯM�2~ʆv�����,��B�<W���5t`��r�=���+���$��Ù��[���٨�
��絺���5�����Q:�M�i^�M&��[*��}�+kD����3Ve�����쀂�nX~�MRԽ�UL���J ��b�F�4ʀ��os�rIµ�\�z�X��Z�S��؆��Y��ua6�Ϊ���U�x+_��.$l�P��9�]F,R�y��N�H�$"�9" ��:��|��o��Kiƚ\�xX��0YU�29���F<Ӂ@�1��S��\��0h�v�یR7E���/D�z���)��Q�mz����؜�����.T�q~Gڷ!#@�Or�/04��
��
���7Y�R&h����.�~��'@zx��������e��ɳt�Zg��^�)RE-E���rT�^l�z2,N}��/@�{R=Jª������ܛ� &���1���@Rþ�=�V�O�d�|��h�缥�� fn����L�����P��>�e��-�/���������#��ӿu."�6��>����SC�pw'mon�	z_P�WA�^��.ָ��U?c�r�����㮭��6�$mnΦ���'��?R����O�	���y�1�1�TjF��
�G�J���0�����K�E�ѿ�G1��
c�np���Z�O�-;0G��TP�f�c��~�M��~�V3��8s͑o�\�j�Zwh�rѢ���v��\�_�F)����h���jh;�]��� �ț�F�K��X�Q*�m}Oo,N6>��|BX�6��Vˬ�O��UT4'�2�L�J2;5�5MV���[�������h<�p@n��B��5�ߤƑ�c��4��b˶JDix[y뱭OG�<\q�TxH��'�.ׁ=a���}M��OK
��>"e�Wdá�W��3ig�̕9@���c����_�jD.i���xՙ���N���XPm9���o�����>��,��� �G�m�934�U��A�h�b��?��y<Y3/h�����Z������_d��+��'tA�J�P~����>f�~9(��S\��	�)Oa��\!9��	��2"-)�_��:�f���O�������<{2�����EN�dOQʷ��}��f��:(/���P>�e �l�s�
Z�ۃ����I�R4*��*���hYO��1���K��kR�-<��m��!*޻z��
����S���qd�_F_U;�¥� �f�~��GV9���K��ۘ�v�	���;�f�V���@�$e�l�WjÂ�J_�JF·����L����-T�x�3zPV-�Z���ڗب<xV]}	s��]#����;N���t��Sn�f��w��~I��ypDL�dBnm�Z�tm� ����D"k�b���x�P�\�Rǜ�>���4U�q��.A���4r�>a2���SW��&%{@dc�ټtQE>�+iqu�c�@�p���2>S�t�f�gtG�CY�����P��k(�#*�� �S^�y�K��Bҿ-�C�r��`�?M�s8�/j�7��<��ڔ�r
/I4d�e������E��
�}�L��0?��!��Oj�0(��� ��O_�R4Q
��`�Q� �v�.�8ʶë��+���RIG�l�a��UG�!�:�=|����u*ʽ����$R�#~.p�]!mB�U� �J�)������)0�8�?��NX��_�K4�Rߴ�u�5���yD��ƩK����&&����7�=�����'��C!�	�@
�>�澢�f�4��MMe��^�E��� �&���uЁ[萷�����+�J�2Hʽ���Ѡ����߉|��z�������ǧ�1��eZ�8&��𘚈�(��ѣ=��ٓ�L��E�f,�A�]���ע\3�Ə� ~^� #�����hvi9�oaő��T��;RU;Aj�����|�H��{y���oꨈ�O`���b�(�rI��њ����*>@c��$ۘAn�\?�g�M;6�tn�V��JaN�R�f�c�S��,�y�*�V�B7���� Uw�$�S=�����`8(8M�i:���\I�����ϣ�\�>��NRp���*�?B� Q_L���:�e&I��YU'u� �O������\ϾO���+	�z�"�8>-��.1����O��aez(p���v@�"��H-P7��^��Y�曔�$�Ӆ|��z���H1L$6M���ܟ��4���t�&4�q{'[���b�RD��h[@�"��ĝJ9��sH��ƫ�^ɱ; ��+�zus��Gپ�M��_�ZT���HI�	K{c%�ʴ�	���z��ӱ���O۸�E*�;��Z��{Y­��uM=N� C��06xk�86Hk?$�I�I#��8m,u�N��Κ�Q�����������M��P8��������������¯��v⚽ �MX!��~o��"h.v�/ub���*C�X���dn�����f��h�ع`a�Ք�.d���b\��z����8ï�`������`��,pm�r��}%k���b�K��N_���V��d����w!��F����p9�nݡ^7W�w ��Rn<#�:$�\RP�2�����Nc|P��h�p_.�H�ScJ�}G��E�b��|N�&����X;� ��O�? �;�\gX���#6�Ii�������XVT��h*żl:�_o��;xUR�F�H�aM �3"�+ըyzq���������L��X��ˢ�l'��q4==���>�T�ZA�.�]�)d�b���`$���Dh��7X�s|A�b�y� ^G�ym�LG���94If��X����Z��nZ�0bS����w���g·�L�md!�^�$��p5��}��h«/+��~���I�*뇬q:LF��l��а��҄�:�`!�[0?I���3F9��l{����0������ ^�<�wY���"��de�&����`��]��۾��A�Û.��
>����U���]A�l������U�*� �V��/�S�4{����~��ڼ���ka5��:[�a���C�t{Îr�����G�!ǡ�B����_��q_.�H���|=��f5���'&����^�P�
�����+����h�RV@����:�I�nS*��+B���~L�G<J{�Nb�g�o�×KKs�����π�	UX��0Z\��ϒJ����I�6��D�yp���'_�.��l�P���+F'My����}S$=&�"{�6:�"D|�Bo\ [K/����XD�	0t�2����!�`�{�v���;�X@�ƅhS2�ۧ��7�]��LD�Y��r�q/QN��m5=������w���TT#�fGuk#;��rf�X0��93
��|w�Y1�(h#��)��~(3@5��Ą!x@I�@XV��t^�F���)��Eo���Q�Ғ �ꑌW,����$��v�J2�`!�����{3��߫�1�JR@������ Vm��:�7�t�����9�L/�����������/��,�¤S�;0���Ӻ^�"�>���>���Q��emJ,�	������Y��.1���c鍿�.B��m�)��$z��f�قHV��{� ˂�3�����l����ණ"���k�������X6�c{E������D�n���P~x�
�;K~��j�f��.�O*����~�6ű�A�L:[\���Z��"r�嶴�M�(��Z��qP��E
vh��qj�� 8q�X�x�6/uF����vPw���uo�I7>\�|}@��G~V����x����� 4B�2"�gJQ��p�i�p[�ņ�H�Dh��^@�rtBko|��eߑ6@à�O]�����\x�u��f
G�cN7��T�/���e.�#�a��H}�T���
Z7"@�Td��jW��3�̂'�L@��j~B��=Y�EVi�xp>���b���P(\����oP��gt,�����$�p9���Ur�,������z+g<�F�/"d���Z?�s���z����ʥ���A
i�P���ܡ f7O(BƯ�n�}�^�'��7	�\��^�m�%�-��%�0�ʺ�Ԭҽʁ2�4\����k2����<i�`��2-}s�� =R(��~��J�>b�� d�as�q�V���v�܄�4ŋ�%���ý^���;�16"�V���߼&U�u!�
�X��#Ϡ����[#U�c��� �Μ~|J���؍�K0�S�V��v�,I��v�֫A�Q���j%�����l��?j����[eą�ط%Vœ�=g��4��o>x��Fz�F�-� ��\r�C�VX9���갿*�#��^"�N�v��8A�f�k����i��Dg!VB���Z��]�;S���Èk�Y�����xʝ$P���RBt�t�ם��=.<��f���'���Wn#& �jd�8R���>��qДٍ�Q4�RQ�/2p[t�Cg|C���ZP�D7(�4Z*}�.&?y'���a(D+��"�`;(ӎ8f/�m$�'�<��8��cFI���e��������	
��*L���?�����1j�T(��s �-��d���QE��`�-L��[v<�8�@�Z<����-�{�}li8Y�P��!V$=7Ҩ��!��8
6���1$���p��X�QB>ji �] �Dkfڙ���{2)ky8�쀶+(N��g׉ރ�̈́�ͤ�PG����!D�֗ƤV�$4l����`
��%�q6�b���J���eg�ء�ɰ�MD�q�Ge���E��̎��&2�@�0��[5+������{]ą���"�� +����o�6Y|�ez@�������@@��BQ;�����<��zF��)P�Q�=j���19�ptDf'�\���,��@3�
�5��^��Ŝ9�+��vdt�����Lz�T��pR�j!Ь&�M���{t*/�ʁ���f�`�Zb9F'M��imD>;�[�G���{ew�gu�!6�=t��x�|%�NЀ����u�?!,�).*h
}B�X��w�j�S8�q�	ϒ`�[v8h0|:)�{�7ΉR!��jTqW�%�ޑpny��#�A?��n,�.LG����?&D2�Y���u�]����'�R\
^O=(�+S�zP�;8��<Ŋ!�@�*|'a�$ps���z�9�}d�H��إ��b�v�$�#|6 ����(1�M���ܺ)(گ��O��42�'�{��R��#���)?�� �0�%�9��H�LLƦ�_^$�� j�c��}��dSо�ȿ���BT����C�	��c%��ش��Ͳ_B���9������۳��*�֎�Ta�����(DPu(�-T:� ������6�����kZς���Ӗ$�4�P/R,sҮπ�ᬣ��e<�������{��w-�V�E�U4V��j����8��M3��|���v`g���Ѕ��C'3s�,��n�)ͬ��!��c���Ӊ�On�dAb�`zhC��1\��P�>��xڻ�g��t�p�h�rP%�%F���'_��$NZz@�H���G�@w��rF����ԩ1�	>�^��B��m�A�<>��:�ՇR+㼔O�҇)�cw�β*��p�Hu�Jp�%�`���h���&����������ؐCOϬe�+\��,��`�6�#i��[�;��sMo��*��luyE_
��;s������Hl� ��"���ՃNYqBz�P����#��ܽXk$�˽�,'�5����4x�n�#!�O��A$�]=ʬ�+�F��UD���7� UwB�b �Y Ɖ�."��M߭��I�(WX�E!�U��n�g�0
I��V?�O!�b;0VS�d�&��bG$�5G�j����&�oڣ��٪����V:����'�#������k%����!/��0�B9��I�F�ڎ���{��3׫����1��;6<]�3��)�}� YG*�A;X�O鲆�M��x��r^Ö�#6-�Б��p� �?�]����|�+d�%�q{����(S�D�C�j~�l��)�&6���pɼX�r�Pt��Nr�<��q6��\�����ݛ�����#��b肇Qn5_��b���o^^���iر�b�f+���㽽V�Z��4�/nNҠ�%����L��J�-8bdFx������'s�\�k C�}�,X�B�Z�H@�l�%���,6WP�`���4����_��F.��lqI�o�F"hiyRuk��B�$X��"��<:_R| JRo��pKz���X�+c0�2/c����^��40�M��	 �_�[hH���7;�i��D#ݖ�0۬���Q���m�m^��4��x�b�*T^�G?5#6D�r��A0��TB�
�8a�WS]Yl��h���$�L~fy@�Qg�ߘ&������1n�t�������)�E*��9P���l��,�7�19:�q�xJx�m��� �C��`/����1*��@71���FVu�@�Ջ�K�v���U��F�	Lʞ{��#io�bl�����f�%���N:2���Y�ӵg"7g���N���h�ft�m%
7	�q���T{�.�?m��܎c1?�z�&�����d_�$������������T�;�҂Eج��:�ܧ9Cϊw��e����V`���N��
�E�o�ὅ|�@F�n����R���S�;f���J�+fdW������:2~�6�T/�%	\��ZmS�r���%ا�밃U����z[� �Th��j^�sQ�������q�F�W��ѥ���E���o"e$>7�|���l�\V�Nu��/��aMq4]�2��	J膃��n[�񝪣0Ah���@�`IB� ���F��q<��jӔX츶 �xќ���?G`�iT�6T�]n.��<aZ��}��z���
�b�"Bd9��WMv�3c����_@lJ���v��� �iWBxi��7l�P��4���-����q,,:�V=��99�AU-Y[䞇��'��Uc�<�y�/���s�Zi�.%y�$��cV����AE��P�����Z�fv�(�� ������f@��J2rR\W�������-�l��K	��\�mҘdm"^�x�����2X"z��HȚ��ʭp�}N��;�=(e,֦�d%>�R Vs�"��Ѣ��Eܿko4`=�� ���B��ߔ չ�� ~��|�8��WCd�p��
OC�ɽ-����U��U����8�* V`~w�����H;;KK�w��ydvͼشzq��L��*ݚ�Vl��j���6�5��Rc������N��M6ߠ��Ox�yz]�-���>���ޭ�VS%�b�z�#�)rك�N�d�s�n䉵~f�ϙtk��$�JD���Bd�Z���v
Q�1bGk��*�TDix�zP�$�R�k�O�%�L�ڰ��.7�����툴!�,0W�X&�~�d�߼��>��q+�o��DZO��2��t4��g��.C��c�CPo�F(�iY*}U �	�yb�؈xG�#��(�`�0/өX�/�,��<G����es �YI�ThePj�#ȑ�;xT
_�L��R?+�}�!0jz`(a� +��E���.Q���`Q�~���v��8@���.;�!���Q���l/?�K��!�-K=��� �ʳY����$�ϑ�Ѡ�S+�B��� [��_"x����e�)�;R82�~���NG��탻o}�H�"�+�X�:�D=�Ɵ����:������3V�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��} ��UWP�Hh1�;�f��l݇�Jߚl�.�u?W�������Jd�WT�VEk_+�o�y�wϢ�w�Yc$�����^�l]b���
_��Dd�3ٱ���k	�9%]���^Al����}���V<�
=��s�'KK9�#�~v����B�I<���[�z��!������c��D�P �=�����:����e��$^�]�]��.�(� ݿ�E�o�hO��z�Sp[�(�혾��K�Ǿ)J;ǜ�zH��z: >ߌd����+|�"�<�H��l�
�M�tc��X,�D��e�b)��n+yL(�f7X2E�3�.�/���1��7��؈MsQ������{�+'|�.��C��@�7_����i�)j��{�!� ۷͖ٳ���U�!�0��\���� rbExy��⵭��T�cUc� �'�a6&~lx/~"\�&���+.G�����k/�~��<�Q�]���/�UZ4Dn��&]�\ֲ	0���+e<�6�p����ꓭh����@��#c	��N�
N�p��Z�(��xmW�wyM��({Cn$�]x�I���b
�^_�Izmh� 5X��.��,���$J�K6��\����ᡊ�J,+%��� ��^�����Brn����WwJaÍ���>\�D����Kq�Ţ���c���"��Y�P(�=�q�#�2n��M�I��6
���d��!N_W�q\[���#AC �+�IR��<R==�b��u@���;�����CE�DЙ@��J�3a�G'�(�PRi�~�Cvw��AÝ��QTa5�~^�,\P@;uM ��W0A��=-���1���f⦴;��ox�"@���jZx���y��Ǽ��o[�9� �%�O3�`������I>Cшmo�Y�5�v[�bA'�����E�u��%^��'��81�V���t�*"o)�}�F��^5�AC�okpȒ��<��	��Y#���I0�Yb��s��`��C7�(��W��2Jq�9� ��Qz�UŅ-�J�c�Wf(V���_��I�K5��U�wo$1v3ûloN��?y_J}d�~�!x��P39��s����l�������%��;��
r'`Ļ9~�_~HQ��9���H�-n���"�ep��+C� 1���7�]I�F�nOe�c�$��j��G�P|��ן��3�2~�i~,54*��F6�`+(���M�"����`�dcSY��������ǭ8���"Ϡ�MP�S
�`>��sg��L|S3E�8�&I*���{ϝ� �Z�,!�`�מ�B�OjzvV��P���`nK�=M�f6Dd��I��y��"�{K�'� ]��{'���s 6�d:�XHa�0g�W��8|�1-`��܉�׽���>��}�]�_���̐f���;Ze"�ց8�%ꃋ���X�]v��"E��/Ew.Q��7�t\��g��kڋO����H��w7�D�LreQ>�7�w<��_����z�� �Ҕs�DH]��Sc>�,�е-Ne�:���ڔϰ[V�'��D�b]���D^?�ă3�{sσ�?���dD���F�o���Q���Zp^w=����"h��B������H%?������]�RD@3�#QŃ���d��L+�Eij�3�� �MR���ݔdǾ�lD����-%�� BC�ߣ�g��0��y�):��3�Q��>~���!�k}�g���y���&�KZ���	O�S~VUT+��_D뒲�L+�75i�`����"S�	�ج�¥���d~��-�Ytn.�`D0��#1��Q5�	���TZ�-��)�/��D����%`��j��Z�-��,~�k,��C�5zڅ���Y;�%�dL�����g��L��?8\��Yn&�Q�����a=&	�᳉�2&�@�'�3��nR�S�P�i���̨�.��i�U��P�I@k1s/���v������'��2���Z*�
����"��5���'Z�4g��?f~=�o��6�\".$����4'Ӯ��|�ww�6�no#�st����~e� ��I�G�
��L|�
!�?cqd����3�Q̂7o��Io���[r)�x��#A�$H�"�eP��#����$�:�B0��k�^��#R|���cu*�M4�v�� y�>��0�-
U;H��!��C�q^�k����K1��η�����¬��Wk�X53���*�-�d�GY�;�V��Q>c���V�z�)2 �h����|{r^r��E5��;,v�yU��'>���wr$��8�����8��k������]>��#�oP��'o�j����s9C ���e8�ݕ������e�&Ȧ�`՘cꬽٓB*m5[�x�7����E¦e��*I"�7ʑ6w�E?��������4��W�����)2L�oMm��?��D�7��UX��m7AcK>ڨL� >���#�����P���M
�2^P��뷰=j�i��Es�$[��6��to��a����T �ǡ�j��4�xF&]Eq� �@�;�)��i ���%���6ɹ�n�hZ�xW;v�N�V,W�35������˧J�(��2Z�������l"ڵ����s��K��#����c�譨8n?4�pS�Bc��a�Y~�8F��%��fto�b��4���1S����?g[-e%\�g�@�R�D�� ?�+?��h�=	\��[�:\���ۭ�� l���5�;v
�hr�����o�Y��I»X��`5О��-q�]0�sl����e7���O'w�:Էh[sT>b��=���N�΀5a����޲���4���/u\�F�� ��C�Ҋ�v_>�0��d�-.[��:D�c����#�vR[�Ҍ��I�O�3flq��÷2^H��x���&�6)�쬺С�;��R�b����L*_�'q6�!0bX*o��1n4��w�x�����*���oL�<� E���Z�a���t�lw"�*|t|z�_1��1Qۏh(肄Cd)�Ip��?�`Z�޺��?��MQ:W1���T#�2�� b�+P�,8/��V���5���Ib��D8룪�4~+�"��r}�~�<y'q�<lF?5�8AT�]k9q�2�^)���r,=s����yʒV��GO�֨�����`�$,��3��� [�2B�C�\�� �ї�	�䊇e1C��p\�8�z2��eّ�u�~�[�]_�tF��ߧ1��f�y���)�
- E�	L��*�F
�+V�6Xwt�w��}��AI6���v����>g���#mm��U�Pl��gS�2��ӑ�����oۗ)Ym�ө2=��??�7>��Gp(t�[���u__��F�ޫD.T���u��tGe�5LB陖�����B!2s���Tb<G��%'�
������7aڌ�!5��f��y��d|r��~�21/�t��-����\�� ���:��o��Qx�����fMJ=����v@�4��Щ�-�@������Ό�b�L�C�F����W����nզ���Q:�0j�AbɅ�����tmA��C�����v,�.��L�Z�@ 3��C�XJ�>x����a��N�9z-�E7m!�w�Z�Cή)�[�{��bc�{d;n�������("HG�}�p�]d�p�c 2��`j�Š|t⍆=lp.~��p��˕��9�3ae�)�L�2���=�9��a~~c�"I��C�访��/����2?�{��u$�^E��h{�nEEi�������9'���$A��h���ݢʕ�Ҕ~�X�zƸ���6���s,>BR�y�՟��q��~�\�cWR��������(�By&3���P�MM�1��:<٥����耼�x��sj����kO�2 c�	$ƥD�j�rw�cxvڰ�d�& כ2Ѝ�٤vDhf�����(���x���D���0���7�YT��2@�Xr1m��o����_s�}�Gs|mY��H��Q+s�:�>�3Oi�4��7j �7&�����A�@�!��8]3p�/�y"��+Df�LVNk>(@�[e�=��A1�W˚cz{�#�T�F���|�j�~b8��h5H~���r�q�ìWK)G���/G��*�V슆#9D~Zx1 �������6��mA��g�p�e�eN/��m��j�4�
��≨��/�8��.�#Nu�3�u�`�L
��ɨg��I?"כA�� xf���[��g���t�iam<�SG�����U�k�JL���2��8�|pY�=��r���B�qg<��`@p��p�B L���ARr�S3�M�Şx�z鬗'?������.# �e�RB�鷏�d�
L�;C�pԀ�h����#G��#�h0�	�y�`	:��=���#QS��>�H���\2giR�y�|��I�K5���D��S�T&.�
j"�Mhg8/7��`�u�!��SZ,Zا����`d9��-�Q�n��M`�5�����KP'Q0.��uC�Ʈ-���?��Z9������*�-����GL5k��T��5���u�u�Y�>~����������BJ���t��م��on��<ϑ����f&��d6�2a�e������~�n�՗S^芀���z?��	U�i%SX��.�@fiL����1"�����[����B�����Z������"���Iؕ	�Z?=�g�f�P�o!�
�1�d"�&����4w��)/�|�:�q�o�Оt�Eq��` x��I���
�5�|�l�!,i��)��*�֬�q7*�I��ێ��K����B�#��9$C�z��^�ޓ��6��̿0���љ�#�ר�]�u�64��R�u�>~u0_��UH�a®TX!�؊���k@y��f��I�����s��h��g>X0��T������b+�;l���j�.��wy��uN)���h� ��9|r��� ���@��v��yU��!>H�7�2@���k��Q������;�eE���N_>D�t#ϪP+�o_a����9~�Y�^(�3�R���j�rp<e������>[�� A*I+�s>
�3(� �6e4�@*ĮV7���6�6�?43[�����A4W�д	�~ ,L�6�m:e�?��)D�TR��c�(;~���#7�L��M��F�޾Eǽ �%�S8����%e^����͢jVTr�^����7I��/�ʸ|���y�� �r���-��?_exA�	E�R���V�j�� �S%Qn���^c�iEZ��;1Za�q���b�����֎���(}��Z;�B���l=��Q����<%�F/է:�����p�ClQ8)��dB�﴿��Y��MF@h�%�Dt� �o�w;����ma�S����2:�[Ȧ�\�܃��*���� Z!Z?!h�gn	��C[����6��5	ls��5a1v��ehM�M����
6�Y����lK��K�5=�>��%dk�^
��;V�V,I'2g���s��}=�	=�,KD<��!\aG����~��xR�֩7�2
�1����_v��4��*����.�L%���:3�á��ļZ�vn)@[@�=��b����|�2�q��r�Ra�H����$`ԛ�ڝQ-�g4q�|8���"b�n=��a*�tZ�h��<�	b��Ao�!Dno)>w�}����*�n�*�=<�ڽ�E
�<y����}w�*i|o߆ɺ�(z?�Q�T;�P��ܣ)�����[����B?�Y�QU�O2#�UB�;�+�5,3(�ޱ������d�9i~�8�q��ol+�l�Z}���<4��®F�~�8ͪ]����ͨ\)�g�͚0sbQL����8�"s�� ߙN`�~���̙���ˤM�
Ch<���1Bxߦ��䅬#1�c_pʫ��SK�z��uߌ�6+!~d�]Z�F��"�죈������ԋ�M
h����-���Fe��+I�X���wC�/����A��%���*3噬^�<�m�®|`#�+�Ţ)2W�ۑ����P~��R�lm��,2���?�C>��0G1!�V�O�Hq_k��3�ī���T�ˢuؙG L�L)%��p�؊c!!�v�'�^T=�a�����z���L�)���I!PS�fW��Vrԝ��z.�o1��������/�ߍy��ф�_'�6�>��M�����yՑʍ�yO�&j-Y��P�X�ɟ�bD�C���4y�ҵ����Ц;Y���V0e�7b$#[ǳ�t��z��D�ڬ�����ɾ���=���@���^gJ�O�tya2�NW��-�����w�
`�u׌�)# [����[�cg�Wd6�\�����(=&�GH��p�1����c�6��jA� �4t�H=�|~Qj�p�+������2a`k�ʧ�_��h=w�]�<Y���D>����N)�o�~/lMK�M!{{oU$�3�E���i��i�㼨[5����lE$j�ɣ
�x�����~�Mt�5g�
��6l���NW�B���p��l��~}xc~���fV�r����ya��˩�NP� }�����wC�cҺ���@�7�Kj���f�2{��e��_��jW��w��5vX]��� ���2+/�q D����Q����7��U@��v�?�?ы�l�,Y)��7e1�3��1�F�
B���W_�nt G._7Y�N��+N%��y�23�8]4�撌���{��� n
�@�q�5v3
c�t���g�D�^��\�N�Q�@�e�����71ݰ����1{t�x�����W��޹K��0�mh0l3�Vi��,�Q�(=VK����h��j;����uN9�L�x����x�q��������p}e�E�Nj(�������\�AJ��֤��e6�)}Nv��3C%r`�|I��B��Iz7��ܝ= s���2����1u�D�؈��� �>:�#���jZr�}�tCuJ~�:���G^ F��O҂���9���g5lz>��f�\x�}fT�OOX[T<���"�\��El)�'��{8\�Usi��|�ìs��	�o��)kF�n�p����8z���-2��|��CG�(�Ҁ��o�
�[�.��#����9Un�<�(Cݼb~;S�u�5�������Rj�]K%ms��������R#���\8=j�e�ϭ�t|��������D���@�H��bx	�8H=�Ñ!PR6���O*iU�lV^��5�����t�+����ծ`c�<�ށHk��.l���+�4��0g�O|�xA�6S�k�9 �����|��7E�����x׵����
Y�Ui�,��(�|�%1#E�̴
��F�G;e�y��s��xhU7���不�;,�f<M����-1$�@Oqy���*$�����.z,�}���S��⌝����V�o�9��v�>H��˫S!J����/u��xB���k�eS��F�������s9��Mp����XN%5���?`J�w�l�O��f{	FE1rb �u�:,>}�`-�r�r˕��u�~����V�m
 -:d�����LfN�M���F�m��
;�����L��N��aL�u"��/�8�M9N&�&q�����&O�2a�� �*�83�<���:;�gf<�;�c3����� ۿC��1H �9��Fw;�����h�����L8�u}b�V�Hff`m2�e�ۼ�9�,���F�v�,`���e
T�|}����Wwp��j������V��'�S����{"�:z����u��A����;)�	�&�%��������~���mZ$�V�Ջ�0��`L}5�z'4O~��[�)7�Vw�d;e_�hhr��ۓE��5�Q`C���&q(�S������t}��ʾ$;/��BՎN}B�F���
��`�Ɓ{}�1Bp��OԺtN��W�H�ؖ�F
� Io�na9sU�®ydU����CW���\\7��CID�FC170�����d�	K��Cҧ�(��~��9�s1vv?��_��0%|���}���S�U-��e���M�D���Ԑ�~e]'x�yQ��צ�&�޽�,�=[ C�Rm	Zj�r��S��4力���i·��նxU��*�@�Sr�x�ח�b���#%���%��"Կ��Ĳ}�gZ�P�{P��6ZJo̮�Zq�"�^U�=g��&�n���7���b�q$�k	����Osu�t4!&�+s��8��W�R.����!�ưs��������F���M-W����H@���A�~<qP0Bڙ`^���2M�^�Ք��U��5'|�Ȩ����q��?����&U���o4$�=U�#�'Q�,y�y��d��|k�8����4�i"��g���-�#^����3Fr��zRy�2�ހfܜ�>�Q�Is��v��"�*MH�(�]�3�'��`&�-N}��y���b�+����D~�z!m�ٶ�B��#Xy�uKz/禇z�I�17���C�2B���8��T��N�9W���d?�	X4�Z�ꔯ8=��t�  �ni_3"*/�p�-��A�{3.�i4���x2W��iV��&qi;X�]���C���D�nd�$���[���>'%/�P:����C�@&���	D�T���(��^�2P��u`J��ʼA�*Ъp���hM(�q]�� �FJ�5��.��x�\��rS1���~�[�(��lc%�_����0�U�CIq��� a��L�w���t>��=��)u�T�^L������+������'f`"����3D^h�Cw�p�,y������}Y6E@�ct0s#��4��:�Ѕ� ��`�帒����;J�w�Ӟ���x��씅 ^J4�W�V���_0���E(`\w���$$پ��l":��R��_��dl��T��P�Y9�4`��&ollx��f��h	��\��'���9q�@~�Og����6��2 �P�>���^���W��i)� �|��Jv�����A�(e�y$C���.#�7 �kaE�<��m 5��JzZ}[��0�j{��
��Ⱦ�Pǡ�&H�lz{{�qH�	}+����m��jB�%���$���X�w{JbNG��3�y��f<�+E/�.S0����k�&
���BsJ]�Ja|{��|V*�.?�(�C@��_��}�{�)�
�{�۴ ��H��(%��@UhV�U�L�!�U� g4�y�����q��9�U�L��:&'x��&㣡/�F���s=�ZdG�L��^
L��*C<Q�~][�[/��4�犁k��AM�	�e�8�<kMZ��W���x�k���5����	L�N�#z�5ĄZW��}0���{�ҷ{(j��r�nA+���i�â��Nrdh.�5We����]������^�2}���I��FXGJ^�+
�!�hH����h�O)E��'`��B;J��J��V�rl&\$!��t��͖�C�0=�ּ&�(��������5�1�l�vaΧт�u|�Z���>{�@*Щi8�Is�� ��90K�]��]kF�=�`�T&{6��|�=y�b�	]r��SK�Q�����E���!��<2���@���r
O~�[�@�2_#���H}��D�+��b��v��4�Ps�2��\ZS���+qO�^��=+ߊ&�꼇u�b�?G��5�#kM9[�`78s�It���&2�z1�8�TWd>[�*1�!]��s���k��F�q���Mqދ�}	�H�<�[�,�q����J�{�M����0�a�u'�+�� �ڵ��?t���W����4m4h��UQ�0'��o,=�[y>{��s��&�i�ȭ�4��L�C���iƥ�`	�I��]H�5˼F؎N�<��R=l.�"��`���� sJ����l��Pz����!���kM�`�W5-�{��=��60:�����zeW�z��B�Z#Ļ���_z��O��w��C����aB����n�T�td���h���[���ᏞyJ�s
��A� �;?i���*���q��A���.�o�!��4��W���i��W��C;�Lj���)C�k6DgH�h��ۊ��B��'�J[PIΚ�U��C-������MZ'Tfx�l�m^�u+P7��u$�r�v�AQ۪���,�r�,��$r���|����rwGx��>�\�B�����=�[�Я��%��������I���˔ѐj���Y��|j�m�u��^�9Ϳ~�|�oOAm�c�k�"F���E� ��$E^�7C;��p���S� � }�Y�y�^0C07���x暼��m����$O��֪0ݰb>J(�Щ��b�ы�g�d�J���W]��Vn�A_twT����X��w]�z$h���ґ$lf��3_��d0���?��X9�/��jl�4r�'��>F�݄��[Y�'��9���~_���u��r��0��:�_�ī[�L�,;��-u- (A��� ���yRe�g$���&�^.�: �3�E�}����N��zK��[��i�aUƲ�^��TY{�RX\�刽H�wz�ɂ�5_ԌMl&+e�i�E=y��B��Z�̶>��;fXՍ���n�b�a�w|�yuh�f���E�!�.����_���j�����ssZ"��Bd{(��|L .�FU�s�@��_x�c����)�o�{ُ DX�����?�U�U��h,�e���y�5qyt��>ԛ���U�O!��C'��~&��/�K���!��ʂG~{���*�g�<���]�u/$�T4�䁯u-� R	�&h��bu<�9M����1�L�� S�Ba��w�A	�,�N���y��Z^��A�����*{��˨�-�2���Ɖ���.㒇h���5��g�g#ٽ������R�TV��}>�c��
��J��+Β���cƂG6���%��k�2�`^�2J�8��6�u\h@���!��T����J�]x��s�⌶(���q�ؓ2WJ�V,I.��6S�* ��]�Z_ �q%�a��J�C	��!�K�z�L1D����\��U_/]��X>N���r�K�G���o��](\��%a�f��PX�/�}B����-I$E�u̿���%�0$�A����{������eS��}Ȳ��_�rĝ��c�����\-�������=zQ�!���&��#�!��n�4�2���u}�ܜf������*oq����	T*��J�D������f���K=X$xB�u��"��%��a�	Գ帀8�2��\Ĉh���A�P������;R7�Y�����a��Ȥ��WiR���_�G�^Dgg��Z�����E,C���חt#�h�t �g �\l0�鹙���6yAQ�r\�t�q�����������A�/a۠A��熫��x���N�.Q���E�p�+��М�����(}7h��w�{���O�m�i+,�s�!�6C�(Ò�M+H��s�nƝ�l�,c�d���w����ǹ(L�XGϬ��P)� �lTG��>*�XE83�Ķ�2�e�p�ϩ��u!C�`'{=�N�j-,��D݁�?~nWWM�6P��9�P��W��=��{Ws����5��.Z\6�^GN�+HmDdg|�b�D��1��I��/��C��3{�i�W]�X����r\W��G;"gj��-���o,�]�1$"Ѿ�/Q��.�}N7�_��g���w��Ox$���$��5D�P�e���7���<莉2ȇ������ �DT���ߴ8�8w��2:�+�V��5��V@rV���b�ɼ�P-,�P4���5,�~C������f��{v��ݢt�u4pꇻ=��������hRx������Ɋ�[�銦�R#�3p�ŏ$�����X�ܖ���?k� 01R󩂷`E�d���������͹r/�AI���i�s�g0X��y���:����+K�Q�~>��8�8w�(g:�Hy�儾��Kf�ʕ4sS��T������~�XhL7�GO`#fr��S���8�u��p�d
[|-���n���`!@ �P� ���Q��κ&܄��(-�k�o��ό��5�=1�ӈ4�L����A��8�uk�Z��`55��L6�F�YGBǘ�_%��x����s����鸦KK��&��n2���b�E��(&��#��Kd2��c�3���R6n^,S/䧀u�j��s2�:Wiv�@�\5�@�=E;#��_���e�lu� ���<;�Z6ɗ�g�"�w���l��61ZPsPg�%f
O;o�V{��":�ꇁ�947�:�|��A�ª�o/zEt ����V I��I�|�
nm|*�F!}�}?W���]�+7�B�I{���5���>�X#M2?$��-�qj������w0�.���#^��%8�u6c	4k�����>�0�0���U�H�� !~���}0k}:�W���Z�`��>�N���cv�X���(�L"�S
2;-)��u��s{��h��)>j�hi� ��y�r���Q�쉑�yveuUSݗ>��i�ʧ������U�DL�;�܋��G��.O>�v`#��gP -$op�����9�	1�Ϻ}�q-ݡС�C�Qe�_�!cH�o>��ei�*y�S� A��F;��}�e%�g*��U7�1�6A�?��4�/���@v�Wb�;	.u��ÐL�[m�0s?�D]8��aj�����o��4{vL�Xq�Ӕ�/\�������|�A�^ܲ��4�j��:���d������֋ [��m��׊�� !{��#<��7,xҊ�E}��O��Gg�$�/ ��P%�=b�Bp����Z���;j��b!v���2�)N�'��V*�(��Z�6�zE l.�bU(��'	՗�6��
2�#�k��8�ZP�|�1B�Lv��akY
��F�ĕ%@/��= odJ0�e�~,�S��҃}[9��\GșLH��Ю� K�{?mgh�5+	�Q�[�P#	�ȳ�lD�5P�v���h~�ɍNe�{5�Ya����ޣ��5������5���Mx�ې\*d��'���q�s�~ny8=P��{Z�a�b<�j�>����&�h`1�n�U��>Ս^��vk�%׼���pr�.����:Ќn�M�ML�vM[N���6o����?�q������H?���i��ln}�Bb�x6Эm"�j�hb%�>�7�*k����&�-�"b�4mo���n�Ŏw	�=���*�<v��+6<����V�q�m��� [
w.2�| ՟�k�`K��Q����y�O��)C�j���~��Ƃ;?�8�QF�f�&7#�⢌��+\ק,���b�:��؄�U�z�8�������+�2��Rm}���<7�=�F�W�8M�P]�.b�>4n)~���~��s3�3����E��S_�4ζ�
�f`IyF��A�c�\�>۷Cy)��,"]%p�H����1Oќp�Ϭ�D�z�n�즽;��ϫ~���]��F�y�����������!͙
�EI�#H���TF�+��X���wT�"��WA�']���-l)��J}Ĥ��m��߮�?ؠ\���y2�Ua�4��p�#ͪm��/2�\%?K�>z�G|���篚��#_< �$.���T��	u)LGq��L�*왢�7�[�!߹�8�Tn\��;G��U��Y� ��}�f�!A�Ffh����rU���>�U� 5�9LJ�r0�� e�ߞ�Z����Y,���؀���MV��Z�Ղ�O�^Rܭ�-`�������Z�b�vNC��%�%z��鱗���mi&�]��0��	b��mǄ�%tyj���v��e�(�:�f���1f�7@�6��O.J#U/��pEa`��N�T.-8�ny/w~{ˉfbf�:+[�R�a�c�~�dǶ��
�r=C(.qGY,	p��N�c)���XuA��F6tn�t=x��~bU+p�x��<��+��a�v��X{�TC�=%��r�x�/�-������P�����GG���]����<�ep]���/�,a4n"���)�=�	��=��<�@��U��Э�ZG�#��x�+	���N�M���.eZ�ހ�b�r�A֖���{�����,��s���'�H��k�3/h�rP5|�$�h�8��F%��{��r�w&������f�J�f�+ϓ��̈́���{���1��Eɗ�)�Ͻ�J�7%�\��y�.��A��Lշ���ݜ���Ó�(��%q��2��ä��mI�o6���4�>�_f�qF�#���Cj,J��Klw�L��D��s�]Pv���RL3m��w� �?��m(N�/���X��6��VKש5��A㝙�\3��%ڴf�aXG��}5��@OI�ӧ��rx�� �%ͧ��t�k�m���5f�,��0m���>���p2�c�TL-ۘ��Y+���Q����)�ٖ�X�TP}�R�%o��7z}���f�mg�k�]��N:��|��)�*w1ϳ����p�f���K�̞x�>�*�����a���8��8R�z�A���T���~΃�I������R��
�:���̥�1�g����R��_%�^7
8g^w���8
j�I,&F�A��t��n�g_Hgs�l�p���H����A$7��x	t�d���9�4忤?��b
/�_Aspn���4~������4���΃Is� ���r�5�4`g(�)���c
� �P 	m�P�,4=���	6v�:(V˺M��Ce!�~�(cR�0���z��F��LD4�K�2��]Pܮ�)�r�A�+�93���Ń��cYf���\ԙ��!0SZ`���!gBj9���&��~S�n��%M^�X6c�M����X��p�w{�72��	��c��<{6�4�,�H@�8g�'̐�C'1��KG�n ��l�����]�"ʞ������$�"m⼁w�ꢹ���JE]U"FV/�,�.Н 7~��Bꊷ�O�����כ6�JDE�e�&|7�w,<�ӳ�#r��������S�D��e��Z֋�+�l!�>u���y��/�Vs���9�]bܲ��4��&���]���mb�}Rvϙv��p[������7p�|=�6I������x����$���IA��0�=��R6�3�o��b�؊����ji�Ĝ��[v �*JR���Ӹd��/���4�ͬg��_�L�V��񆎝0�3�yl�A:ޝ����CQ�E�>�E��^��g���ysM���K�[�ʈ�S��Tj���c��:/+��7���`���eE{Si������MXd}��-eP�n��`�n~�C�D��Qt��9��S z-�������b��(?��J���p��k�,G!�Sk눐��w5��y9��]VkYZH��(��O֢أ���˳�S0�ٛ�nE=���B��^&��( 2��v��� �@h@nq�xS�2��H���*��ͨ�ii�����@�V�NRH�upȕj��֟�Iȳ��/�Z������"�	F4��͙.Z�0�gJgf�$Io��C�u��"M�)��PW4��m&p|cK��öo���t�>	��?� �UIw%�
C1Y|�Ъ!pE��l�7(e�pU�7n`�IN劎��ȕ��1#�#���$� �ք���"���������0U�����#�3��b�uI��4�Ar�ߣ�>�|�0#��U�m��rE�!1�䊐�Sk����*�b��ϡe�A�׶��Xt�&�V,�,v��&bd;`{f����;r�ܹ,)Quh�r����r�X�� �����vq7U�>�G�vyG�cb��h��ת1.�܋)FN�=h>�7#%-P��o�|�L7Q9�}��"��w�)ݴ�%���Oe��#�T���c�X �*�Q���_���|�Dv�e���*��7i9�6�:=?������S�W�V��W5��'VLRF�m~m"?e��D~�tf��l	�B]V�gb*L|&��S�ނڏ�D� ���-��b2^w�V� j�d��"��c?¦��5�s_�@t�׽�� ��B���x��~E�0 ����W� R?�%�����F-Z�B�;u�<�5���ޟ��x�����4�(�&�Z�uI��plI���qd�ՊO&�������ֳ8mk��O�B"F���DY��F5%�M���o�{��O
Ʊ�LSF��vb[��<\�%�_\�CE c?Hl;h�	��j[U����_��*l�ZQ5��Rv�0�h���A@���nfY����ã�H5�7��L�H�K��=��ϐ���*q'vʎԖ?.s�l�=e,}�{la �8x��zU�L1����an���`��T�v~���/��C��.ī���J�:�s��eA� �kv2�[�v݈kmR�B�����q��.`H�M^�2���Y*��Kޫ���@�j�]�bx����e*~�&3u� GbL!o_�n�u�w\R*���|*��G�n�9<�q3ۉy� �ܥ�Mw���|�P�~����Q�o-���⷇)6wW^�������v?�/ZQ�˖F�8#u��8�+�n�,w��uG7�4��( ����8�U�ٳc�+HQk�P��}��N<x���i�F���8�4/]�-ʑ�)1R��Dks�3����QnJ��^^�'��];x`�������֫+�MgC����o_uP�)�jk���5�1b�p���~>z��9��z��~(��]�&MF� ȧ0�Թ^O��8�ԋ��-
�P\�h���]vVF)�P+U;`XV�-w�+]����A�u���S���]Ꞥ�
�mЀ	���A��f���12,��|"�@Hۖ�Xm�	�2���?޽�>NXG�58ȚLG�W\_����q��>�TOS�u�G���LP�w��:7��e�!�E��k_�T��.��i���o���vbٯ�!"f��w�c6rH\o��1���Z�L��������$I�ɩL�����]�	Mi����U���((o�X-S�h�:L�QIb�IC����lS�i��E���`ϸ���0�t�b耧����tL�UA^{��L��X=o��_��F��y�b@� ,�"g�JV�[�8*�aS�yN�y-�v'�z�w�(��9�4�m��[�V'�T��c+�]dzn�0��?(��G���pP]*Ad~c|cv�0;��Wgt�(�=Kk�~�1p^�j�/��~PYa�4��k����9�=��n��Dܚ%4l�Ș'��3�j1��	��w{Db�PR+rM�������9�v���U6?�><L���0����+����T�^�7�Y��m�j>8��#C�P�o���|�9�|��R���9���b��+e��a��d��2l���O�*�f��8���t�Me(�0*8�E7�r�6&�D?(��w�`�W������*L��om��m?�	YD@�r���М�~r�*ڗ��L����8�޲G�tJ��G�,� �^?��놮+j�S�R�����ަ+�ዣf
�pa��c? ��FaK�3�x��;E�Ar/N0�J:�� �hG%��,�Ŵ���!�Z׃�;�[m�eGD�"�ş��=�J*o�ٙ*(�1�Z/�w�*ml1����`���Tպ���.M��PH�7w8�2���BR�W��:vY-�5F4ڹ%#�jÿ�o��-���+�Sv��ҦqG[��\*���]q�sl� N!	?x�h�4�	)�[��<�3Oͭ\=l�^5v�vhA
d�q�����YYD�
G�E�5���|�[xZ��}��_��?�Q�J��'��D��ܚsJl1��=74J82�=�:a;�[� J��Gd�|��+����m��%F��A�v���_ ��s��.�N»�S�:�Õ'��0wjvb��[��w���5�r�^�7q?t��FsvH"9=ǃ���p�Ea�۞��p�K��|�b�4���T*���Vڗ�0��bG�o���n�4(w����E�*�|`��th<�.=۹�X�0�J�#=�w�X�|�˼ɮn� Q�\�W-��)f0r�c~�Ϩ��	�?(g1QIÉ�v��#��Ѣ���+ߣ�,�|'ޥ�B�d���Xm���t8������+x�����}�X`<�K����F.!8��]ݥ���')aS����s����Bʁ�����W��ߍ  `,o(���a����A*�C�F	�H��ߚ`|��� 1��p>�y�G��z!Q��i�֑�֬~X�]��=F�Qҧ`�$�����h{���M
ܿd���Ҕ�q7FYQ+��lX�9�w�>���;�A�V�+DO���{Ť���m ��:E��q2K�&��s�D��Ɔmm��I2,}?��><M�G�m����<H__߬@'o�n( T\�uLIoG��L�����[����q!s}�24T1���^ ��2$�<Z ��	'C!D�f��;�zrx�@���4���̮|)���t�#���X{y~��|�T�*q���M�� )ӇՅ^X#�l��)-��R�Dt�=�kb8z�C'3�(ZF��u�����v���*0��b���'2�t|��q! ��u�݈�1�����v�Y��P@/��R�	J��H�h��a�MpNK$@-�����w!��i;
ΝJ[��Pڄ��c[!d���V[�u�(1>SG��0p�"qCmc�(A�;�^�)�t s={H�~Ŵ^p��`�_�q�Ena�Ϭʛ���`�=�Z�4�M��Us2X�W�`�cI�/����AU�{���$�4E5#�� ;�|�i�>ɨ��f�����+�$��^�lG��i	~�\�ߩT���` 6��$�B��B���dc>��,~@�c��$���~��`����y��˝�EPZ�� �R�iH'��{���T���f����9j��3�ڂ)2o08�8�SM�j�T�w�v�{-�� F�2�/]Dw6����e��8��Q����焳������YY�_��`�'p�1�"�;C�'� �b�G��(Y�d����+Bƒ��ba3��c4��憇8�f�A���B��@�ƕ��V3�kb��H��[�wD2�����NZ�@��ehC5��֣1Q����U�{�hn�f�5�>�K���-���$��h�t�J�s���۬�K�p�\"b�ʮ繝����9��x`�����F��B)��}��I����eV�QN^�^�
�;�yh��Ԋ����J����Kݜ�!�Nj̞3��p`��M�z�6�I�b���7� �4�&���j��u�> �L{��[K͔8�:�q\�7w`f�E�n�u>��:��GsSDFB�DOƄ��rzf�?ag���2�z��oO\l�}��OC}T�3����P��)����	�\���ud�p�����~�6_)_�qnG3�����z�5!2�$������w����x�fS�L���Ih���U�3Ub�x&ݰ>�A��;51!���m����j�0�K��C����Za8�
�
���ַ�'�8��j����!�H|�,>$��%��F@Ϸ<���$3	
�]H�{��vR�wA��i��VRB�5aM���+�̑����I��c����R��k�9l���λ��-0��O�K�x5���S�k�C��3��f�|+��E֧���wx�f��=�
Mk�iT����0���XE�d�
_|h��>Y<�_$��l'7
r���@����,��M#�|�SC$m%�qm�0������[�4-�,�J�э�������%����w����y*�>��c˟ԤJ�<��#3Ԁě���?kH�1���+�JY�ܨ؁[!�����X���%)t0�ʹ�k�$��T��Zd8�L=rV
�ъ)�: �
�f�Cr?d���~8�Jb�~0:X�\�b��L��� ��:?1�o�a�h��s�b�@����na@�"/�ޔ,��9��L&e(�p	��]^Op2a�諦�[!3�����;�-�<WD|�WF0�Xn1 �_%.GH��_Rn;vd�@!ߍ�o�L�:-q��Vv�	HZ�qm�Ϛ���91���e'��tT������pRh��t��9�p�|���A+�r���SD5�	,��Ȟ/���A��\�r}e��Q늙�]��8G�f�&��%�mά�V�l)��d_�Tpw��]�n���^4��Y����iVk��;�Hh\J�Ojn�{�QԆU�w�1(oDe���Ӵ��}�k���E1��o���+B��j�G6
wG��:��}�q�B��O��+N8�W}bC�
�
g�oc��-g��6!
dIn$�X��W��8\��C�7d�蒿D1+ز�s:d 		{^!�7T՜��r�?�TA1ja�v��{~����l&p'�Tr��31��P�Y����s�[��^��͐�{]���f��j%&+!���j=�Ϻ���	�Ʈr��]S���~*�^�d��Ƕ�8��|�@yqtr�.�l���#�d���x��9����6�&B[�{P#-g���"Z�M�̢|�q�m�^IT�=۱{&~ȇ%�ҙ�[Z��6�k�9+�Nsi6�tz`�&��* �8�K.W�m����!z�s�2v��4��2��5fM!Sw�-j��إ���T�q�Īڍ�ٻ+RM��IC��Ґ !'p(�W��eu�?$	����k�f4�Us/'EJI,��jy���#f��P��x��4�N���������SȎ��������F�Y���XR����&O�^<�E��s��^��� ��ˊ�e���x�
*`��c-B$����������� �	D���z{7�*��B�	#�25�iz��߇n�����
��2�{B� 	���%T�i��q���ͤ�}�F�NFN�#m��7� �
�iS�w*�Jp�!�AX7@.�H�4,���WfI�iJ�î��9;L�>�9�C��D���%�:����'��)P��<���C�ҧȈ����"�TWl`�^���P�G�uԡ��!A/��d5s��>���U�m �3��x��"�+xd����(�78��R[`{%��%j�ǃ���YmIe�ވt�+�@/y�=t�	s��,1�}�u6��^@�ο.g�������o�"�&w��+2���^\p�C��2p�T��M����Y��n�-n0�+,�(�w�����Į�Թ���k��`9�J؋ũG��xj^�\4�Y�J��%W�Vj�_$�����%�w�$�EÂ\xlZ��Ҥ_��jd�U��H8h���9��]�G�$l`�q����45D��'g��9e$)~F[�͊"���+t���M�X�����O� �q���	������++e��V$����֒2.�J� �bE]��a��V�z�\�[MY��۲R�S�ꌾ��ǕvH1?zs2M������-+�[��}������
C��f��T�X���ks�b�=+�'m�y%o�f0z�E��].GO�������q��s
�$��2{�6h|�nw.3����@z|�_(��o_)C�H{�� �*j�ϯu�/~�U\j������j�ɢ�["zy$B4�í��U1mL'lU�&W�R/w胰?T	�NS_G.B�R�K�%2<E�L]��/��4]���_����N	�KKʬ�<_J��I��႒���X��IE�'��	@�ND���)u�Z����q����»{�x,�������-�v���7���B�h��{5K$�����Q��k���w��j��o��<�JR�(+~�P�\H������C�������WJ��d��q�\����L���{ᆗ�����W��(Vl�qVq2%��=mI�:6�z�1H��$_�0�qսж���C����GmK{G�LǓ��Ƀ��Z~�/�}X�����K4ā�����6��\pa�%��^f~�=Xdp"}��h�>JI���%�ړ��?%�5h��Gg��l�O�Y��Bj���U}D���MM#cl�4_2-�����l��`LQ6���f���s�����M�7���,��ȏ}���f�ǪǨ�ڃ�9\��	5*4L��ᤴm}If=��K�F1x�J ��}���Xeap���U^8Oe!�5�8���i�� ���3o~宲DR�.��7�<i��n��g|�R\f�_BX�^�4Cg���
���Ƥ��5,�˾A�tӟ��$��g�R�l�	j�Ilq���A-�*t��W���E���Δ��/:�AP�ʆ[�!(,���z�]��v�� ���=ߟ�O�a��k(-�ɴj�g8;�M��m]�,q2��ѦI6�݆(s�M��H���*���lc��������6���iY��[i�\�jPيς]��]p�:B3�O���e�� ��Y�oԖ�c!���`�IO���j�g�ܜդ�;�7n��M[)�6 {��7ީ5�����{�v�\	Ã7[��
N6tw=���HICg,A"��@1i�Z������՘���d�]�O�U9�"���w�"��E�tAz�?�����]2�V"��!/.��v7n�)��e�'�AO(cv�������DbQe�ڷ7S��<�j������7�1l�B��L�D^��{8���ieF��8��1��NZV�|��VA�b�@�� z�� f�7nT�.�ڰZ������+������Yr�p��=D�`�1��Ŭ=�(P��A�b����c�:�R�6{3 n��?�c�;.ї���q֟��z �"�R���d�LV�<�Q��i�џ�M2�Sbt�#��0yI��:[y����QT�>:��� S'd�g�EByPz��b!~Kt�EˌS:Z�Tg��kB�����_7q"�`Ӗ"��S{	�蕿�_yxd�y�-Bׂnj�`� Յ �q�l�jQq`8�֔���u-��R�e����塲�݈�����1qi�����MkhE���5����y�Z	�Y�Z��H��}!�U�Y#��������'����n�������&Ef�E��2bIc�㛢�=u�n��S�r�%�7�;n���[i&6$�r�@���K̲�$�Gz�� f�КU��QZ��G�"JP=q��Z �Igg�If��oB��r�u"�=X�1XX4��)����|�4��r!3o���t���: Z ��IT�i
�(�|ڷ�!-f-<��4�+��t7�AI+������I���Z�#�ޟ$���!S�_ī�v�v!�0rviњ��#L��*�u��4����>?��0@�UIn�ώ!.=�-	jk����{P�
9XϾ�%��lK�3�Xq�}���g�iW���;�SH��(�
Pט�|ܶ�)���h������r��U��>�A�v΁U�\>��ğ��c�@v�Y����,��苆�Ҍ:�3>�/�#P��P�ѥo �՘i�g9�`�7�t���Q9؜�7Ue�\Ҧ�M&����*)�����t�_�Ӂ��eճ|*��7�"C6�G?Ud���K1��>�WzF��ۣ?�Lo�em;�-?�ED[ב�ЩuT��u�L�����93�ߘ`�A�馴��,+��^�]^�s5�jW�l����`v���9��Ii��X�:>� �+!��O�`�Zx���E-�+<����gԷk o)%R�˒�d�׊ZD�;��B�FŒoef��9���E��'5(�d�Z�sZ�*D�l������Q�GW��[�����\�� �8�	��,eB�g����Y��4Fa!�%�!e0��o�؁�B�.�9Sc?�3D�[��\�j��@�s ���?��Yh�m	�8[��� v�x\l��O5��vF��h.yi�����+�vY���wd��RP�5����f+ef^l�(��ݣ·�J'�	��sf�sT	LZ�=��e�!
tSa���e�.��`��	�q@�R���!vb7�l,� ��.Aɻ�6�:��,��y����v�e�[�|)�H;��x|���q�� �s�jH�M�42g�MÝ��(Rn�]d�7�b�@k��/I*SEc����%b�/�o|HInp,�w�����TH*Ce~��jC<y�v��Ʉ�Х�q�w�|�W-�t����Q�qdi����)�A�<���2�v_?5�HQ�4���0n#�o��<6�+$[,t�����q'e�<�*�M8����pΙ+���M��}_��<�5���F{°8���]�~���).��._�s㡻kU[��_���P��T�ߺw`�kb�>b��@��C)�^�M\C��T���J1�ɌpKޛ����zn��V�ؑ7��~���]��iFB"}�m�)�;,���L��M�
iܓ�ŏ�Z�F��+�]�X36�wя��`A�nk�F�ܓ���դ��m�wU�=����ţ�2x""��E���(;�ӛ�mh��2y��?���>� �G,`0ȗ�D���_�~Ԃ(����Tl[u�Y�G!�LM��R���<G!���踩TM��M���1�	?Z�}Fxs�!�L�fHE�q�rv���\���WQ��ħ�"�����v�N��fW�	r@�W*z�ZҷMDx6���2�p	���q-ݟ�q�a�
(b�OgC4�Y��>���v٧boΦ0�Z.0��b��l�4r�t)�i�����d����4�C����@<����R�J�Y�U��a	oNxQ-�TV)�w.z�7]��v�[�zQ���c�+�dw��}���"�(ޖ�G	G2pmNQ�x�c��hص���tT�=(��~ \p{���%w�	"a���tҫR)=�	�X:g2�"�_�o�$�l���-/�����{07�${C�E�V$C���iI���Y��`�-��$�ʽɤ�o���&�6�p~D7`߶|o񫊊6-=��/	"B��ˑ��̭j�~�7dc���[=�3���䉥yb#_��oP'=Hm�v�L��_��$������8�Kj��ɧ�52�5�EN2� ��j��w�4�v�� � �2�\3�K�D$�F�-����R����z&��1���z�YAYʽB�Ӣ��(1�i:+�M��>|��C�G�+Y�繞�:�+/���z7�3M�4TK���,�s(��H]��x@�Zj�6�3,�������ND?�]c��N�Sq@�?�e������_1�Ԛ5@{�5O�ka҂@��8w5޺2Z�Q�vmuc�����I�}pc
a}|"z�-3�9���&��2���,"RO�ĞapѢ�\�3�g�<A�;�}<��7���\���� �yU�zH���造�;�'���{:�5PLM��2�VW�]H[�9mǮb��~9�Dʢ�胋�\ں��q�;��)��<pm�ڢ4M_�PA���1S%z��
��M���	�k�J��A7�'�ɾ/J�z����ԡ�D^����m/KVX�!�Ee�4Ҿ��o�o�PK�H�C�h�|pR/��W�ա{���$"�EI�w%���ip�+����Ʋ�ޠ$�4��+&� ��}&J~ke߽�U]6�d ��)�B9����K���~�Ssc�%֐B�`����؋a�y��8�1d�PnG��[v�}���t����؁x�����jĳ���2��L<��=�j�WKw(z|v����-� Z;�2��1gD{�ٰ��Q��e��4=*��@j��x�V�Y�[��.���}$10�����;���rEG�.�Y�|���lU+�'ɪ�c3r��4����-�zS��/���;@s|��gf3��^��2���8DF>�J-*Nn3x@Q�e|��d�[1eD�F	�{��F��C�I������A����Ah�ق�އ	���2��UK,�n����\�M���9'szxt�>�>a���>�BG��#��\Iej��N�V��L�M
�KL�E�^(��[ZJ���N�ω3�,�`���R{��̻I�=�d�! �CM�黬~��u��c�`�娐]�ͨlH:(�K �/���{u҆:$�!G�FV��OZ��І�Nz?Ug����)m��6�\ ;e}��O�l�T�dš�#8�dm�)<@�꣤�\:���u����!�]h���|)�fBn[���$Bz*m��88��Q�Λ�Q��Z�������±��)�O��i��U���'h�D�=�X�@�.5EM�GT�yMj��K��5�o��nL�� خ��M�k*�8��j���5ҩ|K?�!�g��=�Z�����M�	�1xH�9����QR�
�ġ�Yi�j�V�� 5^�9G�?�ǑHj��]jctBr�fe0k~8l.����aS0���O��xɍ�ۣTkW��G�����]|?6�Ej$���Sx_X��Q��
�"ih"�Ұ������E}5�
)B���]�6��6��sqU� /7T
�@��Ú�,o�M7�%:�$�F�q=����^��
�H�t,y87ѡ��7_���S������`'��>>�5�3�J�{ӷ��Ԕ�φH��k\�{�E���^�q�p>y�oi��xX�:<%������5�����[X��M��hqr�dў�o:�9d���rS?P~3(g��T"�Mu:�vJ�v��L���կĔ��0��GS��猇�����Y�ta�5q"CM���l�9�a{&�­����?�0O �VaC�`���n3c/�/��;a�<k��)�l�p cxO)Y�H���s��;
XP�T�S�H��L�d#^V��*H�h�m����c��9E���'�f��rM�I'�������]��?$�p 	��G��?�z�{��SX�F����@��\ݑ����A�H��#�ɑ����i�w��zB�*�tm⑁Vk􉷸����,'�.���<�z@����V���;�VLh�Z��c���`fQ�:��(��x�C(Y�(�}z�J��<��]I��ҁBM;��[y?
��N��}E*�B�� O\��NLuuWE��DK
?�ow~��su�J��d�暈lH�W͢\����ˏT�]\1�8�򇭍d��n	��A���Dհ�V�I����1��v�2o�����h#�����T�����ɒ¹̎}�ɐ!,�]�։�:�_�`&?�=��=��٪�v�	��r^BYS����r�C�#8~� ��RW�@��frN�e�.�vG#���̌�u��0�?y�:C���P7��\PBZҸ��6JWq�8^��=�-&���9JN��C��u�k�[��$��s��t�	g&v�s>^�8[L�W(��nW?!!�2s^]��/f�ŊR��Ix)M��.�A���ڶ���pӡq�R�!�j�?8�MP�D]��[�%��'�]�k�%��<?89웆Ջ.�4�$XUe'�p3,�y�/��7��j��+j4>���5�^@��� ���Z��!	y�F���Ӏ�XR���f���$�B��Z�s��8�����c�EӴ��Wۯ,v`�4-�;~����z���m�K�L̑�z��v�>��BU� #�����z��t��ʆ�R��%�x�1�B�,��?�T1^�����;7��{Տ�d��7^��K' ���i��.*�����PAl�c.P������xWAWz�tiމ4��"�;��H�MO�C@_�D+�F���F�N��;'��%P�$���Cq��Ȝ�I��2OT*Y����^���P{�u���Rq�Ap<�������*j�ʧ�Ag�8���vBxx����p���@�6?#[t� ;o�%~���[����BZI��h��8���o��Q�J�(ϩ@�����uJ�8^�!%�B��ѳX41̷��xw"
cܫ��>���$^�#�C��?pC��<�D�Y����?J0�����֢�s�U�����t[Jl�[�Ƒ�p�҅��ZJ�{�W��V2"�_��y�³��Ww!�A$��?ÖӮl�l_��^U_E�,d�6���;��؋e92-��[0�l��,�n���e��H�QƟYe'{�9��a~#-���[�6�PC7@�|Oƣ�j�v��p`���Bj lǈ���D��ɈeX��$˧N�j��.�; *��Eq�ز����z���[a9���f4����}����)��HE<z����w>����+)$�ԉ�7��:ǞI��z��0P�X�*���GbրDԻ y9��f��E�A�.۞�#���2���)s��,��$:{l�T|���.�bc��@U�_<�1�YA)W�t{U; ���c�,�Ch7U�����U���;��v��x�y8k���A��e�U����' Ke&k�/��SQE���GB�q��Zm�+��<�76]�/h�4q�;��{�ɴe	=t���XI<���]C��u���X����U�;	�}?NX�'۽f�Z�c���䤒�Z^{�����o�����
@c�K�����rh��5�p�+d����i5���ȂX����]�J�=N+�W����<�����/3�\�a��J.y����\��[���E��E�ŏU��~x�ׯ��&�\(j�lq�=�2Xl���"I�u6��������_�buqi2M����CM�-�[4VK��L�X�]�� `����/!�XX�E��	�Kȶ=����ʭP\�;�%K�9f�x|X�7}��1��I��o�� F�Ҕ%>���˝�R�cj=���������#&���c�"�Ș?-�;�J[��!�Q�}�z\�����0�r_��%F�(�}�Dhf-�FǼA/�n�BM[��L�*H)^��x����0f�-yKE�x�F��P}�i��a����)@�8c�&5�L�M� ~�������l��nR{mX�K���@0���@���Rp��_�5�^ŷgO���s`N��m�,�K0�Ґ�tg�w�8[zgd9�l����G���NA�=� M�t9h�k�q*�q��Y�(��/%\�A�W/�o��/����r����δAz�Qպ�����6�(�5c��J��G�a�"m��C,��6�e��6}�(�&M��4�2Ң��>�c�qC�(ݺJy��.c��>��l�P�g'���?���3���s3��g�v�0�4�J���Ԫ3!a��`�����jʂd�0S �O#n�LMo�B6��n��QK�����{���p����N�x36����H���g@v���1}`��<�B�+��,�c�-&S]��i�X��v�����"^"݁�B��ӹ��3Qu]��J"�$�/�݋.�d}7 �+\�X�O<�&�!�ƛ��D�r�e�.�7�y<��T���Ke ����_�D��飣D�|>��}���oXo�E�b��Vd���
�b�<����h���z�Bxϰ�*Y����P���m��DLp�?�=�[;�E��@:�<ߗ��=��U���.P�N��RgR34�����;�O�����떕�ݟ�Bq ��R7b�$pd�6j芬���}���P��gp�60Byݫ=:o���o��Qh�>��i���{g�O9y�Ǝ�v `K�5&�Y�bS�АT{G���G���5�M�7���`g�E6�Sԡ���ԥ�81d�+�-��in~��`e�K�4�� �!Q�QӺj����-Q���y�������uwÈ��:�"��}��|��k|t{E*�5���*@�n�Y�N�\���*n4�i���H��C��Bj��h(nv��&����&Y��٥2v5r�w
��Q�xn���S�H���!�O��~i�i:���4B@�%�l��Gb��f��0���d��� �mZz��+0�"�[\�4�><"Z!bg�ilf�}oo�]5��u�"~�C�E��4Rk��D|>���]Mos�$t䐭���% "VI��
�#
|nz!A ��N�H�~֡�47�;�I�*�����y���?#�E�$�TEֵ^�s��F8�Į0|]ѮY#���7euz[�4/���P��>Sr�0�35U]��c�!B��k�i������C�R.z��5ק��X����I��}Uۜ�+;�r�S���>S�,����n�)�n�h-���`r��|�+D�U��vb��U�.>=����A�Ԫ��mb����H�{ً"ߌN��>9�o#dGXPDZ'o4w����m9�`&��������
���e69M�����п�)D�*����ȻT�[�ӕei�*�Ι7ș6ǟH?�2�����W&��Mg��S%�L��mO�?V�WD!�N����н/w�M3��`�L-�|��9�s�a�U�
�H�<@�Z4�^�����jk��@��t�~�,~��7��&��N� e!	��5��~x���E�3|P�x͋�^�= s%f0���c��!Z��,;��ͦnA���g�Q�!��ҧ�y�(�	sZ0���>~�lrl�&�ȴ"ڸ�[{ܧ�]���x{�8��8�>��5�B�Jƴ4�Y�{F��%o��u)o(�`�Og��B�BS��^�G�[}?�\������sv �?�r�h<�	���[Fe��kY��LlJa5Q�`vZ8hº��p�����Y%���P��f�75T�X�ݙo��(�O��e^� z3�K5�'�;����sh��C$=���h���a<�ˠ.k��=�z��;��.U�2a��%�"?Qv�IO׀�@��.U�|�V��:����V�s�(�vc��[�*1�ܫ���'Ѓ��q����=H;���c�0�Q���a�<����G��.�Gbi/���*�6Rwi��q�b�Z4oօn�l�wM#Z���*ל�����<S���Ԅ��;�ą�wr��|��	ɯ��}Q+2xԻ���a)��H���� �
�?I��Q�I;��ל#&���P�2+�bg,�\ަ�	Å�A�A>�8;�C   �   ލp�F˸�$�R=�1�#l����O�ToڬrN�'|W�DC�O���]�e�����:Vؽ�Da�w5,Qlڿ�M�F�ilZ���T/f�l����!��TI\&�L	���I!����һi7&�����o�x��f��T8���,O���bM�HR��V��x�Il���>yUJ^2_�Y�C�b|ެTf!m�04Jܴ�M���F}�*�K�	_�ts�\`�D97K�p��T��B�	5?��0�)Ҿ����6`�C�I�m�̵9��]�c�B�L���C䉹|�z���#CR����_8D��C����$h��ѻZ�\�)�Y E�C�I0<ĆDY�*]0�|9�)ˀm�2B�	�V� 4C�l��,ŌD3��!��B�IY �z�ꊘT�\h!���1ݰB�ɯ>�h$3�Ꚋ7��H��ZLB�I���I(�JX�t����`���C�ɖI��D`�YU��=��@ax���>	$EJ�AF�s��ʻN���QD����O4��V�d�27M>}b�ǚ�ug�O�� �J�-D�.ez�,/2�\�@��d��O��L�\�4ᐛ,5�șv薹���AC�>Q�1�S�#<Q4��-}���"��990m�g�<QP�I 2  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   5    މ04�̐��%�R(O5f��p��'l����I�l���   ��@ӌC�A+,ɘ�I'\	~�`%Ϲ>   �   ލp�F˸�$�B��>�1�#l����
�޴Y�:��O��d�����	�����"fŰu�pph��^�wS,�ش>G�6$}�8����
x��ј�R&?&����[���x`&�j�"<�C~�����Y,~(��v��e��W���%���36ڱ�-)?aQ�E��7Xp}BJ�8���D�5{>���N�!��X�Ӻi]�V�Ϟ������ē��.�-!�ph���Ȯ.��x�ȓ�V@".V�>��`���G@�ȓ]d|z�	�i.j�i$e��N9�ȓQ��
��p�GCO�kk�����ZG�<��"��(VX��N½,�V=�eH�<! ��/q��̂0�� n��iI@�<�P��i��`���?��%b���P�<��*�=E�2�:C�"�D@�0b�M�<���c�P�Cc٧o58L�1%Np�<I�"ϧ3��m��->n�a!��o�<���f���'$«h#�+WfD��h�'��Ň �¸��O�=y\������I"Qf�n�󦹤O��7����rX$��N�1^n��6bD�_��➀��I0��B �3b�F�d���
q�9�'t�Ex�}�'�R�j���2������6�|���'�L�k@ ��<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&�   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ����Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �   .    ލp�F˸��%�R(O5f��p"O��Q   �O4���k���W�ID�4��B��0<�bH�Q���   ;    މ04���R0�Q(O5f��p��'l��_��p>���   ����XѮ1�'T�����   �   ލp�F˸�,�p�&�1�#l���_�)��ToڬrN�'|W�DsĐ�M�� ����K�3세 t��7v��Dr��'���'���D8�J� �G�@gJ��s.�MŐ-���ɍEk��A�i��)Ё�J�h�!�)ԊK�=�-O����L&QHn`�w��DKr�3_��d�>1��� �*`�]/,�4��U���9�T�c�4�M˗
U?�V�|j6��X��S���}ȧ�+;n�"˅.:� hO����V�"o*�Y��:R`��FA!0!�DA��"��� �]�l��1k ^�<A�\�[�$�;���|����\�<�̂�y��!@L�W�����G�[�<�c�@�0!�Y�Z�*���&�\�<	 '��s5ΐ)&��y	��Ju��W�<A�+A�5Բ]��̔uH��R�'IR�<�T� t�I ��I� � �s�kZc�<������؀k"��/N�`tca�w�<�
�E�~�9�M�l���k�r���a3O���6)&�>4`�
͔/^��Y��H�n8��T��p�'�ܥ`K�H��뎍#FQ�����D�f*#�d������]��&�fx)w@�?;�h4�׵���'e�Fx��Ln�'��	�a�4�>��@�@UA�,��' ] @ ��т8#d�p�S�
�b�M��M�ax򠋄�?I�yrLV�7�|U`�!�9�� ��.�y�V9*8=0�#	,3� �H�����?�2�'PL1 b������h�N�MX���ҫl�����AC���j

G:Ÿ��[6R�u�������	0a��$ڣϒ/*0,lBE�¾l.�B�ITQVm)�D�w��ѐ&�~NC��-+�����(��[��s�+˿0K�C�I	\̀�'�.Y�XMH#$M�?��?��퓨)c�A� �Z�P���O�!!��ċqO��S�� ��z~�i�"�V�9b�A�]��L{����yBI�*.D�� #S��+�^�y"�� �k�ፇ6:���y��M	���D�%/��0�R��y2�Eyֲ��Ќ�25�p�%����L��(��)cL�*b�*E���"H`�3V�TsDK���\�)�3&.�p�_��PU�HݮB�Ɂ2�����e�*Y�@����O��C��sy�T棔(H���q�ːl.FC�IZީ1�f�,�[��ȯ(0C䉺I�
Ĩ��H? ̑�%J$!���O2lE~��M��~B   \    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�N�6��%{B,!�����`[�nA�`�D�>$�03C   ��4*�ب��P�R�B��eN�uR/�P���N�G(@��������� �5   �      "  �%   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=���w�TM�P������`ŌP_`��7ju�r�d�O���<�'�?)�/c��!���ki,<q��_�\�2��uE KH�	e��J8�(�Geب���4�V�U�XQy[1���h��H�j��ߥa&��[�2�8�wDCs��P 7&��<�Z1)��'?��o���$�<�����D�>)kE�f�0�"B��b��O�<!��*Z��H�Ձئ~2�j@AZ2[�'�7-����'� W�'=��B2�a���ن���ަ\�L<�媐ԟ4'�8��?5rCK~��'�J��5�X�w�^iB��!ː��	˓�����'�$n��d���p���B�c�ayB���?!���䕷!��8��C�k�X����7B���O���(�)���U��H�l׋���!@�ÝZ�@C�3UR6ٓ�i�G{��0W.�l��DP�h��� �?I� s�Ͽ{q!\G��j3D�z�bO�r�'Pa}�	Q%i�u�!΃+�P1J�,U��y"B �9jֈ��&`B�*S��yb $!Lt1�f';�5���G��yR�^4������_,Ā��o!O4�Dy�̱ Wl}Pg���мX��Z�nw�D6�D���S�� ��|}�a�s�eu�Ǳ ���u�L��'���"�@�h��pG��j�0��cl��j˒��>�TjX�hDe� ="$��ĺ8&�
���?���?��A��?�}��2���&#���8�R{d:���,CH!��K��dH�#B�F�L4��J7�r�����L�'��Ӗ�2�zuA7��=={��쐮�~b�'���'�ɧ�S?AuR�[%AB�%���w�>9��ؐ�9��"�nC tr�0D@%V���""G���B��!v�tQ`P�ʌ:�T�p�F��(P�d��O�����z�.�9IP�M���pi�9�!��ZQ�N-_����׎6WqO�lZv�ɰ~V�A9�4�?I�4�P4�ǡޙ@�%"�����b�'����I�|2���[�&,�g�I��X�¦����ʭlҤæ�0~>���
��F�<yC�I�V>tt��͒�'~����۶P��	�F=�=�/b
u��k�o�x�<�v�G̟��4�?��4}�`1�ļHe4xv���!!�'+��'��'y�O �'��I�ե�"p��wm�9  jy�	�'Z�g��H� �
� 1w�����R?y+Ol�[��Ao}"�'����mڢ �̽3vW#4���pQ���-b��?1a��5;7��#�:?�-2T�Z8��~���168�)g
�|��!Fs�.�D�( 
H2R2�Ar��7��c?Ń�,N�K= R���F���"�7�D�A��+r��5G�����A	��&Q�e��M�x;��8���SH<I �U�}�rTj��-n��� �,�q8�p1��d�lۤ! �h�U<���`�/]��
޴{��0���?�'�s�oZ�?}�	���ק� $��`%K�2��4�4b"�Ņ��(?V����V�<1tƏA3$��|&�$yu��6�p��C���J�pc΋G�(�H�Z��y"H��=8b?O*��F�=� �C�3]M`�p��b�7��My��	,�?ͧ�J�}R���>P�1�EP��Z(��C��y�@7t��ge�
G����ь��	�HO6��'��I�"��	xci -jH��u&�>4%v�'�*m�f�'R�|J~2�I��=��ܢ��\)HT��E�Q�<�u ȍJ����`^9��v�u�<y"��8�H)�%2 �(c��F�<a1J���0i�L�5g&�rt	\�<!�r�B��k_b�� ��PܓyΑ����k�O>�(CG��HґRW���N�@�:�П(%���)�gy�/�(#Zr�C��(`@H�g��y���'i�5#�.% ����T,���y�E��2�aڷ�y��<Y�O���yB�ݔ&� �)4oi�U�h
��Px"�U_:
5�#N^�I���u'z�E}RL���h�v5�#-
�a��;p%�.ITX�2i�0�I|X���D�n���[Gʅ���e>D�����A2�a5�K
e�rx1�6D�p�F�I�#�:��qdJIɚ3��2D�|s�	
�/�]H�@ʕd�D�sb6O@�Gy�/^��x�SAM!���ؐ�W�~2�#�O�i�O:���>����&i�5zЬX����H���<��A�7?��a�J�`4ĬPtg�|�<� dsi���'�>Ta���Sj�C�əXA��'6[y&�
������C�J���5��81(,ʶ
ʶT���'��#=�R"E��
�ʰ���)&�H��]���{���O��O�O\�%y��Tǫ�]�v��'�/D� 4жY�b��rMG7#q�q 5�8D�@����0�и׏ƹ��y�'9D�H���l.%�S�!�jup��#D��8B�
��DH�v�D5=J����"�I���O��S��'4x��ғ{C��X��b@��O��O���<	�Eں
T�������(�b��c�<y�)"yVD�ÅL�%�����]�<�Fj�v*N}��
f��c�X�<�Ef�x����*�
���D�T(<��Z;N��l;FE��5I�	H�(S��>s�I�Ow�	�T��Jp��֊�Iú��t�OX�%�O�|ZG1p� [V�"��"Ob�#PA	��BAT�bI,\��"O��3m�!?����A���9̺���"O�(2�0)k̤V�Y&\����'?Z�<��������=S�0u͓t?��!�`�����'�r\���!.���1�@۬\	Ty6�9D�����ؚk@vt�m΂�����9D�TIcG�Ku�HC��:~,n���9D�����HXz��4Q�袵�6D��{f(42
�ȸ�HNr�Dk3}�".�S�'J4|��bC�T*��#rhxA�Ox�R���MC����S�7%��4\ [�K�N-:
C䉢<�J��Q���F)@>��B�	7DʑH%�B/Q���E]�V�B�I>��y��6}�4۳g���"O�qB���1Va���l\2m1�m����FI�'d�h��h�X4���I�C�v��`Ŕ�w7��v�'�'6��Y��{���4xJ�S�K��c_R]*��/D�!�j����$Zf,���)D��i�$x�@�� -�gĲ	s�D(D�$S%��P�:V��S
�A�"�"�T�UaN+��۱��XR>	IV�(a�Q�HI'�5�'|=��h��CsR� ��G��2*����'>"֧� �ЋG��s���f���0P� "O$����37f��,]=F:�h "O|u{燚7H3����'9߼a��"Or����25ք���Oۚن�Ʉ�'4*�<1�T��	��C9{��K�B�~?yp��I�����'��S��I�a_��ޜ��-�2��1D����s��0��F4T���P2�/D�d�p�T�a�H�k5ÆF�n)�AO2D��L�5F"1�RE>~d��;D�� ��� ���V �&
�=��+.}�B?�S��3�PA�`6�9H�� |ؚ��Oإ�g�Op�?����J�@�T����T�n�m#�ƍ�y�iR�t�6]C&I�(:�*,ӣɫ�y�ϝ3Z���	$�5��ಒ^��yb���P+e�M�3��J�j�y�gQ�N����8� �%A��'�#?�������Z�IP�&^�+�@�P%�Q���?�J>Y�S����%k0�2D�J3:�� 6G�-OP!���p��X�Fԏ>���e�6u6!��K�#8�`'/�_D������!��/m���iL�.b�����&"���R�6�P�����22�#Wn����ο��>Հ�n�5K7j�C�ɦ0�(����K��?�����>�4��I���)E�M�|9�VZ�<��%R!i6� KÃQ&e�Э�oV�<�0���!㩖#C��L; �ZG�<&��7)v���LUD�C�k�Z8�X#���҅h[�-�%�4��|V�6�����n���Ο��	W}b�Y/ZԠ��bC���!�tG�4�y��F��\i���3�%�%;�y"��5?zP	2d�P#9R�/�y�gL�n��܃1,X0�4��Nڠ�yR#4p4 ����'{����I���I�HO�r!���L!4ȣ�Ki��1q3�>i���)�?a���S�ӏ��@I�I�0=�Q��,��d�HC�	�M����� #a�U� g�qz&C�Ʌ.8ɲ�GB%2f`���ԇ��B�ɞG��A�(G=TK��Y秐]�C�	�c�F@١Fގ`�z-��͂i�㞜����E��jEaD�as��
&*d� 3�J!c���$;���O>�/꘸ b�>fylq"�4g*��Nz��uB�p��,��(M������)�#�ҿ�� ֬�
v��D�ȓ>�p]8%�#Xt�����xk�G.l0�	��aQE鈔s]�
E�;�e=E���8O�y��"à��eA�9"�d�O��D���j(�% b�h��k[0S!�$�)h,�&��@N���7���&�!�X	c�`􀙕=/�L��"�!�T5Z��tS���B#
3�>k�'"�<��U�!�fXR� �E�9
�.J?	�,MU�����'��_�К��.[3L���O5TA�d?D�p�b/�8�
}��擻(� ���0D��@���&O�p �
d��[�"D���Q,֜8��!H�>g�|qڦ?D�$���ٖ�t�)�(0� 2��=}"�-�S�'#�\9��F�5(�D���>��ؤO�t�$�O\��2���t&ĥVI9gO�YILi��C��y�e͋@����Cf�0y	� @��y��< �>�	ăm�v�R@�=�y"HX���u)�7T��pÌ$�y2���da��@l�1V�D|�Љ�'�@#?�rh�$GF1������d:�ԋR]��?�K>��S���?k�1#�a87`����'�!�� 2��Ec��,̚�)$ӽ`QT�3�"OYb��ȢiE�X"�Ô>NMB�k�"O�v�∐z���SΈ�A
O��8��ʸph�ڄ����湨AZ�ƨOVq ��S�.������39T8��*�!sߺ�����?��׀�Ja�B�W���v�v�C�I�P��,)�)X ��"R�QS�BC�.!h���`))^����5�Ђo:@C��+젽b��\�f����ȑ0t��d�p�'���
]�RdZY2&�	�OC,%��'lhٌ�4�X���O�!�F��'lܞb;�<��"Z;E��ȓdH��$�Nd�NT��慟/0�ȓOS������Q&���CCV�0J8�ȓA��1r2 ʃK-�� A0��B�ɣbF���	�������D���'�"=�BU	8[ƤQ�o�"4h+��}�� �	�$�d�O��O�OӺ�E��;M�@u@>cA�\
�'Kp���%�%m��(�Tj�:%6���'Cl\�)�/*�-��B�M����'iL�a�L��Zo��C�`�u�a�<��dēIBb��,��Y�u[��W�S����J�O�E�uBC�(�*�@�&�N���P�%]ܟd&���)�gyBi�'��-D?&ɲ���Պ�yB�̸D��dAÅْ+�SQ}�C�ɖ �6P�Ǣ�]�t��7�҈uzC�	'�]3�&�=%u~Z�,�<q�.B�I, ���ˁ�T�'.�X�CA�tmv����	c��}��$G�L�YS��&	� j��jI"�'�a}2��q���kA0Psjd��+��y���J!�2iʯ|,�%a"�'�y�l[�!�v�ʰ����y��[�������Тd��C:�p<9���{�N�	@!.^F$��jÐe2 �Ƀ7��"<ͧ�?�����dU�N� �)�Ψ|���_~�+�'���@Ĩ��8_4�X�-��f����	�'$V<qV �3*���p��(\����	�'�X� S�����W�P.z%9�'��u�XeU��[6�Y�\j����<}B�/�S��=�H�6DXN�@P�N p���OD|[!l�O ��0����J7���R�X
	��ty�@�#�y"�I�`�/�Vu�E!��G4�y¢��e�X���+�6Kf���c�y"�X.@��E��;���6h��y��A:
a&���_�P*4�ekF:�'��#?af��ɟ<`���Ji��,)��hd��0v���Ia���"|�' i*p,@&3���ꊏG )��'' ��Z���T��!)��8�',2�8�$�-m�鉁H.s�����'�`�Z�� 5xI����.?�����'O��C�'�j����S��5���A�'K2,���)N���Q�@�!7��JJ-��`�	ן��	�XX��ɇ�'j4Z����u��C�Ɂ�<�!F8k�Б
��xF�C�	�B��ä`ζxI!٣EY	߀C�ɴ<�Ԉ�b�6;��`D�[�p2F���t�'@�s2�� �V�8c�_;aY��'�ˈ�4�T���O��W[$-�T$�� j*�p�E��$w 5�ȓ#�̈��#	7A�b��C�L7� x��
�%*�d��'LpC��@�n(����D|���B�K��"'%�!��x��=�v�J��i�0�ӥO٬��O؜Gz�����S���e%I>y?��[�����-���	ǟ�%���X@�ݢD�� ���PJ�"Or�B�^�R��u���a"O� J�����=�vBO�G�Dxip"OT�Y��g����0B*V� �"O�z�� #:��r��5B��H���^�'ά���	�����.��	����&qp�p!p�'��'q��Y�8� �wt�:�*�	-?
� � <D�pP-��ufK�J^��L@��.D���3	��)��(޷-4�0 ֪ D���(�M�:��Q'�[�廠�2��Bа,L|���
�Mi�P	F��Q��05+8�'44�m�#��+��(�V���C�I@S�'bB�'��}H�e�Tu&�)'���&*���'��Di$'��H�	@د$*�{�'��yЇL�'cE$����Z� yd��
�'.�u:�bىC�q7�­G��h��Q�t�p$������I.�J���lV�<I�#�E~2iW�I�Ox�d�>1§[$7l��J�擄R2��q��	3v�2���5��$�-�F�~&�E�����Ko�'Sh��#�M�f��c�KS�C���C2=b?OXh�)���arX�P%d���O ɟ`�'�L�j��|J��d�y���sr��%iö=���� �!��
]L����.�:ы�/حe*�_����S����'�\�$&#z��Į[v,p �^H]�D6����O��O�4����dfCR��tm��|�֬��c�{vX@B"�|����ϓSg�)����+\��1�P�ҋn�&��2"�Xgl �&�T
;���ϓ[dȜ�\��M�G���� �ׁ������X�'a�OuAѫ3��l��q0	{d�<D���7�F�=�:̋���d��L�4f=��M����ā�4`h<mN,)o�dƈhB����HP��xP��>]������d�OV��s>-r�� �L 2�	���c̶9q�0��Z-)���9e����<qS�Ѯl>N��p�E��(� �na)sfP3V$�u;'� Gay�d� �?�����[�acy1���V@p���HB
}'qO���%,OV��VIߺ@s�p�ҡ�T�&��
O��d�^4iw�%��C��BA�UL#V���d6�	-#|�ݟ?1l]��D���z�$ޯ�*����?���P�:��׵N3�EԂSv���FJ��y�E�sG&�I�JͿH��ȓ�����T"RJ�yɆ��:'N��ȓ{��z���� �:���5)ְ��ɝ�(O����)p��DR�U�U�X� S�O�|0��i>A�I����'0����,
l�� a�f]��'�Jc_i�q�Q-`��)�'���;�P:�L|�ШB�X�*t�
�'zzհu��(H��5Mj��Z
�'8��3f�{���&zw�I�I��0���霴_�.�*Bǉ�!H �e�� U�t��m��?N>%?E���<YS�8��'�~�0�ٗ&D�X�0���ed�l�2�� A�+!��j4X�h��Q�h��-Y�`�!�$Z�KV�0g�MtǺa!�D))�!��T�`'r0(êDod�H���� �qOZD~�o��?i�S�W�d�� 
�-C�Z�)p,ܹf���|b����I�JKZi%l�
wReC���9��B�a�@�BZer�c#J�Kj�B�I�J���/��y0��0�½R��B�ɳ �����֊�\�Za�Z*m>Bቿ���¡B�IG�I�O�)��ya�ɕc�j�}��hT�J���;�&��-�;�.ܗl�R�'{a}R��34�L�ZQg��g��e�ؠ�yE�c�����X�Yj��]�n`�ȓ ��U�v���d�\�1E�+	v��ȓZh�|�	-��@r�E)�Ʌ�ə�(O�<1슝�.IQ�(�5��	��"O�ɺ@  ���gθ(CmN��y��N�5��9P����i�Eϝ�y��_)��-yŋ��J��Ò��y�A�4L�#�ܝ�� ��y�F|�u� ��t�T0R,ۊ�y'� ���)n�%r�9q톦�y2 �:6�up�/lc HBa&�$�y2)�.Vv@�F��-~�Z����y�B�(~�xCT��xy����#8�yB�=�"m�w�*_՜ȋa� �y2�Y�gO�\Y�j�Y�J�@H���ya�>{ؽ���'�A)0��y��7�j�q�kO�J?�`t�
��y�B���@ D��:20ś mM��y��!����f��+:`�I�gG�y�&��,�bE�w��05t�;�]��yR(U*�D�eO:u�1��#�y�k�3(������'J9:���y�E!ɪ�`U{���CO��y�!���̚��	t�|@��M��y"-ϻ"����b��X�>�顈���y�OW�^���P�o�:GR�Hi4F��yB���>�ʤ��,�4B�h��"��yB���� xF%6�B	�Ʀ���y
� ���v�Ę�B$�ԥ)�f�@�"OVi8 ��6pR�K�>2���i"O�I���F�,�l8�c�:|�p@R"O�8� i�.x��i�X�b�
�"O���2W���W�M�(@X�P"O6	z�
9\��ZP��$K:�}
�"O�m"��Ȼe���"�)d{�Ԃ�"OjWnڞ �#0�ҵudvHs�"O��A��֘;
ȡO�zD0Q��"O����!W�\;�MS!D2���"Op�l0"���1��O M�~ �"O� ��2H9���89�ԐSf"O��)b�W��0X�Bk�7,�
�s�"O|P3����������O�R���"Oru��*�zP�<�
�&tEJ5�"OPd1�N�w�J�ǋD���u"OP0�D6E��!Rċ!i�f"O<��'�ر{�Ђڰ
�mK5"O\L�B�J�sp��VK��t�hm"O�� ��!{z��SJ[�v1�	b3"O.��SJٰ䥸�nĂ(:�"O��ࣦ(H�V<x��V�xU"Oj 0��λkچ�ɦl�6;� 4�"O氉 �Al����4kN�S_�a"O�M�V�Ҟs��T��W8YAK "O$L�o҂x�6��〙I�1ڄ"O��ѕHh��0���ķh�N5��"O�U��a�"D����ˉ$_��P�"O�`�	ܴ=�ʳ�L#\��]�3"OT��F�+�)��l�*�"O��6+Kw���0�٬�x���"O>��q�.�p�+5��?�~ݛv"O`q�`W<<�l���>`�ZX:�"O`a(��=y����D#&����"O8|�ׯ� I���ڠ�V�?���8�"O�T�P_��"���0k���v"O����[L���1f��a�"O����+��M��895�y6Ʃ`�"O�J4h��n��AP�c�`'�Q"O�q
��֯Rv�|�g���"O���� ۳v�,,{�Y�R�8�"O�Ö�����8T$*����"O�\�d��L��l1�d�>Vh�]k7"O��@K�<k��a$D�-EVD��"Oؠ; �?��,Ţ��+D�j "O���F��X}4�H��<v%��c0"OLl�ueS9F���RkA�D0�;�"O��aF���LU�L���<^��p"O��0��W�?$4���+Ѣ=�BP��"O�D�s/9$Z���%��q�ݛ0"O2H[�b? �j�;�&�Lmh#�"O��"g�Lˆ #�CO.\N�;F"O��)�d�*J�tAT�ZgF���"OJ�I��C�6�Pxه��}8
��g"OTZP��)h&��o̱)�4ằ"OuX��/Ww��(� ��>�P�Ib"Ox����,.pP`�� Ա"O�-�G��+��"��[�ԕhW"O�\�����~�8=J�J�(0�Tѣ"O��K%��z�zD���N(���"O�L�p�)!0VA�Dh��-4"Ox=�Q�N����RG?ZK�Ч"O�qhVI\�R*J�buE��$Ap�ڡ"O(A�`������S��`�`"O� �Y{&aO�F��(��ԩF���A'"O`��TD�1qfxY{'��Z�1�%"O�T�e9J�vi�g5<��=��"O��"A���S`d�bd`�XWB�#%"O`Q�N�I+���hF�1��峓"O�Xx�+��q�@<��GZ�J�,�"O����-�J�65��� "|x4(�"O�< M	;9�̙��Q j:0�2"O��p ��\�����)/��@�"OFij��� %|!���X"�Db"O� ��J�^)JP�e��+�h@%"O>�4�SP�ᚷ���I�p%S�"O�q�WDQ9K�p�DeQ29 ���R"O �jDB�-ɳ���7����f"O��+�2�0	��V$	��0��"Ox|ZҤ�R��"�a�#�l�۰"O~�Ј��@Hk���7�D���"Oȵ��܇o� q��/�_���I�"O&��D���!�|AC�8��u�"O��p�ѫ.~��2�N�%{v�;�"O:�3 �)!𨫲��0z]�"Ot5SHF'jޠA�D�l�ж"O0 g�m�n�0T"�8r��ur"O�Q����V�Y�$k�:a�tL�"O�iS�ڈ&� hr2�H�V�B��p"Of$�LP�"�v}dL�
{���"O�&n��e��(�G�Y�	µ"O�D����;|Nq��&��Sq"OҘВB��/��u��F�<|y�"O`��s���/·>��7"O4D���5J�x�0�`��_���v"O�c��� ��S m�}�@Q��"O�����QHhJ�#�e�.�� c"Ob�CeA�!�2��F��F�: ��"O&�)�"�r\0�[�d���Щ�"O�p�3��?<d,��D
!F��x�"O��N�,��lp��R%s!�\p�"Of�:Q ˙;-Z�7�_%�cb"O:܂S�ɷ]�w ^�$D�X!"O�,�C	��>�� �IL��P��"OD���L�Q&��0F� S$"O��ӄF(&�uȦ�����z`"O��q�'fU�#����� �"O~��g�\���ӂ7��;�"O4��¹��)r�! }h��G"O�I���G�r���h^��"O��)H��5c7/�S&�A��"OV���A!*\��6�MzyP��p"O�E�s�Ϊ3͜�*��ݕsr�y��"O������0$���R�=({.�P"O�`�q�֝u�Y�2G��Dz�(�"O�����u��"aM�w��}��"O|���m+1���)uZ��ei"O<D��aϋ�a���G�Xq�G"O���k�N22ǈ��+�"Ot��3ʐ2&�䐣���"`����t"O6�xѭ�0K�.IS�/E�)�hp"����zt��͛N5YvM�^i�'�����[l��E�B�N)�'��g�*ZV^���\&|�X`8�'�ܝ�ơ/t
=�c�߮!����'��`�3�e@L��"n�i�X�'B���t��=W���#aoG�
G��	�'��M!�"ПLN��0�>L`����'�����	o_�{�.ԏE���p	��� �T�4搥!��Q��='z!�P"OR������kH����>3|f�pR"O�]���S�.�>���"Άdl w"OBx+���U��dK�2PT#"O`)B���UM<u��ȓ�1J��ɕ"O `�/��y`����|��"OL�������bv
�m�dt �"O�M�A���"�pJ�&	���"O��SEFN'�Ը��c�a�:�P�"O(�2e/՝
�,�r�kP��b$"O�4�S"Ӂgd�ٙ���unt�"O�u���E=Y��o1p�-�"OjPX�h�-\��]��i�@O -�'"O~���*E�W�di��/X�6D�a1&"O��h5�ؐ?�zՎ��\�r�� "Oq0���"p<� �������Id"O��+0,��i.��Z"E ���@R0"O,����!7�\<��AB�u���""O��(�KÙ[�fQ�R.\33���"O~�z4�?S���c�+�$lj8�U"OV1�à��x\!%�#1��A�"O6��_&s#B�u��6�"OZUJ�`J��tAk�F@�Mp]��'sj,��b�,Xb�yjg,ߖt^�Y��'��X�����Z���
�LB�~;r� �'���a�lҨSq^��q$ÈHiLPa�'�)Z�hP����4���.!@��'�����њhQP�2����'�t�)D�Hj�%�s��7*c.l)�'.TtS!̢ɺ J%
\q�'A��s��A%B�ATj�.��a:�'̩C��t���┫�� ]�,�	�'`��ǂæ5�����W�.P4�I�'��Lծ�;�9!I�)[(@�'���!���FgB�|�j�'f��+/̥VjX3�#�9�P���'�<��C�_�x���gĴB�L�'�8�@T/:�D���.�K�Py�'4Π# BѠ��Q�C��-0=��'&��1����oI�%�Ȑv]��'za�	�ZfB�����|��'���B�"DL�9ϗ�M.$;�'w���Ứy��С挒q��r�'�ZMyƃ�O���a`XY��T�
�'
�	�q�Q6�bq@�Z�[:���'A�e���<����3���pX��'���F�D����2(�*=-h��'����" R'N���B�7�l��'���CM�8���+A*�%
�'5��AC �/\uh�#Wo����'G���N�>jװ�4��k���S�'�\� �ZC��-�h����'�b]ص��z��k��ϓc�f��'��)!�dG25�=R���4\Z�'����RH�4l'($A��S�"��:�'�`�A�'ϻ}(��4!��LBI1	�'i�*�W.;�:%#�G
.H�r��'��a���	!d�Pr Ʉ�ډ��'��u��&�)a���ʆC�kf���'l���G	[�=���ڑk�2�n(��'N:�y�	"���B%s'&�k�'��	�2م	�P��p�^��X
�'&pyO� �"]�!��H�����'T~<�Ύ�/{"-t�U{��(���� tlu�L3q{b�#Q�@b�2"O���Ưv}4YB�k��
M�)�"O�� ��	4�>�EhM�y@�m[�'XV4XtE�2c�;�EC�_�fIy�'�� �鍲K+\�@�]�
<��'*I#�T���V(2M�2)�
�'Z�b �?�8f�V�Kj\j
�'�:mH&�M�xy���߼RP�u��'B���W��j1lLm�E�'QșQ皈R�vY 1d��.��ap�'~&i��,��ԑSuF��-��J�'���!]);��Q�']

�	�'}Ԑ�����@�`�aԋP�a����'ȡ��N��%�GmZ'`����'yؼk@H
�1�`-Br��8�{	�'E�ٸ���"�M[%��.ZJ��	�'�"`�Q�[	j+�� ���"AH�!�	�'� �HB�)<y�@�W�7A�Dlj
�'�jq�kY9$�(���̗v�$�' l�rO�&-|����A�;h��s�'�Aȷ��7utB�!!�ܞ,�$�@�'���C��^�~�H�bJ�$SF���'���i��_Z��� ��*/�v]+�'~����A6� h{ B�p��)��'ڪ��]6�"�X�ϋ3@��'��[P�T�s�	sǊ]�4t{�'2H1s��A��qҫ�*Sg��	�'Iܩ��_N�xy�'@HE���
�'ۜ�;d�y�\49 B�0}��
�'�9� f[i��M0e_;dxP,3	�'2����	F�8��B,U��|	�'42 ��TÚ�SE�Ɣ
d� �'w�P'%Ƀs��|�g��9�eB�'�
��
�I3@<�I-��a��'��Œ�JQ��`C�1[�L�[�'�xa�5��t�D���^?%G��y
�'��b5K\�5������#l�$��'{��9��'�z�+ �Ȅ:5�e9�'�����h	I!~9p#$�03�%��'��\�����}۲ˇC�_���'�܍��h�{場�WLėPǶq��'#:l��u*oޫ2�XE�	�'T����o׌$��'R�*���X	�'ǆ�Y�KȳXdlU(�`ɺ%�����'���0&b<h��ㄜ�"�ݛ�'x������?d�R��e�H�@���']��bǁ��E���Zb�����	�'��2���z�0�T�P�W�Ż	�'HT�A���*WH�t��R�I�~���' ̬���K1LĞIITf��}M4���'s<�rk��a��Y�ǥ�@�4A�'�@P�N_+F��F�7A����'|XA�\%9�|�Q�ͳu{z���'5<H"�	C�!I2� oSԬ8�'�H��擆-8ƴ{�΀�l��%��'������م���nD�`�~�:�'�u��'�E��mRR���l�'Ih,�Rj��S�)��D9}G��'k�īSl�(b:�)���:�8)��'��4��Ԁ#8�1�b��N��1�'��K�84 �E`�$ۮN����"Ol�q�čGv0��ʆ� � Qc$"Of�!H���	p�䅟Y�
�!0"Or}�7!�Hg�c���2��}A�"O� b�[P�
8x���ʡ!�+X�^� &"O�%�!���xl�S+˶D3��5"O��$�3f�䪰��Q$:�p�"On-b�L�"�*P����q6H\P�"O���e!��az@�Ŏ/"�H�F"O��Q�E�8���2��ز9��"O���F� /%C����ސO��zf"O2�J�.@��J�1�Q�l�B�"O4� ǋ3Y׺����Q#t���"O���Qʎ�(��� '��~~�8D"O��:3 X�%˸��P₄u4���"O�pR�Ɠ(p�����>6i���"O(��`��&a�J�St�Ҙ#�Nxx$"O��b�G�	Y��Y#I
4�V�Q"OFi��/$m�#Q�&�B�z�"O8�80i5G������Z���"OJ���'Y�5vRp�2��;w�x��"O�e�w��s4ʩh���7j`�y�"Odh���O�XheC%��f�Rq"O���N�V��ʂ"C�J8�8�"O��0J¦H���T) ��(;c"Od����[?&��Dt�-,�����"O��YSG�3�@ڕ��!8Q^�r�"OR\�"j�!Ǻ	F�Y�p�pm�d"Ol�CF��>�ĉ�a��4^nB2"OV�@��A=Uq�iu'K)x��d"O^�h�2��hs�fL4_A���"O���4�V�Sp�T�EE�pm��"O޵�W�H�>���ۀA�]���"O�`XfG�=�
�Co_�Y��(1�"O~��U��6_  �,��~V�"O��s!��'��<Yc�M�Q �"O؈(M�=��Pea�<+�!��"ObH@u��$V�xѩ��&uDp��"OT�B��	N�|��N�O~�	�"O��外�S�֙6�SPK�Ѓ"O4�x��;y�&�B�d��5���"Or
��"^�H,��E�.~��`�"O~�5��6d�Ѐ��[�ʥk"O�d�Qa��S��yP��'���Q�"O(��Ė!!!Rͻ�A�s�:�r@"O�p�@J�l�*Y��/�
����"O�q�����A��&&��e��"O��7M�,�p���E�p�D0��"O,�%&
�4�Xd� �U�.�&�j1"O�E�Ŭ��S��� G_E�~�YR"O��Q.�%�n�8"�Q�o�Ƽ��"O� �eڇr�~���� =��C�"O����ޫ'����"O:v:&�Q�"O���UH��WB��tD�)H$�4�"O��H�W�@��K�/D�=p5"O�����L 2aI
��<�|m��"O��y@��s��!`�(e���3�"O>(2H�)��L��B4O�Ҭh�"OҌ���B�PI9!,=Hoef"O�0W䛀H�F�Pp@�ZZ���3"O�m;���+[�B�s�kU�T����"O"�� ��ԘZ�*��L�ٗ"OtɁ�mM�rM(%* ol,Ȉ�"O �������@Fׯ	���;%"Ox(�0���"�4];@���;��������o�l���G�!�4x���"��'�LmS�դ�05BA+I��ح�
�'�j����W�Z���BG����'��x)�"��;'P�1���?'�h��� �jŹlΰ��!�I;@W��v"O�m�d̙!<NAp��:Fv)��"ONp��.�!7���9E!ج�0�e"Opp����r���4��s"��P�"O����i��\!���TH�+r�]k�"O��	B�*ph!G�}�u�"O⩛���w��8��]	�ĸ"O��[�BX��Ph�$�m�0��3"Ot�V�C�(P]�Bc�c���1r"O�����[���Q"��dxڈ"d"O�$sыIg��`��=
d��B�"O\Q$��2D� i ��.pZ�R�"O^U�"K�u��P�� BX�`"OZ��wR�6�Ƀ'#B&AZf"O^�ك�b�b@�#!
�'+0��"Oʌ�b��8�$��> ���"O�]�@�#/(P0�:8�0Q�R"O������*��|���X�9:�"O���/�� �V�1C"O4�)��n�[�`EmS��xQ"O�:� ��j�<<���#�嚅"O%Ň�89EM\�r���@�"Oq�bZ./[�HA��R�XA��"O��yH'W�|2F�^,�Yڶ"O$A��/3��4�7㑦j��""O�Ջ�N,l��G��u0i�U"O��҂�6NX�gAC-M$<�!"O�u+#Q8$��p�Q*ZN���"O��)��ň�!�GW �iS"O&�jvf�'EXx��L�s$T5��"O�X�!��е����;x)�A3�"O@���'hE�t:��7J#�IH�"Ot���N�IQD��$��m
�$�1"O*t�5�	7|z�Ű�����$"O|���D͍B�b0�ւZ,<�M�q"O&ũ�؇m�|�$@�Ht��"O����cx#P!H��� t%{q"O�P�է�)V1�C"0����"O
�!�O:A5N�L��A ��d�<�ERZo��e��)@(<�`�b�<����2ѦA�gȁ;N/�d�E�F^�<����-Y0�����EH�öM`�<Iw�Yw� �
1��Z����d�[�<ّ�Z�j���&0�b7i~�<ID6
����DEɤ
��q㦝z�<yE;/�T�i�$��}Ԩ�I�E�]�<q%kL&Jcց�Y�L����[D�<�"
�4"X�Yb�Oӄ����c�u�<��=tļZe��>p�I�[X�<A̫Yx�5���/k�M��*V�<�O�0"��]�&��eHAi7!�T�<���� 4�ݠE̡N��5��F�<�ShE�n_�
%�6
|�{d�k�<qюD��D����\�F�:�'�d�<1 ����9�X4�bС���k�'Q?
�)I(=�`ЪL�
aPz���=D����Ȳ�|9�4
�6+�9�$�;D�PK��<�"|s¤ƴ$�x�@d�?D�@r�gP�qUr4$�`������;D�	�f��`�)�(J���15F;D�h h�W>p�+S+O���y4�:D���)��
m�&�ÀYU�|��h;D�̘�oC>��ӕ�^���h��&D��y�.L�w��S,-��1Ҭ&D�� @�CGΒ>���T�G-i��"O$͂���z5���H9�"O�9��U1GS<|��`�7i��q�"O� ���Ha��K֏��}	�4k%"O����:3�H����"����p"O��"R>C���x#�!Dʎ���"O� A4iɱ��=�u#�f���H�"OLt���M"dy�A��hP!�h%!�"Ob`�w�@&�$ �5��5Z8����"O��c�/�.�bH;�/�!S�`bP"O�q*��,q�`Ccn�LCPI�"OQ�U'�,#��(�!��G��v"OT��TdŲM���r0��B��[�"O$)�3���q��,y�@��pC��u"O��`�#|b��/��N�Xp"OT�j&/G)5��a$NT�$h�j�"OD�� nȥYT���r�Y�k!�t�"ONe�+�#)<�1� .<�8��"O֨���Jш�����T怢4"Ov���$މ?���[�$O�,m��"O���t�fj�4�a�J8�hd"�"O�K�^�o
�ͫ��HUu���"O:�b$�ƥXC	ԅ s|�+�"O�	���Ul�)��G�MpL0�"O���B�2�b%���Ū]T�ّ"O��Ê�h��zeʑ�qW�Ū'"O��+'�F�t?�p��k��I�Z�;f"O�`����f�(�k�'ОZ7����"O~$H�-ÒFN��fD2Y;t��"O�*bgZ�#eb�S���s�:��"O0equ	Ku��(��P�,�� �"O"�����(�Eт	[��"O� '/\���90tA[9$yʔ�V"O�3��%[�� C@�g`���"OE���C-h�183*;_�1��"O�Lj�n�:��x�5�e?�U�""O��Ȳ�K�yL�
I��5ȸy�"O�)x'Fɛ`R\�h���V5����"O�X�1�N�\���B��G>�	�B"O� �r!ؤ���nt�"O��Q��F��y��

VP�!�"O��YbO]�|,��;�G�]8��Zp"O��pB/rC*c@�j�||��"O�YeIY0C��lx����$<�c�"O��0��KU��U��)1�\+"OmY�^᠔��хh��1�"O�.-�>��ӯ�OP:u"����Py"�ց-�j����
E�b�Q��KZ�<I�-s}�}�D�]��p���V�<�6CQ�;l�У��+~6�0�jYi�<i�g]�K{F�X���[��-Z�<� L= �lQcs#��:���ѵlXQ�<�0(#b8�X��aX $ìzr�_T�<�A,�K���Ҡ]�) �Y6j�P�<��F��Px�y!M�Y`��N�M�<Y�͆M��$��U���+��1D���s�F��ˢ�Ӭj�ȘR�a5D��� ުw� 񂄍Тi���kw�6D�:�g�vhLŘe���fc� ��9D���Ɔ��~�C�'s�Uː���yr�%�:T�T �&S,B�@�W�yr���V]ա3�,_� )�Ŏ�y�U1�6��f�*{����G�7�y�*�dxi��9ykv���M �y
� �}�r�32L~)�+��+9֩s�"O�X�eaC�*S������-J.t�!W"O8iXt]�R�2�R�)�����ac"O�0��DP����"o_L���"O�Q�F�/J�f)S'�4Lvh�if"O�y���D��|���T#qj�أ"Oh� &��jU�:A�� Ag�x��"O���E��}�# �2G�*�B�"O�+V�$ ����3��d�`"O���I|"p�5M$1�*d(T"OV���� )��1��)�*��"O�I ����.�2 +S�V��Yx4"O.|S!�E+b���1ʋq�t�*5"O6�k�ُ,�F@�R/D�&����"O|ԙSlO�oB9aڅ8�ZP)�"O�JTIU�@�����`F�p-�y�3"O����ھ�\���aC�(/0��&"Olժ�ӾQ���2��],��H�"Opd��@�l�%)� ��!:��"O�j��@g�`�ѧ���QPz�#�"O�E7��Ba�	!�Ղ����hL!�ğ&?צ�w�Tz��	d�S�`�!�Ro�^���A�=d�p9SaO?.I!�$֑"���A�Y2)ZU���Q$?!�D@=l�d��R.. ���cD�!X�!�մ�H����W�f�r�ā=S�!�Da4YٵBW�C�2���d
<�!�Ĕ��0�-��0����}!�ߦ ��� gɑ!��XD��2!�!��+-�����=$o�D�t&�:�!�$�t�j���&K>cM�!���@��!�:pk���SK��H��#��<!X!��RA�$��S�PM�T����-y%!�D�C/
�@	�-!�H��/!�d��B�pZ"JՕ:�k��(j!�Ĉw �����\�|@��P?$!�;}Rp	��>8-��SEN�T�!�ď<^��1�ȟR*v�y�C��%[!�d� b;��B��8.1b��O�!��1H8)�b ��rWk�59!�ڴv/\]qE�F�!ZR�qEH[�I1!򤂟g�A��L> A�Hz2g��3<!��>�Z�����<=0�ك��}4!�$-2l��Fk�$,��	��'!�[$�\�p#״<�xB�Е)!��g���آhƞ7�4ٱ�D
!�$�4Xޠ�Z�M�j޸��"ə'�!��C�3�Tx���+���v`�	,u!�$VXQp ��ER�I~�R� �]!�'Dz�9�C͕ NK�.�>o�!��	X�y�T���$l�7-�6.�!�dK�V�^ࡢ�O t�~��W��1c���Q2%����G*� 	�y�ƍ�K�\h!��Q��`)��y2ɐ�a[4aR6J��F�vQ�����y�$]�vu��1Oq��j�5�y�E��9���c΀�Ha��⓭̲�y��~�4-�K;O��T��y�X�dfDyh��+�R�+$��y�)X�T���H� �+�
�yRaTv���n�a����oܱ�yRV4�2�Z7	�V��%*�yB.ѝC*�;��ǊK�hA D@I8�y�Ő�..��
)q������\��y
� ��3�ˁ',�|��T�6��3R"O:�20���)��H�#��/�
�"O�;��>.0,Д
�D`r�QP"O$	)��,0r��
l��(G"O��Rq�Yte�e��!Zv��Zs"Ov����F>Ґ� ��Y���1"OB�Y��M�?�2�;B(G;|�ȥˑ"Ot���n�Y�T[���L���5"O�١�� �*�U&"+�vh!#"O���fQ!�%Ҏ:��ܺ�"O �z���;X\^U
c�T�d����"O��zq�!��U���M!p�*y#�"O^�[�� vv ��l�b "O"��VKC�_�Dp�2�K�Y�}:�"O���G!CF*``&lN�&6�� "O<��mBi���딵 ���v"O44)C�w��9s�0���C"ON�AP-A0{^�8�S��xMA�"O(1a %��l�Y`-���D$b"O�p�%o:��Qe̝�n�%qd"O��� �6y&\Y�1��#��4"ORA+�!9�୍�Kj���"O��R�&O0מ`�u��!Q�F�@�"O�q�b��dx�PBʨ)��Ht"O��k�	E�8�<�B���9wԆY�"Ob\R��Pl� 5%��^)�"O����":,xH����5f���"Oz��f�Z�~���&��j�b2"O�P�"��t���@��U�I���"O�	�ĆWdI[Ч�	`1tX�"O:5���J64���E-|�
�"Oj`Ñ�ٛO�~m��E8���	�"O2��Ȕ)��i;�jJ�{��2�"O���"CB	"�U���_M�¸ s"O2 
���TM��p�_<)�H�&"O��A��wla����>�@dc�"O��¤,J9{�Ta /N�mn�e"O�E;V��R�,-ђ��eHL�ڣ"O��b���AK���N˨6.�a"O �z���i�t�W-�}��l�	�'0��j 
'"I�0��k�D�V1 	�'PR1O<I.�۷�������'��؋ÃC�y���C����$��'by[��� ��y"���8�2�'H~}�r�>z�����'V!x��'fl��}/����J�G��p�'�Z��dF�c����!K�;�L��'�ƹ���ڟ?}H�"�9Lp��Clli22E�#�Y�����*(�9�ȓ<@H���;#<����@=k~�U�ȓ<z`ј4@"���4�Q5Bb��ȓ4�������7~�&�ᆢM*?��هȓ	�Z)���$H�Ѫ�z�4��q:�-��aH�h"��b���-Ņ�K��1��N�F�{����p��qɦ��Ug�?`�]v.р��Ԇ�Lr��q%O��IZ��G&ZO�цȓO�F+�/E��¢%D� ���ȓ~Z
(%`�:ak(!��#[SX⑆�5�`qp�++ʹ��j�	�:��~v<�"���j�t��!C�X���ȓL�鲖-�-d� �va������'�.��6S�5
Mi�^�`����ȓ1b�EJ�'JX����P�|��S�? �I�q��0XX�QE5lL���"OX+��ւ0�Q�BʱpiL�""O��e�O�8�|��N�{��A�"O�	�p%�
�b@��o��`-.� �"O4aZ��A0L���mF-_ ={"O�H���5��"��%��uh�"O��Q![�b�ܰ�UJY)b|�9�W"O���&����p0�IY(5mX�"O�=��+��TX萦�Vtcj��"O:1�f�-��Y(�'a��z�"O�,�aN/r�H!��ՙb�B �"O�lpvjE� `��pq́�|<:l��"Op���ِ[7��i��4e��q"O8���L�7Ϙ���mJ(<�^�ҥ"Of�y� �4��,hcmW�<���"O�����U�^$b��ј /nt�1"O ����T@�PY�F֛m�<��"O4��)��>U3��C����iD"O�%{훏=J�����d�s"O��@��(OB!�G&ȚH�B�"O�Y۴�A���t'Q�~�Ȓ�"OB�i�nR5v�"da�*/��諒"OZD�%X���@��d�p���"O�ȸrm��9?� ����3"|l��G"O�ȉ�ňu��Ԭ�1�"Oj0�A��0oS�A��A|�4*�"O�����)�
#FL�.�.�S"O�d���?�jq��Ŋ�M��tK�"O��	#N�o��a&5yb�R�"O<��/�jlag>)x�Y�"O��gm�t�0&\�J�F��"O��J4��X�"4�$��t��!#�"O,̻Q	;TRL$G>`ؼ��D"O�m�U�ԓ��5
�Ě�?r.�!"O���6��lԮ�+�$?��"OB}���Q�mm.|q6F�C��9A"O|��d��{٘�C��R�R�Z%B�"O�d۴A^�K�q"G� �r|�"Om��6���"������8�"O�%�G�9"�^��W-��N���B�"O�р��O��0�T�T��"O~l#����$�j� �P gςD��"OT�0�(E�r%z�Ȱ,�/Q��{�"O>����PT�ʤ��"F|��"O8d"�bJ�h�*�V$R#�$
"O���0�. �4�#d%�38����r"O�<��A;���:"̙`��Y"OBȑ0`�7/����d���)�"OB�C#N�^���֧S�4Ő�"Oh���
�ۊ(0��w���"O~�Q"$4~TY�Q�]�� :�"O�l����?L�ģfM�f�~��"O�Y�L�=5'h|0�,ճ4VH�T"Oj,)��_�@�h!�U��7>���"O���@}:�P��R4��9�"O�}Q�\3-��}C���S�E�$"Ol�H�VFLp��Κ+
�#"OZ1j�%��qXX�0ЏN�l� �"O�x ��I�"ۆOL܈�5"O( ��	ӷ!���� �O*��Q��"O&�pW�H�w�C��k��RC"O�$�V	^��,�q'X7Β�9�"OT��`����Ԓ����x�6E"O�p��i�hÀl�$��$/@P$s"O� (K�äy	�%��W�`:l�I�"O2�SԮɉ*�X�X@`�.9�<�"O�T�B�B^���1勨[*�IpT"O,ȥ�@�JZYB�uh 1R"O�EiTH�3c4��aaB#M�%�`"O��;��/C��,��j�08J�`1U"O�tJ�흠|�j��Ɇ=�Qʰ"O�YCgȤl�|	P�MRB��@�"O<�@U�����O�T��U"ONTD(��f�`pB��P�I��*b"OA��*�O
1�+I	�D"�"Oz��p�Ӧx�R8���T*\���"O��O��1����Ôx:��"O����-Oz�`�fb�!9v4c�"OȄ;&/�h�F��"쁍{ �y�"O�+�ȉY�\`rT�3\X���"O��'��?	�!1aBP�0��<:&"O������a���BG�[��I�"O6)s׀/<@��b��|�~@��"O~�4o�<��"@�o����"O�L��W�q&�\..��%��"O
�+��ո/g$K,��V���"O�у��
�P�ؐ3���NuH%"O~��0#�0�(l@��Z@p�,��"OrL�N�Ao 0��g͊D��R"O`�	F�&(� t�D;��@b�"O|EIR�O!/�(Q�p�Ȩ�y�F"O�U�&%O� ՌE�'C!�=1�"OH�2U�]�u�2�	�Ş��D��"O����X�4�l���$�& �"O�	�2i@�Vqf����6�@ih�"O`L�v@�8����*\@�S�"O�!f�I�"tKߩ\�� 4"Onl�ˎ�^��j�'Bd1�"O�=��K]`ae�1(-��"O�D����+)����cĦi�P�rD"O.!	���`��Qb0 ن����"O@�1��&!XeB�� ��Aq�"OV49�;��Q� Ba�}�f"OP-)�L��N�F�E��AD����"Oޅ	��D�o�T̹�f�@����"O���A�4c��hj���?n�X�"O�)c��:A�x[��M�W$l�"O�e�X��L��#2*m`�"Oh�Bq��1iKʰ`R�#qU��"T"OX��L�j�ʔ�t�\�PT��S5"O����+U?�vd�T���c��J�"O�4��?W��2�mݮy7��j "O�)A$�&),.hra�G&�(M��"OFTZ��(NSx�a�����JQ"Oڥ��j
z�|���E�U����Q"O�P�(~�[�V�m�:I�"O��%���
` �A�kd�1��"OfajĤB�~��Q������[g"O�p�b��b��X'h�c�.��f"O�16�W(3q���a�n%\9b�"O:\A�.ɹkPޑ��A &,r"}bd"O�Th0&�V�h� �'1`z��"O�� �� ��pBs��W��U�6"O�-����=F��n��fʸ�$"O�$�歋/R��ؓC�~��B"O�`g�&��y!��/8n���"O>��R��+���X#�VY|��"O2���"�7��)�6��65l%1�"O� ��"���1��a`#�5Mvd��"O��и����p�A.%����"Ob�a�d�R�պeL�*�5�0"O�`�Qlˠ&��ps�X�����"OrTk$���=����f��[�D2��۟��&Ҭ_s����r,�Űw�W�nQ��S�!��?�]�P2H>����I�6@��iS�U$#���XE�=���Q��(h.d �!잙V�8�QFS��II�7@�{S/Q��*\c���e�'M*iI���?I�����i�����紴{��	R\�����O��Op�d9������m�yI�!SgFiu�d�C;�O��m�ԟ�n� Z�hd$D=�y�jM6xۼ �V�i��tbc��ĸ<y,����Ob7-
"s�h�OO="���&�(\�丰a:E�ph��OD�'��<�aDׂ3�`D�"K {�"(H��Ϧ�������IT7Llq���3�H�kl��x���:�\`�E/ :ݛ6/��?a�����'�?7�@8{�H�E 1V�Tٱ�â@����O���(�S��(T�J��~B�\Y�$X)Z�<Y�id�6m)�SϺ+��:oM
1j ��84����L��I�s2��ڴ�?����?IO>��o���`�)��k�,����Qc�����۠�5#�O�1PUke=p+MD=x<�@v}��O�o����2��xb�7'Q����"�ype�`�Ԁg6��>/D���OXx���	���'�����ڗ�~!'щ]��y�5n*$� 0ףԠ|8�`�Y/#��� oӄ7-�Ǧ]�<��?ݕ'�,-sr�F),k�iæ�u⎍c��U�����'m"�'ɧ�4�'zE�.O@��)��n׌�*��dc� ���'�� �ir\��;��C�~���I����t�ju���p�����.\��i��(0��P�z��E�S�>�⑁�N��@��h�S���գ,�>�����%bۄB^��~�A%�S�O|�An�W��y���N35���(�'�x6_צ�'�J�K�f����.�)� w�h�3z���We�33���?��o5ԙ���ʊ6Z�I��x�O����D��w^�Ԛ� ͟�JT����H�N�d`Z�.Գ*yj��U��ŀ �J���Ϋhj@���HO�����'A��u�B�$�~�AA&<�����/	4�Dए5n"�4�|"=��MI�(���/p�<,���s8��Xش.���i;��A�[�����敺z���'���ĩ>q(O���<����e� `�4+������T��z�iT�Q�"�x��'��	>Tv9�!&Xk�61�@$P=�7�F�PW0��Q�U>?x�)��̄�H-.��%��r���¤�}Ӏ�P!�'�op�2�$=���2WWM�tE��'�
j�V��T������Oy�'��	�M��4�f)�7�X�Wh�����{Ӝ�,���6M��"��+���7���׊�N��&�ȅ퉂w�� p   �   �  �  �    B$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�U曞@�VM�P������@��P_`���'4r�'d�|J?��f�s^hy�&A�x������ b�8�`XTv�|2���,�
�*��ڹz7"a��iRȖ:[�Fi��	�[ڀ3�F�\l����S�
��0ɂ��O��d�O:�d�<�����'��ر`�W�z�n���iЩ7�� 
�'�jpQ�,��t�U꛵{|l��{"#e�n���<A�b /�?�����fJ�,���Y*�ڥ�EHO� $����?Y�U'�l��'z()��-���B���H�;`k<5	�h�){��?���>���ň;ByF�Bꈥoay2,���?������v�\��3��~e��ɓ���0����Ol��-�)�S�?q��/ۓ���C4/�d�C�	=`�Й�B�_�t��	:pF�~E��`2�韜�?ɢj�@�Ͽ#�7p��q�NP�J��Q��6R��'�a}b͟QI�`�׎B�Z�*l�f
߷�y�'��Ul��[����}�@U���y�B�f��yz$��:}�j��ej�%�y2"ǟѾd�#�-,�@q��@���p<e�	<}�� ����`?�tza�DU�:���O\��O���'��I��4�C��Ū3t�( *M#��b��+ �$,Of0��&���*T�U5�\(D�$�mbay��Ⱥ� +��Z3?�&�ա�'�����O���RP���Y��I��fV�$K�(�p"SO���#��&$��	�͞6&n�p�,($Ec��(}�&��|�����$��::�i�V�%C���e�Ԋ!�lK��O4�$�O��d9��~r"&F�L����� �45`� ��A%h�d��o�&=���1���Gl]/.i�)����Z<)�j��c]>�ň>,Fĕ2��	^vx�IX؟ �`d�Y�P�{ � T�>�@� D�(1! " ��Eɵk��<�s�j �M{��$�~��A�(���4 ��7�*��2��y>���=���O>˓ I��"��ߣo��u�)9?Ԡ��F��r����y � ыU6��ȓ~�p�k%��^��1� �
$F��ȓN�� ��啦 jN=H�Aއl�І������(����� #zy�q��K!�2�"MF�����X���KV�w<�%2�M_�I��$�OD���B<�����J��`9���)�!���r�¹�P�D*/���2!�ah!���#S_l$�f��dQ�ݒ��߂*L!��F
�L w	�zE���'�@�H�x��#���P�P��Sap��M:L-���J`eEx�O`��'=�)� (仃'یBx��"���6�˰"O�q@�	��@�aKb�1h�Lm�"OaP����`��\���3��"O���lr��-�3|�z)�u"O��vJS�-��H+A��usp	A��>i��)��1j�L�B��ΥjՈ��1��+���'*T��d�'7B�|J~�A��99�p��G�fp�3�C
Q�<Y@��d�f�B;R�&D�S"ML�<�#ۼ|����#��(���H�<)�MםB���5
�=bxD����G�<1�Ç�;i��aڡb`�Ց��^ܓO���u(�O�=�S¤�BHC�e �s�۟�&��)�gy"lG",*Ȼfc�7hs����)���y�Q^�H��0��#�$��y��O��z�1�
��} ���qAϬ�y(RC��U�?A���I2F��Pxb�)�Ql��\�pH�Ĩґ+��F}Ҁ�:�h��=a0�A>�R��g�*� �ȝӟp�	lX����O�N����ql �Y�b@��;D��SvA�zb2��Kߺ�
T��=D� 9`�_�#X=R�H�8����'j8D�8���_���K��X�Y�(�RT�5O�DyR�G:nJ9XC�+����W�L��~2'��O�)�Oj���>i#�\��:�b��Ǒ8���k6`�V�<�fM�iH��&k�T5P�Gi�<y��
i���uA�&/<�� �Qy�<)��8
;�9$N�Y½�eQZ�<�O�3��2&
�ڵ��QP���k���O$�9j`&15ʱp%a�m����I�h��������v�)�i	0�
�ː���3^�M��LGk+!��;m&yBQ͓�`���k��H!�d�,PD
���/�|��Aɂv%!�$
ZO�9eD�J�΍�s
B�!�$PGS.]*��;��xH�jqO��D~2o�:�?)�O	�s�  ��ڙpmr���[��R�|�����I8)a�<�7.G3@O�t[�/�Y�C�P�2��¨-��X�΅=g�B�I�x��u��
�&%^��#�
�T�vB��*H��!(9�`"E�^�hB�ɛ0��!�@��� h�BD�H2�Q�'7�-A���L"<�X�a!���C���&3���I֟P����#��� ���9�h��(�+T�B�I�-m^��qJ\�{戔s�/	�ZB�ɸT]&� �Q��\�Ї��LUXB䉌v�>���Ã6Lh8��l�p�J��D�q�'���c��ƙ��%P!�ۢ��(q�'�0�K��4�����O��[�$%h����$u��	��[�$`���&�A� � Gt�$5.]�t?F�ȓ|�@9�e�-Dy���L$A�bф�b+����`�����lr�ȓp��$0�&��i�w�>�ܴ�O� Dz��4&ɖyy�p����>'˸@
�����	��š�O��$+����m�����.��"��b�L�yRD-k:i�4O�.0E(%l��y��X���놆�
}\yQD'˒�y�g�m}�p䃏�z.*)�����y���==u��AK&q��ih GȊ��'*�#?�E����ܓ�L�hFa��]8��!�=�?AL>)�S���'(���Z#��hi,���f��MG!�	:��ѡp�Ĵ3&|���R*!�$D(7�习���@Jm:�A�Vv!�d��>�p�$ =J��9���+#�𤜠
�\+%�3y��D�G���m?\����
=��>q���^ j�`�v�Z{ج)!���?q��>� �8�G�?��L[�"�)b��""O,����s�����E�<��"O���QfFI�Ѝ��:{*�Z"O|��ä:/pCs��~����'B�<�ޯW5� S���2.�H3L�{?Q��Fe�����'N2]��`d\M�֨H�@�!qg����:D�(�GزV����j�+��E� �#D������;%���s�f�$.A�\I®!D�TK�b�+0���딡!v(I"�>D���hB��(��EƬ8�<�!u� }"�4�S��L�����J�/vJY[3D͜<�q�OiIAI�O���3������8���Y��Y� ��������y��E���[�G��jP��!Ð��y"/��x�P)X�e�H�R!�Q�yJ^��qႨ��a �1бnD,�yBeܜyd�� ��*� ��@�C��'�*#?� �Ꟑ�g�J
�pt�2��4�>l�V��?!H>��S���DX�^�XCB�Q,�$2S�]�,�!��.�B��#$Z:a�*�w���W!�d��~�U
Cd�=H��e���v�!�DM�(������E,<�Vy�Cm�F��ā+M����G^
xL"6%".��$�>����X�s�, �W�W�}��5[����?9���>I��� ��p�j�.c~��R�cGS�<��C<o�y ��w`R�+�J�<.�Qھ�Jć!�b!�*E�<�2 �gm~�`Fĝ`��;#d�\8�H����-�L�ە��> �ݡ�m�F���I����\��Y}��Y�5�آ����9��9{����yH��E(
%Q����4-�Ա��yB���J�`��)�$4RJI	����yB�[�g�X2'm&t�H8�hO;�y2�6Rzp��Ag�@بCoA:��I��HO�$�zwΚ�����$}}�=��>��֑�?y���S��q��yC��1S��Vi��C�	�N�NhT�X9T30��Q�ˣ8�bC�ɆP�ɩ�X�"`n�(�+�%tB�I���B�aҀ`
t��E�I�"B�et@�@#� ����G�U��X���<I�� cNxԙ�	J���:U�C�4���%���O>���M1��%?|8�a4�������E����s�Iy�G5�&m��[�>1�5C�D�Xu�QF�"��ȓJ8���J}R8�3D˺%����~��m�5L[�\��`6���҂�#�#<J8G���
,�(���:F�x��Rɨ�$�O0��:r=��@�շ9��Q{�M�@�!��]1 ���q�+�9`E>컕k�NK!�Ev�iP&�%Բu�a@Gb,!�_�vpi�CV=��1�i�-%��xR1� ��M�pk��<M24⃋��\�X��$�"Fx�OL��'���9L�r�&��v84��H��$�C��$q��
Ѩ�9#fԨ�j@>1C��"h��E��/לA�����%J+�B�	Lb9�ÆȀ	#8t�V"�x��C�	�q�z0�e��#�|5oZ!P��'�"=�z����2cj�Ј7�ʕ�F$�R������OH��-��	V,MQb�ɍ�3�24A��5�y��٤#�4��#w�H�jA�Ҕ�yB%A`�V%�q�Зo*���
��yb*K$���΋�R����m���yr�B���\C��#K��$C5����'�l"?�rʟ�˳��8D~�� E�MF8��O��?	K>��S��򤗗g��AB�˾`{"(��Iս3�!��  1��e@u��8���H���@"OԌ�e�^�2��KE���+����"O�Q2+_�F	f� �H�#�ܤJ�
OV�k�3+��2@@��8��e�����O��H��S+�~ ���ͼHqh��v��!+Fȵ����?	�	<t!�̇�: �A ���E�4��ȓF��dՋİt���Õ���q�����$���7(ܣ�����'�
@����+O�UQ�*�Qo���r܎- � ��I�(OD)Q�*�)>��y�5�Y>}~����O�rb�i>}�I���'\���צ�1�P��-P}R���''�e�T�;n�z��Oչcb���'c����f>w�j	����X3�1�'x�`�􇎋@.��%�8f�t	�''4� �=/z�B�.�3W�>�N�h����)&U
n(z��N<3A��IK����|�����?AL>%?��S�T��bP��N��@���?D�$�f���T�b9ص́�?U4Aa��>D�hơ��b���'#˷Q��v>D�V٘ ��) E�s���	�Z��y��Y��r㨚(g/ tȱH���'��#?�0G�ן��$DٚR+��3�Y�&��D��?�M>��S���=4.� �偙�s�0%�r�X�E�!��<A��#wA�9��h3��be!�S�c�%�%Y�v� ԩؓG-!�d.]T��4�hr�`M$���Ȼ.������-7VP�1�D�_���䑞u��>	sg-��"�u�2��!���7똰�?)����>qV��
&�(l'��#iv�r�jc�<��aA S5Z�颥�\�>��q�_�<�aP� �n@�6��$����K[�<�C�x=\H�&�P��0jN{8����dF�q��)�7G�b*����L�/����n���ϟ(�IC}-'hpZ�
(!�[*C����yBg�0�,A��R8&�H����$�y2�Еf��͛���+"P>%�!�\��y2��:�ɥ��lr�@p�ۥ�y��Y�"�����m�+Ro�� ��3��	?�HO�2��4�S:\�ҁ�&$s�4:1�>�0�ϵ�?i����S��/�ё��~\ޠp��Rw��B䉝2�8d[0΄ifzR��bM�B�	�p��a���)C�j���k�Am�C�2i��5mޡoX�Q�gŏfKdB�	4%�]H&/��IDT( !D�hJ���r���E-/��8{���#vî*T�ç!ͤj1��d>��O>�|��������pL�Vc�=�y�ȓbTȁ��N����q���T�O��#*`88soK�F-|��g�1m�,�ȓ��e.؍\�nMb!B+=L�a�rt�G���;jd�!�V��e:�=��r�D�Td�]�8<	VX+8�*\��j�/XE4���O������t}�DÐ�:z��!���M�!�$D�g�����?q�8;�-g�!�d�U��i[ �F&�ƌ"�m߬b�!��ں�Kg\;� �6Ώz��x��"ʓ{j�P�S��)��a�D�5W���E��Fx�O�B�'��Ɉ8�
B0���!�dJ��g�JC�ɪ�AH��ep���GKǋG�.C�<7<D���>�Ȱ�7!B.Y��B�	�i*���M�Rf����şz��B�	RYРs��P�P�wiɸ ���'�^#=��얶g��m9T�X�	�.��@cQ�D�7� ���O��O�OW�s$��)b�����?&��'G�P�&�"���a��,A���3��� �]ytG[�7���V��To�i�v"O4P�P!M{�h`���h_���F"O6I��*�<6���냁�E^z�`��d]�'�fX"��V���R��T�l�%���Jb�vje�'��'���Y����,J�,�@���ܖ.X����*D�� �mδ��S�Z�65�'D�@c�b�*դ�%��Mʬ*p�#D�|���A�,s�$Zu��k�֙�'�+������v���IcN:9�T��m�3XQ�$�@F0ڧH��Y�)Z�Xl���J�J���'���'�~���$j��`9�c��z�0	�'aRX��e��$��Hi��F-Y��1R�'y�Y���%}�DI U�?_h|P	�'�f�
&��F.�]9T�P�Z6�9�
�Q�Q�{��s�u���"i2re&�i�'m�Y��h���O��V\�ؐ���%R�t�>o^c4c�-~(�k��OpTR��j�g≽[т�H��F�w�� ��@��Y�v+�6.�`j�'R&�A��4�3�$�_ Y�%F8�$)Zi\�|��	y~�jҸ�?ͧ�HOL0D*�a���8bH��Ft�4"O��vH��29�g&�\2����>���i>���_}b��h`�hrV@O �zH�m^�I���
������䟀'��O�\�("mV�{�DՒ��ז2��r�N����4OP�{[��X��'�d-P��ҽWh�a��s�h��Eʟa��]��8�J$�'��	��i��?ҙz&��
L�2�m���?	��hO�c��(6�l<�|��a[9��Bi9D��4 X;��sE\���Q��`9�	��M����'k�����-`d��BW��Dӧ�V4=���'1�'��Y��!�{Q@�Y�'�<l{BJ:D�h����355�����	WB([% ,D�(B���i*lAT����iiG�/D�������L�Y��T�&3ȕ���.�� rFD=�<���`��C��1���LdQ�(��#<ڧ%�M ���]�Dmz� ���1)A�'o��'�ڕ�P�H
�x4�n�@Й
�'P���j.X�F�B
�{�@���'�b�Z�m�O��m;�I��/����'�����t���� 8�(�Ǔ_Q�D ��!\<��d�m`���Sͮ���)��|����?y�O ���h�-eڴ����L�1&"O0��Ӥ� {v�q��øq)e(�"O� �2͛1���րQ�(�4x�"O@����$GM�[��[/u�|��"Ox��e߭lh�QP.G��p("U�>QT�)�S ��M�*�h�´���=����wb/}r���z��'ɧ�'>/�J� �7=~th�O*�,��zLi��L�j�x`�u�P3�D�ȓ�0��1eӘiA���g�?�\��_��*���K�����+r>1��M�BuҦ�"R<f��clм"6܍�=���I����$�<C�!�JE}��J��"VzBL�Id�I�"|�'���vDL@�pPq���Z���K�'|X�顬�.JM�)���E�R-����'��H�B�	 P*�B�K	�BY4��	�'FŃp��3L��m�$�B�:��
�'\@@��ӻ+6�Q	A�ۡI�0�q�{�'W��9�'_�2�����7$zj�)�K>pQ ��5�'��'ߠ��2*(���lY!zc�0
�'�\k�ǖ�pL:L����wt2MB	�'R�7�Ļ5iʠ �l��}8@��'��X�_9�T�ʡ�F�!���ǓQ� ���V�����(D'�p|Ȣ�3D�����  �    �  �  *  y  �"  �(  P*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms��a?Aab��jD�O�,P���$�0y�x�����A��j�w��}�n�W�R��&R~��YBd�*���$� y�~`#_|X, ��o��L�#hZ�i$��`N:�`�O��t��XF{b� �v5��-��.s��c"ճ�~�Ƹ�R��!dH���J���7�ybf�9b��a��Ƿ��P�F&�?!D�V��|�¬�,�`sgb�i?�"�%̓@_����duP2��%�y��K%i�i�J�PLQ�ALR�>T�D��f?i�f��."�O=b@�V�DS ?G������_�h�n��0?I��Iڂ�8�L=*���ؑ�]�s�z�*5�X�L!LԢ@K��=)\9��_��0=�F�]�"�vT�YI��I!G�&\5ўԡD�U���T��*]�QHh������]�p�hQYB�G"{UlՊ7�#D��ٴ
L�K䱱"�D �2-94J�O@��@Bδ �)ۂc�T�ض�O���`ӣƠP��/0�jD��L-D�ȹĬ��s��+�G�����-��k�ڈ;��O���b�/O���'^�~(�<A'IL<{.�Y$�j��ط@Hvx��ٵD@&T�D�2��A�!,V9H��Fe�r�G���D�f��$� �`V"�q���S�˓I4�yb����l�V�Ha� �"�TA��`M���#c)��5{��!�L�����ȁ�g���ȓ�rP�5�ڛEC��!dO�	&���	%}(�X6 @b��a��Y�;���)��40V�e
�Rw|��&�C������4�|���62�V�h�����8@q�'`���I.�5��é|�D�ۺ��'�J�(���j���ɕ	��s:}@�S^�}Aw�ܟ2ܠ���� 9�
7n4N?���		P�8	����P�v@��l��VCY�-��Q��[n E{ @@6�QTbóX�4� �Ɇ�~2�J,")��"@a�"� IZ!L�-�y�	]5'�ҝ@��(�Ҽ��"���?q�(�$^����*Ż(l(��Ue?�r�K�}`k1��Pd(��f#��y��{�ir4�
hjR\���=���5
�v?Q���f��O��@Q�$��@��r&�d�f�#���1�}"���$q�Ț� �����G)~��%*������H�_HΌq���(z�bi�C�'��4" ��k��)�(����EI��$��͈Ȳ�Œ8'%
%K2#4U���0k2�� ���������O�]f!� �a|���W�;M،i[��IW�#�^% �҆ɐ��J��v���~���IXFr�8�Q�)?
@��l�E\!�dٛ'i�*�KCRi:���ͶZa�x��S��~��f(6�)��ii@.%�I�{8�ԏL�$�����2)B��"!i�d�����Ed��°��Y��1�0�+T
�YFB�=,�~����)�n����3�Б���I3j��rd�6ў,��*T$n�hЈ�!]� �6����ȓ$�Z��� bBE�&��d���$D��7=:N�X��M3��J�i�	��̞^4�2P��6�´���S�'QƀRp��;R���P'F)H�.!��'��4���R01�g� xt|�8�*G��x�#����o�Y��gQ1O�٪D��:R\��f�/V��4�""O�b�@�TY6�G/\�]� ��"O:P��F��'j1���20���"OR��!�CY:��-ƆO}�<`V"O�����+]�Yr�͝�]�5;`"O��C��,���R!�*v4�@"O���e����4���|V�\ۤ"O�P�#/I.��zU�y@�M�G"O��iҎef`�b��z�41ia"OL�P��
eڰ�B��>h�Hȡ"O<����&�&,�Co��`�����"O�aQ�ٮAf���ݞA�a��"Opy����L#��1BM�4%�U#"O�,�l�>p���$/^IwbA�c"O��؅��&Q�H�aM�>?�dr"O,aYgi'A-��BR�:=���Qg"O�����gH���S"ۼ#�H�5"O��@�#S��I�D�23��_�<�MG�:�m ��/x`�hq��W�<��hڜ&�|�3����"@p�"V�<!�o�?l��aV`��a�j�ծ�Q�<�uG�\W ��𩛔mY�iNTQ�<��l k�8u���֐<��%y�e�c�<A��DIU���'�s
ԡ#$JX�<���<�
�H�I�X��a��o�<��\�-7�!���>Uɀy��C�<�ŊҞ10h��> ��Z�j]�<'�H��z}�Ì%�� t�M�<Qe�9��@`r��5<xt؆"CH�<�QW9<ī�-�n)�Īs��\�<)r�Q��,K�� +���
3E�V�<1s�=f\�zu�7�Ig��m�<�uF/��|�4k�+22n�t�b�<�pbV�D���I�Dg��|;A�a�<�W��3��s�	�t��}ZG��h�<q��ƌ65.x���k��5r��K�<)s�
	�j���zP`C�<��h !�4Kfj,i5��ˡ�@_�<��;yFy�dϩ�l����S�<YÈPV%Y�@ͼg~9��OS�<�5BZ/Bf��{��Գq#�!���CQ�<I�i��9�X= �)B�z@0��Y�<p/D�'"ȍ'�%��cU�<�4��#m8d���K�jn:<{�I�<ɧ�
T	|}Х(īL��0�A�D�<Y�j9�p��q!��ܹ8R��h�<�q�W
��:��$^�ʙ�EF�a�<��e�,gV�l�����\XȔ��B�<1��ڦ"�䛱�ײ��=�Z��ȓ<��(�Ǧ��*<��.)a��E�ȓ-
�CF ѳ5a�c�Ο?q�����S�? ��@BC��B�a��c��h�"X�"O�a����4�@K�B���}��"O8�ā^!Of>p�3�C t 9Hp"O��G*B�zD�4!��$BY��"Op��A #+:�� ���$._�D�"O�9����8�Q�M�DE��j�'��*H�9�4�fEE�_�6P��'U��8D!WQ�\HQ�^nU+�'���1`��	h,㰭�Y��Ls	�'����͂�mϲd@@$C�V��r�'8��ʃ�ޒ;e���$�EO�>��'Q�H&d��b{�0�T�p˄�	�'s�PC�-!Nv�h���}�Y	�'��};'�@؅ic慭t�� ��'���s#�G���k�c,i��0��'�Nx�" O69J|��iׯn�^�K�'�l�z4�R�2L��` BH�pN0�'!:̩s ߷r
��3@�"|ծ|p�'Gmh��6�^�B#�x*�x�'�+o�61h (%�.!�U�V�/D�` f��L��0��8T�Y  N:D���� ԛH9��{� ݔ�����&D���M�mJP8�癢k���R��%D�t�%!Y�,@�i�v�X�9ž�Zc#D��V��Q0����o��P2�<k�d D�� S�@G�����Ֆ.^yȆM.D��A+�9Æ8��F$�>��`�&D���5̏�u[̑�Fj&2[4A$D�D'���+J��p��#g�2�1!-8D��+A�יఽ�T��_�m`�1D�|�t�;;8.<KAM��ۅ1D��p�B��JΊ���",)�<�e4D�|�*V�Ghn	�R� V�t|��(D�h�T�\��8R$����K�f5D�x*HѰp�u�@�b���W` D�j#���>p�C�D�|8���"D��� �I�q�M��Gn"<q��!D�4b�)ރ�f!���P2���j@m/D�4�P�Y�Q"P�2�O�!?,,��7D�t�J�!>T^+V��5T`�i�6D�<É�/�nhhuD�#B"��F�2D���I>���S3IC�	��4J��5D�<+��1i&�ɡ&l �L���E3D�tᦨ	{�``2
ϯ`?|�!"�1D��xR�^�����O���"s�?D���!!��m$�I�ɉn��B6�!D�`('�M�N��p#d����M�W�,T�pr�*�@����2hֺuؕ"OVaʰ��t�`��p
��=`"O(��LP$aVV�q��<]��"O�aJU�[�?�=��L֋xYv�bR"O����*,�,@��V�
_J��"O�x��k�X���"�l�n�Hq"O����+��"��vȶ�Pq"O���O�%��ՑD74�|9�"O0���x/)��O�2���J"O��c�m�ϢAc �H7'�2� "Or�y�̘�{NѨe&םUBB�k�"O|�
��%0�2� %	&@ȑ�"O���𩇡 G.<�&���t�"Oq@�I�l�\ �B��r���#"O�<�7�ɞm/ؘ�oƱP�%x"OH)H���@�Ne9.��sz����"OĔ� �ק�r�{�NS�Fx��&"O� �X��N�C�j��5��vq>��P"O��a]�- ��kN
*prmi5"O��f�/�X�	���2F�u:�"O�Ih��B<&�
��6`<ƒ�k�"O �r�Ā(�5��-T�G&��W"Oz0���ә/"l�L 3�Ģ"O�8v�s�NԺ��:����"O�A�&^�81h��t�ڏ��$�A"O�A��dY������GͰTy.�֎{���/B_X��J��!h�؀i�̋ ;���@�=D���I��xz$��:p����<D�HL��X����ؘ��=D�4�hC/VD�(��׾�\����1D���c�*����
	�N�[�,1D�p�T�N���l�e���Z�,,�e`2D��@�J�q��(`!+�z�<�&�1D��P��w��XD�.��0��*D�H�
��q -H%��I��;��)D���g� �?ab�i@E�S��}I�,(D�L��	�_��9�6#
��:D��)��˱H�Hd���D�RJ�S�'7D�S��=6Y���E>aT��'F!D�x"��ѐ�j�zjN�M�X��� D�3��A�z�$��%@�8���+0�1D����ջ:ڢ�B��wv�]�� 2D���	g	Ƒ�wj�1�#%%D���b`F�gyn$�fǋ�q�~	��I8D���T?���4(=�����8D�1�%U�{o���*�C�f�X"D�<�%2BW��"M ���K"D���eN�']*mBC�ðSx&��!�"D�<��X=Lu�d�򩀼-�"x �@!D�T��Hߺ�HT蜔W{4dB3+$D�����={�Y�"�P����!D� �r�¤��K&g�q4�a;SO#D�0�2�^����ĭX����ej%D�t�c�F�<*4�&�@��׉!�$��(>l�2�T�<[bI�.�!�ć(hЄj�-�t �S�!���[��y U���`��M�@!!��!#Lv�P�ǒ���D�c!�Č�J|8��_7����:{�!�䈸�h��򎊴 ?8\�[>�!�]+�:1"Q�I|%��*�+\1!��M�U��JE}	h;Eܭn!�Đ��x���~�B��E�Q!�$�_u>9��A'�H �&��!�DL�,Hi��f
�~ɨ��U��!�d]�����N	~ D ��%v!���������3^�L�Bp�	d!��-�}�ģƪR	��Y�J*D!��ҺsY�H:�'�
S�@��e�,V�!򤎿b��� B)C-�QY�D^%N�!�d��GG�p6�ͷ>�!�5^6wy!�M�-P�G�0k���4D�c!�D:/t�Ȱ�)�]�@U�c��S�!�	'�T���Ȱf��DI����#�!���}�$�2�"�t�`̹��1	l!�Ǜ.������ծC*�j$�\j!�#�$���n�q�*�qFe!�!�ēq�"���'��v�L,_�!�ǣy�$A��DK�X���fd�6�!�D��5h�q9�LY9i�m���Z�mN!򤐖q(�����c��	
"S2!�� ��YC%N�o�Ha$�_��-Z�"O
m�ǩr����cA,lF$�V"Ou� ��T�
��ͼB+�Q��"O8S�a�HoFMA'FF�$�<��"Ol<!��[4H� �g�'|g�|�G"O��qA�hS8g r@E��"O�`��F`��81����:;�M�e"O�y2kӜ%y�,�����u�S�y�L��0!v��-�,�xt�K(�y2�F$E��qeO%#�m��,S�yr'�)dH1���I�$�h�� �y�ĝ�*9�y���mn�Kw�Z �y�n�
s~Cbd�"j|X:N��y~"����
^t�=j���"�y�"\�������[�h��˻�yb�L�k<ܤ)��N!U�H�f��0�y"DՍ>�D���Z�i��4��N��y��*ֲ�r�j�b���� ���yR��0�p���m\7G�t��)	��y����44����ד��X��mP5�y"�R�
�ڡhӄ	z�24s���y�oY8NJ�aǠQ�_N��j�7�yB�˭7~)�Ώ
w(�����y�K�ml�@��L�Jxu���y2DT�%v�!����i+.�y2��>��Â��z�����H��ye	/l�t�D(F%$)��ē��y�,�aH5(4eJ"xp!Cgπ/�y�)�Vvx�n���8�q�[e�<YaD]!5�СG��eQ[��z�<)ƍ_$1x�]%�PL����Hs�<��`�*��Bg@?Y�S��g�<A���cĸa���)z�J�de�<Y�*��26D��N-5�P1F�Yf�<I����Vd�Q,C7����&l�<��͊X�@�q�P�;�,sÉFk�<����C�t�2䞅~�)K⢛�<��/@�R��|����LdB�*�*�f�<�!嗍i�L�Q����Y Ѣ�dZz�<Iqi%v�*T �K�8�r��Nt�<�s�QY�����/"2Mra��w�<��%�0S4�jf�0Ht�Bc��]�<�TŃ�[;TTA�Z�7_�i��i�r�<AB��5q��i��g\-K.n ���j�<�U����y���ڏ\��2#�M�<� m4���cM�Y/TAb��J�<)���/	z���F�'t�>����G�<9$�Ƃ�ph�#Q=��Έh�<oR�}1��镎�D/�I�Bmo�<���b�b�B[ .t샧f�k�<�&Nƴh`���"p�$��m�N�<A$�	�:��R�	C�]��� ��S�<9���2&ּ��k�>f ����a�t�<�@JVj-���!��j��(�U,LU�<���?���!�Ο3u ��w�CQ�<QF�Y0��`�O�tl�"��M�<����?Ճ��N���s���J�<�c��$�j�Y��;)�� 3�@�<B���q�y�VMA�6���"W�x�<��ME�'�j�뀮�0h.Hԛ��v�<Yr��r�D!�#�,J����g�<Q���)��4��l��Q��{���w�<u4
��ib�ʇ�72Z Qb��r�<Q�'P Y~`�&H>'r ���,v�<� 
(	�GɈe����M/T�ӥ"O<���CF7,��
�6\��A�"O��a�NS8V�j�s�H��/� �"O|j��"�%�?D'x�yc�A��y"m�L�X��4Rv2�dY5�y����� �`�)Lš�-��y�䍘��艕E��Q�tY$+��y��է=זѲR�L8:�p`�ā��y"'�.)&����9�`A��`X��yr	�<0�J�QC74�Hg���yb��ZLɸ�8)j�#�M��yr��C�8��c����9&#�$�y�@� ���m&�6��I]&�y�B
CE�I���M����k��ɟ�yr�X��	��*P���V��yB�I<B#�)��D�>U�n8V� ��yJ0� �86&ݶ~1��h����y���=äI(���oJą!Վ���y�#N�#��/Ċ`:���f@
�y�)�9U9�s�T�QHErD��y�o�>�4Ht����P��D�y���8M�5cnB et �H��y����
x(cAK����F��<�y�JK�,�B�˵�+���S+�y�IC�:m�[��ҫ �j�9�,� �y�D f�%�C��x��$�3(�
�yR+��	�	���O�h1�廇�T�y2B�T�\-��	ozT1�J�9�yB���Sj҄
eH�{�l=������y���5y.�A�u�΅c��%X���y���"
���1��Tm�FEc�$�'�y�	�>�x(P�OY�c�f��@"���y�߶[plْ� ��u9����yR)&?8�䙑��X��1�r ��y ��`��iK��M���1	��yb?�P�8p@�v6 	��)���y�`C$P�)Т/4�ZH���y"���'�<�襎Pc������y�ݙ��Q,U��A�#���\��F>l�Q�]�o�� �n׻�FĆ�#ڞ�˴%�Uk*�k��l�(��R�=���׆>p����H�%���ȓ$���+7�}�A+p ɐ�����%���>k�T(���^.�*q���jM	��ٚ 5��A�+-{����+����@�fYD��	�%'n渆ȓ1��ņ�(��h�I������)z����P@�#fD�<���ȓ7$���>z���0�Ɲ A� �ȓN@����M�'�6�C����$�te�ȓ�D+�L˓��\�D�V�4��ȓ0�hx#0��,QN\�'J��&�N���ҺRF�
^F��9mH<��5�H=(qcA�,���&Y��l��|����#�W��т��O/U��ل�E*Չ��N "��XB��èC@ P��o�6�aP肍Z���1�	I" ��-��}`���QiA�d^R ����t��i=0�
GaI>yLl��E�ʘ	(d��R�Iۧ#�.�U������ȓ�~�۷�^0z�m�Q�F±�ȓ^z���"I�q���c0d��Y��ȓ��@A��Ch;aJ�5�؇�l�|�@�(���W�G���m��S�? �T�W�G�2m�p�K\�vp�R"O��Ô��*?4�<r%��
�x8�"O��SRk��
.A�Af
�M��i"O�,��_M�vL[d�M�PQZX[#"O~�򢏂	X�(8��ċ=o4Yj�"O��P����B����3Ȍh�"O�<�Ǥ�	�F �գ=�N��"OTM�ğ�>\�1y��Z	�,�"Ob,�ҁKZd� ��@�2>}h ��"O���f���<��
۝OxUp�"OD�fm�v�F�����e�� �"O�}� %�6,a��3[RV-9e"O�(�F���{��(� �J�ɲ�"O ��`�  ��   �	  �  �  �  B&  /  �9  �D  �O  |Z  de  \p  /|  Ƈ  ܒ  ��  ��  M�  ֲ  ��  1�  ��  +�  n�  ��  ��  ?�  ��  ��  �  ]  �  � � i   ' �- �3 : T@ �F �L "S �Y �` �f Jp �x # g� � �� � 5� L� �  x�y�C˸��%�RO5d��pJ�'l��I�By��@0�'�F��A��|�^{���OM4ؐ�Їv�lh��Y�&7�C1Jɜ��AP�Hj�%+5#]/AT֝�ҍ�"�x�S(#�t�	0�� �Pp�h�� ���rI�	cUhm���>>O�|�6k�p��`Xw��dU�O������q �P4b�d��A��$lkL`����t
��Ia���9A)�9��=n�<;� �I۟P�I���ɘ(ɼ4��M7P(� �c<w���	���I�x�'���t��ϟ$�`J�4j� ���~���eFşx�	J��ß�ɵO2�y" �l/>�(fLѓXi�q�Wf��y��+N0�*�XҮ t���?I�[�qV��q�՟>0�����uH5�Q�]:ʙ�襟8�@dܚ#�()`�ҵ�,�B��O��D�O<���O����O���1�S!O2�A��>b��'h�/6������������'E6�@ڦ�޴!��	�1�Q�V��9q��w���b�ԭE{��O��=ke'ԥbhE��P�o9Aϓ�OT����f�9���������G�'wў"~z#m(@d9+�nQ��"��u�è��-�O`@����]w��"6c��M����[y��p�Ҽ1����2��W��8c���)�n���3	���B`�I�OѴ�����:�	�>���@�QS�.+g��Rte�'Jt��9�D�Ob�?�'+zI�7��4���:A�Kx��!�'�By�ЭB�XE��,��u��+�',��k��0��I�m1ܩ��'rʔ��b1{W�^������B4]<�}ȳ�Q�l���7����hO�U{���.;�  X��"
��	�$A���m�	؟`���)�y���PtFi�/�1*">C��g*@�I���}Uȡ:��I0	�(C�I�d� �*��Y� ��M�r�ȭ�JB�Ir>��!w�Կ:0@����J�V�?)1�S�c��jshޘuZ<L�S�Z���Ix������	c~��{�r=��eY�� �$��y��˅"ب-�`y2�,��mI��yB�:_���kR/I�n$(�r�GG��yb V�"C<$R��G��h���y��E�=�hY��
�����d+��
P��(���1��3B���1vz$��S�lp��ǟX��K�)��60��қXQfY[c�˳+�VB�=`߼ �%�S�>�M
�q��B�	�?��[E#��'z�p�u�ɿ{�C�	qR*��4l
b�`H2È�@�rC�'7���(5 ҙ?~���DҠQD�O^H�>Q��U�<��O��9E�9KQ����/�.C邕���'��'��6��1�7��� O���T-T7*V"��Qi<J㚝��A*O��1�cd>�;L�,X�@#od�5�rLߔE����*O}#��'�r�'W`��D{ȸ�V(N<;$
4?�I�X�?E�4A@�O�pE0��/ ��XB� W���?A��'�6 �� }���M�,/�Mj����d�;:���$)�s�0�'@�P2��R�vk�!�����=��!�	��t{��/�|�"|2qI�#>�f��h϶US��Ӗm�D~"cX�l��=E��E[
�`��	A�[��8��Z������@���'��O�1��Q�E��1/R$%��
�' h0��|��'0az,�V/�A�t	�*{�dyr��O�@G��h �*w���&'J�p�H��?Y�(�3��'T�4�'.╟�"A��f�(��2d���҈cM9D�dcu�P��x34��2�X���$D�LS@��M�^�:ԫ0�h��=D�p�Ňhܘ���T-z�|X��'D�� bl���֡T�
�`Dꗈ�<�1�)�'r^���J�-�$�.�%��0��j�<����?����S��ݡ�<C��1G8@&|�.)i7O���`�׊R00��IW�ܸq	͊J|!�䗊4؄���F��MR�c�6��P���'l�'=BX��g�62Й�C�\� w���q��K��
�'+��˕��!��;a�I�G�VM�I>���i��S�\��O�j�Xa�+3����DV"o���	H�	��'6�!Gx
� N��o�!5��4S��
�V�����'��Џ��	�X�䅐�I�k�&�S��Ǎ4paxR���?��y���	���5���ʬ�����y��g*. r�I��",2&a����?A��'�D���6Pir�H@�8^i\�*��d��nA���(W���Ǫ�5�< �*ӥ$���Iɟ��ɽU�t R"�"��gk�r��B�qT��5�W 8B�}����/��B��9%�s�ݠ2S�ѻ��T�K��C�I�wĵ�%BB�B)di�@� V\ޣ?� 퓍h�)�� ع�b��!+ߖ3X��NS����D�Iz~򏒟,e��'�L���������y����5�T�B�v,�"�y���R>��A�!RZ�!�f��;�y��Tkj�!��<�8؅�=�y�,�-_��S1C�42�%��P���s��(�7��i��p($(�-Z��(PZ��h4N�����Im�)�S��.M�G����".Si�kI3D��Q�F�P$�a��њe`x��F4D���%#Ю��И��.
�~q���0D�� ��
�1l�thwb�=@Ht��F�.D��� ��w�@�x@Oį d�Q�L.��P�'MU��'
�A���w�C��]�������?ɍ�L��JfQ�)��x��bV0p�`�*��!D�8:#i�!j��)0��Ӻq �a%D��b��-.�b�卆z 5 &.D���)M�j�Rq0��.������-�O$��Ig7��+�7��s��_PƢ=��)r�OT�X�F��B�t�� �O޺��'4B�'�F���(\�R��š�a�z�'�y��U),*p�KSq����'Q�P%coz���銫DNr)��'��|!f�R�i�L�S-��-��
��dGb�O�j,�p��:tDɁ����P{�u���Ex�Ot�'��-"d���%��R�6L�%D�B䉔�+*׆L0������!8v���'y荺a�c��y�e� ��u�'�T�r�`�Sd��u,�u�Y �'�x�)�N�W�δrga�p�$+O�0Dz��T&,IL����� }�F����5"c�99�
��I��%��>u�â��X8�{sk�X{��3b�*D�li�I��Ut�����3*Ȅ�h)D�,S��/qÄ	���[9����<D���'�$��r�O�}���&D��T�;���S�KH����&>���r�'�:���' �@A�צ���:���&'{jqb���䓧?a��L�\3�ޮd�z���ET�=�d�{q0D������0^�'��Br���/D���	�Q�`)�QcLr�4��,D�PqAψ!8�I���8���P�e(�Ox��I�ls$%�R)��N������0q<��=���c�O���c'��=H�Z�bK�|T^-���'b��'�jx+��C4\��[����
�	�'QP�;�A�5��x�%*�
�b�	�'�$��E��t�t`fC� N�N0��'
�A���r�@y�֡-M.����d�~�Oo08FC\�0��Q�v��"K�����:(Fx�O`B�'����C��	;��v)n��e�!_�C�	�P<�R�X�DǤ���*�;,rC��&��0g�ˁ}j�s% ={nC�	�t��X#E�#M�9���$:��B�I�h`���ľW�TYG�Z�mG�ʓl���|�Q�f"�<yN�#a�DP;�LUyʇ6�B�'Dɧ�OK4��G��`ʨd٢­d�40��� @��D%S6%9�)RE�2S �P�"O|E�3��&��`�����C��	"On�V�I�/Y��ң��b�|z�"O�� q|�92�kN#K��`࠙|�1��΍�W�E����e%`mx�K��~Q�I`�	�����ON�R l/��i$�^1v� ��V"O��nV�H	�r�ۃ�$��"O����� `6�iӳGU!xᆌ"5"OL�30ʑ>��|qQ��&b��,ٶ�'Բ��Γ&C�Q1��c�DxR��&�ўLIK6�'!�ݨr�ؖN���Da�5^q$	C���?i�j�lx1����V ���a/׭%�D��1����ͩ�jȃ7&�'m�m���0Eq(�V	�Tc�fR� l:�ȓb�d9�'O�/$zx+���j:�D� ڧ�$Icf�6n�0�+G��,�F}��-K��"<�'�?����D�"*&<�7� ���!�ƞ7!��J2b��w����Nh0�G�I!�>0Ȉ�҇� eR�,b�`B�u*!�dH*�"��Iţa���DJ�6�!�d3`�$ٓ��t��ъb��{�剽�HOQ>�'�<!�X��dg�C��U�BA�<��M"�?����Sܧ9|Ѡ�\�0��M0�eƪP���ȓTp����r|�X�2�C>U��X��@�n1Au&V9���J�9��t�ȓH�p]��G��j��� �L	5P��$���.aY��lV��
����$�D0��$�71<�$G"~P���F�k�^���H�.�|��'N��Oծ1��5V�,�F')
I�ȓ+;�4�*���r؁�l������).>��G��@�f�:��(���XL�G	De�8�P-�;<=�Q��Ɋ�?iƉ��kX.��Vhڔy���a�Xt�'.d�َ��N2��!�uJ)ق𰫉�-/����O��d�/7b2��%g�]&�0���<c!�䇗=Cd�:D� %�`Q��u\!�d�!���
�&
B����0@L6hR!�˹;��ŀ��Ph�,T��?">џ������2G>ܨk���,�����<< ,R�O���O���-?�A���=-)���0P�b�D_�<Y��s�`��%�[g��!E�Z�<9�I=�tX�G�k գV��W�<c$S5�
�� E��eF���Y�RB䉪(�nE�󣊺�PX�#� �U���|��LZ�A,������ ��K�Sy�c	��'^ɧ�OY�Pk��!x~����ʗW��-�	�'~��ir�Ӭ�\E)`�PDd�b�'p�X)1�֠�ݣBO|N̽�'>zUC���cY��1�Z�%�b���'�H�cE쒛U5�m�6%V�2�܁�M>����">��t0<q�EK�zĀD����45���1���OB�?�''�����j��j��H�C�(K	�'s�	�S[�,;F�V&@1l ��'��8�sf�8
~$��iG�A�4�	�'����A�"Ore�׀c�6��� Y�U�fPc*X�CdU`��E2�hO����Ӫ<زS �hvD*'��'vcxD��韐���6�䲗G�5A��I�#Z+vB�	>�=���2i�t��냜n�B�ɶ`W�`	A�H*z�ah��*2.B�I�Z����I���@�b�
!ܢ?A�5m`��$��'UV͊s/��Y����"2���S��,�Ib~B��N��k��]�\�R͠DCִ�yB+�6%�dy�&	
�,���+X2�y
� ��	�.΀y��o�Ը�xf"O8T�Ц�1g�*�x�0]T�
@"Ot	�n\�ȉ��)dZ>���Q�����哮\�%��<Pe�g�]#}�0ʓd��R��?AH>�}*�I��*9�0�n�b�����
�]�<�5C�v.�j`�ę%��mc���X�<���(z�=ku�?8��m�%M�U�<�L�bP�\���6+)�؋%M^M�<��
;F�E��
�W3 �h���d��1��O�� ��OȌ�G�G����)�������'�'���>��GO
e�������t�4�RWkKQ�<�!C<`����%�ȑ5�۱�V�<ё��j%z9�6��X8��U�<�%"E�'�%I�)� �~���C�Q���R�b�ȼI�/��1"�&�D���D{l�͈�܄bFоhϸѡ���t��1se�O���9�O�I+�F���@׮D��"O\x�rF���0%�sgM�H<p�"OH\ȰA��p!���s䌲y'�yc�"O��ٔ�� iiT$ #�.�<(�g��%�h�|�	1�Z�3�<�8�Ʃk�x�$�'�Rh���4�H��O@�)�Ո�B9$l���?�~\�ȓ4�z���V��B�[e�Q_����kP�}����$LAJ�;�aJ��d��o>��p���K������Zذ��G��5�Gn�*�<٪w��|Ӵa�'T�#=E�Tb͍_��Y@���i���J������ƈ���$�OƒOq�<��sƁJ"�� �O%{�<b�"O�U����J��AK�,�t�p"Od 1����L�2��c�Ɲ'�>�*�"O�X@ƛg=
���n�(���"ORs�ٵY����Eڿ$tX�(�|��%�ES�i�9�4��'�!*4;!g�W��(��e�П���O$hp2� �7�<��+�;V9B�"O$!�E�ՁZ���S�TIX�Ӱ"O����bO%���1j��:ij �"OԸ�G٥JaHвh�F^�M�f�'y*�$n�ܰEί5��@3�$Dvў$r�O$�Z$^�	4�ʀ/ƐZ�"Mm������?y
�M�$�M	u�dP��T�[�&Ԇ�9~B�B7��_��Q2�ȇy�Ȇ�I��AQ �37��L�w��Vt��ȓ1Ŋ����Ak/��p�O�-��HF2�-�'![l	Cw��g ��T;����I�H�"<ͧ�?�����AM Dz�&�#[�����m��X!�d�3p.~Ic��_?C�̭��k�`�!�$K*I
P��$×6¸���a�,�!�d�	�Z�@�B�+,�*ڒ��9%�!�� s�Ԙ��+ �X�����<�創�HOQ>%���S:K��s7�/M=H��<��#��?!����S�'z�ހ���)\I!mͺNu�]��Eb����h�G��P��&_�^�͆�DD�)�b�ԉi�Fe
L��[3vy�ȓ=���H��ڃe�0b�D̙��d�<�!'R��t���B�:�d��g�g�:��O�#D�O�$B䉥���2m�"�&���'Q�'���>Q�
ӹa��S�0Z��-�`�i�<��L�>=�p`���R�B���e�<���=gj�1��M$n�D!K�B�^�<!��1�~� �G�t�D3KR�����f������ (�nzBȒ#~�E{�kF�҈�Rqq��Y�b/x�H��IH�y���OX��5�O��b@�͘�3�ڗ
5�h��"OFD��ɓ	"<�A[ �`�)�"O� @�8fIP��h�rr�H�0EY�"O���p��m��H���`����	��h��B�M�n�c�ʚ�6����' &IJ��4���$�O��3�V`�nLq�&2���f��=�ȓ��1£Q2M}8Tae��*(��ȓ=�L	��iÚN.�$�Q���Ԇ�0���E_�pIH�
��V5���uz �2L�f�K7O-�$�'5�"=E�Th�M��lX�iB�l���Zb
����v��d�Of�Oq���S�A�Ct��	��O�o<N	s�"O�q��@�(�Jj�4�J�"O�p�"ءiu���ɘ.V8Ȉ�"O�2k�2Y�� +،~�HXf"Ot�SF��	�f!2c��N�
ĩF�|�,*������M�c�;�f�鰅U�T�L��@�	�����O<x#��&aY�ɢ�E	�)r�8��"O�p�%N�w�2�TNNcS�a)&"O*�Av���E���c�Y�O7�h1`"O��#��0G
2qp'I�C?���c�'Yh��Յ-tbhҵ��(c��	
 ��(�ўЉ��4�:8����X�Xk��W�t�����?�t`�X�ă?"�ڭC��]+YB�ȓA����MR�~�
<�'j�*g��؇ȓ_�8�S��ݫ�r9�'�	�{WJчȓƖ]׌��"�,Dσ�
dr�E��#�'c�60�H�0����@�S�°���q�#<ͧ�?9�����^<U��TBSj��T���� lN�u�!�� 	���vmD�g_ؠ��+�22�!���Uo�P�ǫ�U.P "� ��a�!���2*�`��ǌ1���`gI�!W�!��͌]BxӇ@
4�VX!���剠�HO>}�WՑx�� ���)r��]��nY֟�O��'{� I�O��'���RU��&h�^�@Fꖫw%�����|R�'E��4o\fу',	@��	3���O�!1ub���KWx@=S&�z8��Hg���(a�C�Q#��Ozt pB�d��š@�Ȧ����� ��'&1�R��uK�H�4�j��[�U���pR�����=+�ӆd�:6��ab!&��	�(���OLyr��	M.�b��T&n�hUr3#����D�7Z����O��?�	���� �/����2c�"���Aޟ0
O�Hp��,��Ku�X��S�O)�HeG�, �5�&#􌩜'&*Ѩc�l�Z@�"Ă�}N�?-���׷p�Lia�	"W#\�(6�s�`S '�O���#?%?��'p�hI�*ʿ��a��[�4J�@	�'Hz��$�*6�\�y��ܸ���1��$�m�O���R$LK+jr�(�f�!��V.D�:��O4�i�O��/�Dۍ2�bL*��[	ˈ�y�IO��B�(vb^БF��	?�f];�
��ܜB��*S`<h���2Z�8��wE��]_�B���đ���N1���T�&=~B��&[��C�M�>�y`��T�G����B�����H�`��62�؅O�d]F-�U��O,���O�d6��ӹUWh��"I��K���YR;Y�~B�	�`��Li⌙�9�`� *��.h^B��	-�H�	j4=��X�2B�I�
�����* )]$)B�ɫ,^�B�	>��c���\Z��G%/;˓`ӑ��BC�6}�@�;/K��p�f�9pX�g#�'�䓓?��0<i`ߍe��� �q���A���S�<i��	Ǫ�6�f�hDO�<	C�BAQ&$+�O >aЍZ�-b�<�,�U� a���`��|
0d
ax���/O@�X��F�IT(pmާ!�f�8 ���o��������n٫,:�����u���������� �f�("CL�L��!CG�}:0,�ȓtҸE��� 	�8D�UX�l�,4��S�? �eHchwѼM�dbS<_r�U"O�Iٓ�CJ�Z�i�&^�C���蟆,�J1�t\���.e{l����=�O��)�O
�$ �56ȑ�sg��x�V�X�A��6�zB�	*\�]z�BAg��(5���TB��
�^���d����Т ��qm,B�I��\�!!UQɞ!���%v\C䉥B��Y2�!�J��	y���vj��dCZ�������oT,�^�*�B�1i�cA�O��:���O���,��5LL:�r��}���F �sLvB�I�"���RBM��#��NDC�Ɂ4Vm��5��ج?~:���o��|{����R�ƥ���<W�t��ȓN��T��C�0[+@y��%�5
`���'<�"?	Ӧ�g���,�������H�b$��ꓧg>�'���'.axB�T`zl�����^��pӲ��4�y����0ǎ��KƳWD�"�ۍ�yR �����P�KN|����n��y�j<Rf�a���K����E���$ry���i��1�G��J��3�@W����O&��<���kz��3����l����)V����O��xKB��>�©S����;8�@q�!�����&�d����|B�NЗz,!�4�W�4��ɠ�~��W;���|�t�l��R+ �(h�E"P90�0��󢝣���DD�d��KR�F�O��$2�n.��I3	ˍ8�`Q����]��RB?ٌ�9OR5�5�6n2X{�їg7b��e2[��-��"�PD�O���On�I$�Q�^Δ�j�.�a;��F��O4,�v�S"u�>=�]���"p �V��8�	�:�.�'��'xHآO����4J��� �Nז�
�KN�];�a�'6,]�I�x
���٨^ �aRG�2U�V����W�3��5��,̔U�O�s�X:�+>?	@��p�N�t��>��ٻ��AV�/O�HW���3�ӲB`�E�%&�?
'���ܘMP"�Dۇ�~RF�(���?�	:6����2���zD��+��@h"����'lba��	h�����*��=<)2#�1_��B�Ɏc���ᢍL���}Ba+
?@�B�$^Eڍ���Z�"��%�2/�r��B�	�s�`���ՅT��Y2D,%fB�I�~;����i����27eBB�	C���̝�yN�;Ӥ �cB䉸qU����N*@v(k i_	PC��,A�R-:d���J��ɖb9�C�I��й�MZ;.B����nC��L��(�� �v�>�P�$ԥp-C�I�e�
@+f+\/�t�тc�[��B��?'��]�LΖoJ�M��ĲR7�B�I�O&��+5&�% �9��8lX�B䉍��lJ�)]/W^� Â���!��#?����?���?!�[p e�� �c���<W��)�i�b�'Z��'>�')r�'f��'�0��֣&���aƥO(jغ��e���d�O����Od���Oh���O,���O����̟|�6��3!&m��X���¦���ǟ8�I۟X�	ܟ��ğ�������#��l0n�AS�
>�d�K��ז�M����?y���?��?���?!���?	��ZI�X���ϦJO8���0����'�"�'��'�r�'���'~2��8���ps�^8(~�	3PB��G��6-�OD�$�O@���O����O��d�O��dY�B����ʲf~i��_"9!BAn���H�	�����Iӟ�������	�0���ٱO�#Ӿ�H�	��?�~|��4�?1��?Y��?i���?y��?	�E;��nbԍ��K{N���ÿi��'v2�'lr�'���'���'��ഩ�B�zL�Db�	Jzp�
u�j� ���OF���O8���O���O��$�OT�Aw'ٴy�<�Ec�_C@��`l����	˟��I͟|��ڟ������	�i@fH�B��4�Jb#հ;xt��ٴ�?���?1���?!���?����?��qZ��t��]xμ�����3��i\�I��'?Ib�̘�CA����P�f��D�6
o}�T�\��D�'�?�'LZ���e],M�J`,A����s+R֟h���<��O2��L�8#�'���ÝA���K$�w���-�28O�e��.X�ў���<lǿs���I�������'e�'��c?��	|�? ��UjФ)� �r8/�L��"��<)���?�'$�.>0dQ�B�N�U29:�ڹu!(ʓ�?�e	�h��1���ҟ�cR1O�l*�n���V�B�
5c�Q0Q���'b"��:&�  ��d�g�:K���c��O���'��I�p�?�'ڸ��v�^�����2�D���?i���?���_5�M��Ov�Ӆ��^w(�\0���0"�TJL�"�A�����ON���O����,oe�5`�m>�0R�<�rY�x�'���	��6^͊D+]�dp�A���Q�.��ʓ�?����yB��h����i��8�<x��E�"a�oܠn����?�p�O8�I>�(OD�[v��3�V1��ҕM�l�4|O���'���y��ʒ����=G�"�'��Oʓ�?A��y��{c*���S�����%�:�)��4��$��i�֘S��O�"�����ݙ.�ּE��=J`b,
�:���D-����dK2|O����'p�H�`��O��$�O���'��S�`�<�㒓=�|x�K+B���G���<��O��d�O���P�L46�5?��5����G D�K<�I�J�0����g
/�?��)�Ī<I��E�:��� 	�(�L-㶄�4�Oh�'��'�r�?�y�([�f�V�C�N�cRp��u�<1,Op��O��]���>���d�9d>1�Z	R�X��?J>D��Fay"�O�4�	y��'Ny�O�)�vHKTK�;�t(���'�B�'���'��O��	��?a �Eg��T�^�{1R�����T��ݟ���b������O�KSl�������`�yn
��QJ�O2����7I�7m ?���Ƚdf��Sc�D��Z�bͺ�,K��b�9�?�-O��O���O0���O4�'9z�c�jF�*蓀$����O����O��$&���O���f�g������]�2>(��G�O��D8�D'��)UN87���(��HP�x�vyh�\7l�(�U��OE+v	և�?�V�.���<�'�?�%���:�ڶ^-K r!��*̀�?1���?�����dE}}�' r�'n �@3�R$J��1k�6|;$�j��Ģ<���?�M>!�^2}�����i�	v��� X)�򄖧S& 1Q7���e��i>)j��'��5�.��)�+l	B�)���U����ʟ���ɟ�	w�O����2i^=���{M\x3s�#��"�>I���?����'��d^�n��� kB��H�M��	�'(�'�j�H#�if�i��I�V�?�Y��ڨ(�X�)&H%/�{CMS%�'�Iş��Iџ��I�����>:.ĈҖF2������"��'F듗?���?�J~Γ4M�@#WH�`�p�e�w,�/O ��OړO1�2|�蝅p�R�a#�\8}�y;���3:�7MTHy���LƜ������$Ŵk��(�s
�HkRx3VJ��-�D��O����O4���O�ʓ<��	�4�X ��ah���=נQV�럀��G������O���t��k���T�d��N{��d�/��6�;?iP��@��i4�㼃e
�2�=�j�>]�@���ߟ��ڟ$�	��`�Iٟ�E�T�ɯrp,\�C���87�;�$[�?��?��Q������l�	O̓j�>L�A��X_|$��(IF��$�$�Iџ��	J
H�n�T~������D˖j��cؑ� ):D"�1��Iu?�H>�)O8���O&���O��KW�z�ʤ!��=��ݚ�F�O��D�<)�Y�8�'B�?m��
Ƈb͘)�W��a��<	/O���Od�O�c�v��gܲr�(��m]��9FkG�-� oZ���蟖ha�'��'IjL`�b95>\)"%g�_z��A��'d��'b�'�OB�ɐ�?�b�� �%�'Wb؝�v��~�Z���O����OF⟀�'�b�[� � ��k���(b��'G�(���i`�	�ED:P�r؟@�'/s�pr��`��JE
��t�����wyB�'�2�'�"�'��?��3�%I�DU �	�	�%S}��'���'.��y��'-�DJ�g�k�G��H��(IRj��!r�'{�'��O�BS�i.�$�H`�z���Oc�}�'�I�dz�Ƽ�"�������D�O���3�L���V�L�`�ue]*���d�O����OX�g���Wy2�'�<9���,�0=�7�B;C���1���<����?�K>ٗ	)j��q�V��H�  [bm��Z*k�x��K��(	�i>u�`�'[�ΓZ���E�<bۼ��7/dFjX�	韤��˟l�Is�O��dY{���w��2h*m����@f2,�>y)O��8���<�Qo�9Yk���΍�i�7i�֟��	ɟ@�əCx%m�g~aF�Q�]�'Wn���W�,d�~� e9Gph�I>	(Or�D�O����OF���O��p�*D46Ȫиa�5��͍cyb��>A���?i����<a��B�V��ܘ�h��4����d�O���.���!�|q���F�D%��� Q5��T�i�h��'� ����a?�I>y+Ol �D�@�1�����"�?"6�+p��O<���OD��Ox�ī<y]���IW�? lj6g�s�J�pPV04�,rD�'U���<������*�$ԳT�ݪ�1�e��>ix��x�i��Ɂ?̤�V�O�,�%?=λm�⍹�	�[򖌱gB�����؟��	̟���ɟ���j�O�xt�n��H�ɢ�-p�� ����?A�������	ʟ��<�T*@0^��j��B����a�K�|�I��T�i-7���R7M/?��¬��R�I�(�Ǜ�l�f�""G��?�D	!���<I��?A���?i�o��M�8p 	b�NZ�M�3�?	�����|}"�'u��'!�1?���G�ξW��glB�.����d�O��(��~z���0����T��|�FYȷ-K�UJ��7�H��z���O
�I>q�M�h�2|����	j�8�
��?����?����?yM~�)O����2N�(�u��-�($�fA�%M]���Ol�D�O��|�'M�N� �DȘ� ӂf���.ɘF�2�'��a��i���(&���i��HA,0�SK��m� ��'�8P�T���I�����՟��I쟌�υY��@�+#CM�JA0� @��w���ٟ\�����&?Y�I�Γ^�fH1S+\x�ʐ�ɓ8����ğT%�&?y�����y�����E��RR�����4!D~���^ʼ�)��O��O���|�����}��F�>{YpU�#m_�Bz7�'��':\���O|�d�O��V�|`^��7m+Li"[@nV�kE��x�'����%��kIץ)0���Q�EjZ˓]���Xp�Ѷ(M~"P	�O`�' 0��n�',�8��eX:C�����?���?���h��	�` ���̟pn�%�I�1� �dq}2�'M�'5�O:牒����!��Ap�mR�A�g6�D�O���O$�� p�Z�Ӻ���^��� L�?> ��A�8$>����Y�cT�O4��?���?1���?A�I^r�@Ab�y�.��J�`�(e*O~��'�r�'%��T�'x� ��e��d�g�4�����Q�������&�b>�����W���'��!� �j �[�v��s�]~yB�o����ɺw��'��I<;�x��g�J�+0�Pr�NG�n���	˟���H�	��ܕ'�@��?���܎	��ai��O��)�s$�7�?����'��������<�¨:5���F���tE �B���秊�'O��$\azJ~��w,j�
X�<�и�����Q���?����?����?A���*��$���f��;�bּ���1�'T��'e:�����O�b�8�d��� �q2�[�LV�T�q�=��O����O�,	�E|�N�s�^YQ�(�m��E��!�/+#d��v�H�j����X����4�����O�����f���Mϱq�Ȼp��9�R���O��t|�	jy�'��Ӕ)ߎ-�
���%��.vJʓ����O���8��~���#��ЁO���E����> X2�A̦;*O,����~�|"IH(~�LH P�DZP�I)��	M��'F"�'Y��4T�L`��|aj!�Ѧԛ5<n�(@�@:8��������Ɵ��?�)Ob�dQ�0�Yȳ�>�N�cc��8lH�d�O���	g���A��˓��� pص�5�T���O_TD�c$�'~� ��䟨���x�	Y�4k �	��OF#y�V\�Gc�g��I������&?�����ΓF6�)"�A��D�!�Ϲk�z��I���%��%?��f��A��\��DKR3{H�����hk<D�	9N�$a���'5��&�d�'���'���Rc�s"��C���)�$�'�'��Z� ��O^�$�O��D�Ck�l�t�μyXTa���qHr⟈�';B�'��'{rԸ�*�>}��D
�KF�[�K�X�l��+H'&�L�lI~�O�����y���bR���e�>D�p�k ˉ��?A��?)���?��Iq�\�$�F:1�(I�K�\��D��O��'[R�'���$}���i]\��P0�(8 �U�Ba�OV���O>���	6�??� ��~��	~�Q�jY">]m�HÚ#�� ���'��<����?	��?���?4�A�=�~$���Z�
�ͩ�O�?��Ve}Q����~�'+��1��''��S@��1wEJ�#*O�D�OؓO1���*�e�8)�lQ�4�� ����Ri B��6m�oyoΆJ� ������Ė��&e9�eP�yj��36/��H�R�d�Or���O�d�O˓��IΟ Z'E�>/?�HR�B�FG8J�W��h�	I����$�OF��`���4Txx��a�eB0θz��؉Tu7�"?)��h=<�I?�S���GB�X�ĠU�L�]�`Q`�@�	ş���ɟ�I͟XD�dB/}eh��.�<C\47`L�?���?&W�P�������r���l�� H�lQ�D V[;�&���I�����{��n�M~Zwˎ<�CH�af���(7���3���6�fVk�	Yy��'�B�'⫏�s�"Nu	`jN��@U���'h�U��r�O��$�OZ�<Z�-��)�F�`aM��fҮ�z�yy"Q�@�	Q�S�	�qf�4:ω�@6� S� yg�Y�֜� �T����f"�LP�	�9�m�⌌'������^4�%�I⟈��ٟ`�Iv�MyB��O� �k�LMW��:����Ym,�g�'��'�����<1�4�I��ċyh,B��̙������?1K\��MS�O`��b��zK|2�
�O?�	����Z���OKɟ��'_��'
��'B��'��ӣ5�z�z���F�,�vE\"O����'�2�'�R���'�23O��G�ÿ*$����ԓ7�\�s��'�b�|���D
*��6�O|�TG���Y��aQ<"j�պ��'wt���P��#2�|�Z���I`��6�@��K�e�����I̟���|y�G�>����?a��YR���E�(`$��`�B���}���P���I̟X$�\ʳH��vK�����V=�{r�wyۼ[��	׾iZ�i>Y��O��ɼHd�t��b��&�O�M��D�O���O���0ڧ�y�͖r!0���钐- �p3���?Y�P�d��۟(�Ij���y�nO$t�����nC�X������?A��?���z2��P�4����?
�RxI���u�hw��c�
&�n%/A�o��p$��'�'eB�'��'������,6L�p�M�*Д��P�HA�OR�D�O ��"�i�Ob�I� &ws�9�(T�w�6�Q��<A���?�H>�|B��؈Qɐ5̳iZA0��]6�l`��Lx~r胶(b&��	2pC�'c剐r�ܲd*cQn�h CHڥ��蟠�	ǟ��IX�'QF��yr.��<�ЄӇ�#�I+����?����'r�	џ��I�<iR��:,�� ���:Ppu�rF�=BZo�M~�%Ke���E��;��A���j��-�7LW�+O��iE�'���'�r�'�r�'�>����"� �__�a�w��(��I�`��Op���O�D"��="�t����P�P�QQ�+@�:�O���O>�ŵB^@7�5?�;"ʬP�L�	��u�P� 5� V�\��?ɰ+<�ļ<���?Y���?���i"�k��D���k���?A�����M}�\���	j�t���>���S�1d�4��\��<��������܄�0��6=?�MQ�hϡ2�LA�X�* %I�)����?�� �'z��'��`�I�!�fqKrl�+P�l��U�Z��\�I���Iϟ�&?��'�D��}m�c�%� �@���S��y��'[��'�O�˓�?I��mP*�q#���y#�A�2����?���kθD�޴����!蟬A�ʟ�Ћ3�[	!�B\��#�|h:ucC�'��ϟX����l���� ��H�Ԍʇ �B������G�o��IП��I֟l&?��	ޟHΓM����C`Y���m�� /�,0�I쟄&�0&?����ܦ���!�r��.�u�ѩ��Q�p�	9\��y؝Z �|%��i݁�'�?���M}�t�T��4S 8cJ״�?����?!��?���OS���'eb�'��m�c+ �b%�p�>�PFJ�r��':6mK�g`�d�O���G}�4��I�B(,)�T�Aq���@���F�'�rK����c������:��{�*�ə$�r5x�ÂnN�H��6)����O��$�O���:�'�y���,(��V"~2�駪4�?	�Z���	��0��Q���yr�\�wU���!k��_ؘ��&Ƈ6�?y���?���|x�D��4����,�[&���;T��/R<x*����df���f��������O��d�O����O��� _�>�J6	�;@~-k�oZ�4,B˓~<�	�������&?�,l�R�	%'T8dZĢ�H1>)�1�'A�'�ɧ�O�j����.-�d��t�؛>V��3�:�ź�O~�h��W"�?�uc6���<�uS>�
�3�Q�i�Z$�q�-�?Y���?)��?������w}��'h�h��"H�q#�4'za�0�'L��$�<���$�;( #�ꑗ5�LH"եڇ7�՘��i��	�j)�ț��O�ȁ&?�ϻ@H���+�#x�����.z�4����\������	��	T�O�(yB�)h\��&�)� � ��?���YC��XyR�'�1O����C�.��h��o��@ו|��'KR�'�t	H�i�	@=���5[J��.Y�[I �2�Q+�$>��<ͧ�?����?��*9x�:E�HJi���G)�?a����\}��'��'2�ә%�3cA��E;P 颎ĹQ2ʓ���O���O2H,2E�ȩ9��Y �)Q2	Q
	0 C�"8Y�y*���������lA��}{B�O�c�Oм{J 1	���HP����OD�$�Or���O<��2ʓ)����~�@��iá�dݩp���?���?����'�I�������K��
��u���S�d�Ɵ��I�_wZ�mZD~B��� h�a�9Ɣ[���2P��ڄ�^/���D�<Q���?)���?����?q͟ Y2f ��j���r�@�;=��e�ʷ>I���?����<)���yR	6W�	�aJO-u���c���?a������'xΕiڴ�~2�zj��v'�'kڨ�bC��?��`(hv��IW�Ity�O��k56�%X�,,���c1'�X�"�'��'8�ɇ��D�O|���O�$aeC��M��b�
���6�	Jy"�'n�|"�Ӭxn������YW�* cмR�	�SAd�Z���¦!���J�v?��'8L�W�]0|���2j,��h��?���?q��h�b�)� �`�$��H��=���OP�4X��'͜��?���?y�<Ox$��ʅ'<��p;�U���@��'m��'h�iK2��&���A�ᄺ;�4���q�m�*�V���E�>od��|�U���I��P�I؟��	��ː�+�p�Yq�\�K�V�ayң�>1��?a����?iP/�n���A�&|���ߗ��D�O��+��I�$ElN�Pt%�Fx���`IA �����@:�	� h�y��'�t@&�|�'��P:u�?KD�#�JW+Yg2h�S�'���'�"�'��Y�l��O�$�Cir���T�G�P\��j����OX�Ȗ'hB�'���'�V|�U�R�!���U�[�z^N�#@�i��	�o+�=�C����jۮF�a���O�eh*ɔ������֟��I��<�I���D�o�b?�0�G�-ĭ� ���?��?��S�$�I�\��E�`޵��+��^���E�A��" '���IƟ0�	�[<l�a~���w��u��GZ,W#l8�ߛ��$�k֟�r%�|R[���쟔�	�� )�fH���ռ�
%d�ߟ��	vyB�>��?�������J�A1�Wq� �Ʀ
`u�_y��'��|J?��Bŝ( �&uY�f�<?Qx�0�IT�DВ�U�p���z2��O��J>a��*�Ĭ;'-��uaT��sM�?a���?����?aM~R-O���I�0��s�k� j=�Q�H�-����OD���O:�$�'�b��nn�)�CIѹ> ���F�F�IF�|lZd~�f/:���S ~���5�h�J��S�O�^@�
���(��<q��?����?���?A͟x�HG��8�8)��CDϒ93K�>q���?!��䧝?��y�a�(,�PS�̞�!�j���?��������6�Oȑ�5��t���� ,Mb�'P��ӑ�m�6� �����O*����Px��b�&9ǈ����<���O����O��,��DyR�'���a�F��);�bF�: ����<���?yI>�*�|��;T�!49��{�[���P���x(t�];i����p�l��IEB������k%�@�O�M���$�O��D�O���$�'�y�ڹop��`T���1��]+�E���?��U���	ٟh��d���y"d�0m
M�4(bb �ȫ�?	���?���=�F�ش��Ċ�0 ��)���uا G�,#��N!.���87�����$�O:��O��d�OZ���9Hp��+���`���Ȝ'�6�!�I��d�����%?牽G�^5)��V��-s�C
3
�4��'6��'�ɧ�Od��	��Ѿi��+v�V�e���3gC.:��OTu�fN[��?�-�$�<I��Ŏe| ̱�Ŝt�:`�ch#�?1��?���?)������i}2O|�FfR#�=��I$q4Pyq'�'BR��<����$@���:���!���Qa*1U����i��	���,��O�M$?	λk�V��Æ9C�D���)\$����ܟ��I͟���ϟ��Im�OB��q)O�RZpe­~�|r(O\��H^}��'8��'F1O�ɡ��
�B��ŋ\>Y�4�`��|��'s�IoLou~�@:�D�+B%t�.48�E�o҅9�,՟@B��|�\���	ٟ��	���3D#Q�K0ܝ�0N�bV�]a��G���Imy�A�>�)O���*��͝�`@�!�q%TAϺ�@��cyRR����ӟx$��O����CY�j`��Aa�3Q �c�K�&�F �fD~��OZ\��I0)�'Y�i�HaJ�ꑀE�(b�B&�'b�'!r�'��O�	:�?��h��B����0ꂬ����c��㟸�I�P��|������ODEA�+w2����2C�
��m�<�T!��M+�O$
sg�.���!��	���<�C��4@Cֽ�"P۟�'�r�'M�'���'��S��hC�Ƒp����	�	<��}�'6��'�����'�;O��;W�܉`5����	��q��'U�|���d��4���O�4���m	��:��!����1�'ɼ ن�[�8BA�|�Q��S�d*��6rm���3o��hb���ߟ������syR�>A���?���x��E�����R`x�$Z�1�����T�D�I��&�DJ#i3Z�ұ�2Ie~�1��DByBKG4j�(� �Ø%�O�,��	%��$N܊�1��!K��a��%�c���'��'��S�<Q� T����f�����t�&g���$�Ob���O��0���<��+�1u,bX"�ˉ  ���������ş(�I��r o_~�-(�����+�-�
 K�tcqō)��p��LRe�	iyB�'g��'���'��'q�L��V����h��Ʌ����OX���O�������b}�
õH�VСe.��;����?Y����Ş�4��G%�|Xl-) ȁ
�|�����M�_�P��G��8��$?��<�*
cID]����&� ]��9�?!��?��?�����	m}�'�4a�Un��z�+4��$� ����'�b�$�<���?a�'��X��R:Ix�X&�D1Z�U����M#�O�h�U�J9�����d4�x�3͗�,T:6�,�����'��'�B�' r�'�>� ��U��%Lg�yчw�n��_���	?���Oh�D�O�c��cN�&^��D�T�X�W[�hz�j"���OH���OVx�	bӐ�
�d�3�o����9A�K^�*x�+�&��S���������4����O�� �̈��n�N-z0yC��)ef���O��M�Iӟ��I̟��O-�Y��N� �
���!4��!�.Ob��?����S���8�8Y�7��%bd�ag�;V�L��A>y-��3�O��	B��?�gb,�d�� 8��rB��m��q�mC�8�����O��d�O���)��< �'�8� �Aκ8aL91�����?���?��^�t���uN���C  |�	�c&F�n]|��'s�Aa԰i\�	:
�(��Ocb��O� \1�����c�E�/f�U	�����O����O
�$�OZ�,�#,\�[^���G.Y�E�ܜ�&&��$�O��D�O��?)�I�<I���)!����=6�!T�����{��r��L�anZn?�eo)Mо}!%�G\�0�e	 ԟ�Ҥ�[SWbLq��RyB�'��Ȁ|A�eA�+N�EP�E�͞}!B�'�b�'�I���d�O0���O��t����6lˆ\���5� �	wyb�'���|b�Z�qE�����9U�<� ���5U��	3�T��B̚��L~���h�<%���ɴE[*5!a#"�l���؟���۟��Il�O��D �SN�8�/�([C��G'׎ie��>	���?!����'i�dZX}J<Z�DM��*��K���'���'�� �4�i���z�J�!�O뎚�|m�Y�bOՕq<�;B��'�'��ğ����4�Iٟ�	�$�(�l��Pǆ�k�(ߞU�8�'듼?A��?�J~J����i3i^)L�$�89D-�/O���O�O1�b���eX�U�&T�J��؆ŏ2.�V��H��?3���s�Zy��9C���E��*i�A�BF�2�'}b�'M��'�����D�OiI����P���@���:}6T@0��O��:�IXy��'�2?O�*��;B~�� �7	����6@����,`4��
3��d��g��ì��tYRu���A�!��O(�D�O���O"���O�#|J7��r�L8�������a��\�	Ɵ���O��'�?	�y���f;t�3"m׷(��8I�� ���?I/O�
ujb�d�la�y;����VK�4��*R.Cbx��_
5����N#����d�OF�d�O���ӊd?|�o�vҰ���i���d�O@ʓ\�I柌�Iٟ�O,���?��4���Q�WHdA*O6ʓ�?A���S�)��H�@���{(�0�3ea"y�D��n`U��O��)��?��I ���j�c���EnMy�@�!��$�O���OL�d5���<1G�'��cS�D�"ľ(qW�:H�������O"㟔�'�� /�, �׹c˒��Pf�";�b�'n���Źiq��9%�Ƌ<��
�0ţDi�Ā9��e�%��d�<	��?���?Y��?�ɟ�I�����sĦ��AػZ�$R���>���?����䧌?����yRHL('��}�t��w��H�/��?q������ڤN뛦�O�i2(ݵaj8����D�����'�҅6ƃퟴK�|V�|�	���ؿU1����ް�B�%L۟����p��ayҪ�>����?1��qX�$��1Gf�d�g+Q1+�� ���W�h��S�-V  id(=3���3	C�� �A+O�l����BʀT��,�)�&�?��!m��#�π�7�|!ri��R�R�z��OF���O��$�OТ}b�'�X(�#P'yF�1'�L��k�������I۟ �?�'"`<�G1:�I�w��	�LE���?����?��D�)�M�O����B�I�3vn����@�Hph� S'�x��K>I/O��$�Ox���Ol���O���U��,$�mɁ�o�a�B�<�TW����ڟ �Iu��4S~%$���>%�	F�I�k�`Q�+Oz�$�O��O1��� b�7l$�M�<�d���2n��`)㗟��a!�0e����M��qyb�Wr�A�#�gm�W��'���'��'B�����O�`Bd�ȥV��$��(Ġz]
I�w��O��-��Ry�'�?O�dҀ�^B��Δ�SMȭ�3	�
%���<!�N�"����@�S��[��@�g�B1:���U�~��������I�4�	�\�I��F��ݍ$���w �q�b��tb��?q���?i^�|��ӟ@��k̓[T�b�*_[:��0�x��&����ߟ��I�Gp�o\~��m�$�'I�<z"�K5��x�k1@ӟ�C��|]��S�l���pc�Q�8F���`�%������I}y�>��?�����i�0%j�ه��s���as.ؘU��Ieyr�'^�O�'�e
5J2�U��O�j�-����J�нCrGP5h��ʓ�׮�O�E�K>G��,�VhpcC�Cx)Hd$���?a��?����?�K~+Oz��ɠ] >}WZ)f:)�|�$�<Y����'��ן��s�ِ���Qp!�����"Ee�ş,�I(~@*�lo~�d�nkP�~
��:H�bA�PDg����&
����'X"�'���'���'��3� r�3�%�82_tqbvk�'��ً��>���?	���'�?���y��,��%�B�b���Y�]4�?������'7��X�4�~↗�_�x׫V�] $�p�l�?���~�b��i��~yb�'&�eZ-q�0L{��Ɩ>��(u�\"s.r�'"b�'�"����O��D�O����$��z��Eo��r���¤(�	Uy�'��|��,x�j�)]4o1Pd1A��|��ɧt��)Ф�G�wM*��|����O�T��'��i{�̆T-Tx��G���Tq���?I��?)��h���ɚUT��Y1&ܑx�̂2
3V���CS}W�$��F��yB���X��ᛆF/��Y���?����?���sX��ڴ���J#w�ؤY����k�OQ>�L3�dQ<J���|�T���I����	֟��	͟ Pc�=o�Ҧ�B�4�8r�*�ny�>Q��?�����?�F�F� MB k����ũ��_����O��2��I]M��X�ÔU�F�&��dMrQV�%[T\˓{�&5qq��OxQ9M>i)OL�j Ê�	2�X��͙��x�Ä�Ox���O��d�OZ�$�<qX���	H�n� �j1�`&��D��ɟ��?Y(O�5?Q��p�b�K�)��cq�OZ�Xl�Y~r�E8?qB���:T�O�#s������ƩF膤��*F3"P��'w��'�B�'���S}"�p`A�/s,���m�/
����O��S}"T����v�xBJ}Aᇿd(ԕ���q%�$�����$�	;O�ln�a~� ��RP$�hvaP���ͳ�&%�&�r�n�̟L�Q�|�^�b>�I�s�LL� ��]�=+!/X
h�0��OD��O��9��%��E�Q���a),� �TBy�[��I�0���Oâ@d�֟z���̑�'֬�6l�>Jm���Ϋ�����B���?�`�OHȡ�o�V(&Az�c��5���O>�$�O��D�O.��P�-\r.E��HP�R:)\ă䮙��?q���?9����?�+O��ĝ����	<��2c�� /�2���O�({C!a���Ӻc􉞔�bc�1ʃ���a��vΜ�h��9��F���ȕ'/r�'���'�b�'��ӏ8:=�s�B"N;hpu)��jD�'r�'$����'7�7Oh��B�ȫ=$�	�o:�J��D�'D�|B�����2כ&�O�ewG�A}xq�F8J�^=��'u�Y�A֟���|�V�D��ܟ��r+�F���N�#�6�S�k�͟L�I��x��my�e�>����?��
�X1A炠 оTA���Eh�K>����O�$$�� ���S�B��ۆ"R�g��ʓ �}��h��M+���T��?1�'���& λ%u�!�p	$fB@U����?���?���h��I%�t�{!-�	��B��P[���O�(�'���'wr�|R�'i�M�ih��C��5=n�[D� :T��'���'1�K�i��iݡZ���?͙��;a�� � ӣiz�xB�Ϡc0�'�I̟��Iӟ�������I�� d��@ΊQI� @<~K�x�'I^��?���?aH~���C�N)���͠\/P �stz��/Or�$�OʓO1��tbRǆT%(�X�䍌Pil�qS��52 (���<��F�o���������"`X����%�� C�vF��$�Of�D�O����O<ʓ��Iԟt�UI�~��!��ڙ7�P�j  Iҟ��	P�П��'��'@��B�����
+@�a��I�|�ði���$$eS$�Oir�'?%�;?4�R)��T�А��� ��H���d��؟��	���^�O���i��/����2�0@\�����?���
��������ܟD�<��+ @�@@�����5�Lq�6��T�ʟ���֟����B���'Zd)��@s-.�Pj�/>�1f�J$C�0����'G�i>��I͟����6@�i��� DG}(��Do$��Iݟx�'t���?����?�ɟ�� �'L��w�:#���S���'c��'ɧ�$;�pJ%�͒d;)�j�+OJ@bMQ6"�,f����S l@�̊C�I���`�T@R�RV�����^8D�	ß��	֟��	H�ByҦ�Oy�%M�Wl�t �#��U)�'���'&��d�<	��H�j�І$_Ȥ0H�'��jW����?�!��M��O�!i 'v��D�S�7����@�:y~P��ӸM�F�d�<����?���?����?qΟ�[�#t���[�H��I�<}�j�>���?�����<����y2�[ƒl� ��;����s!L�?�������'7}h,q�4�~Ҡ�IȘ��_��t��o�?I��	d}8��O����4�����?F��L�U�D�1�HY�5&ʣ-$h�D�O����Oʓ�����	�DI�.܊9��(�GСIRU����l���d�O���1�d�<|�,�7p ��ru+$'�˓ܨ�F��7D0�(���� Q=OhU)��=&ޤ�,D��0�'b�'�b�'�>e͓o`�����|i�G �*E����$�O����O��hΓc]��:�j�ԅ�(M
���s(U������	� �z�o�n~�J	2u��O��y�� �dD9�� ��9O�1#K>�,O��D�O>��OJ���OJ� �]G�"F��iY �Վqab�T���O���O>�$7�)�OrtHHISx
�%�ύL6�d:6��<)��?�J>�|�$��z2тQ��
Q*�zŕ;l",kٴ���@�|���'1�'?�	�S�6l��F��(M�2��!v�`�	�������	ܟ̗'��ꓹy�%�1J��_�l"�.��?����'�����I�<93���־�JDC(������$o��n�L~r*�>�@E�0�r�
�n�oN�� B�C�o��aٲ�'�r�'���'B"�'>����k�⑐G��- �4��U
�O����O�d�'���'���OI{ � �>2�v��ց�#��'���'��'�u������Io��
R� �v�n���H�"Z��en�/!q pR��G	}�>�U8X򾭲҆ {�T�p�j�K!�Q#�l�%5Yإ+�Q2Rİ��3W�E��M�kΚ��JU.��҆
\/Y}��&-
�eZ�d�%��%{��%2�H��\z��Y$}�����(�3=2�h����;sOn��-�5w� ��Х�����7e��K�*�v�T�i�ȪP��1ggęSe�T1IW�����N�[^6�p�ʒ$o��r��Ǧa�6��&�=�9�Y+}?"�z�E�wf0Rȗ.{:�����B1	�15Ԝ�z^<�q3r
I�x�(��`�xM�2)��
�XT"	�g�9K*���#ꉓA��T��Dհ>����� @�f���N����㇝�S�L�,%(��DO�g��X�Ԗz_�0`�	I5A�����Fɏ2 `)9��	|��$����x�LH��ix� 6L?U��8@A&�.��ge�*@��;F��R:�D��j��B"�a���i�0��eL���J�`��Y{Ǐ�F��@@I�,y7��U&"L�1 ��9�ď1BA���D9|�&h����O����O@	�'@���pAT$��e�G� �69H��'��'���'Y�'��(U��Y@4͕�|����� @���1�Jޟ��I�M[��?���?)7Z���'���V��NYH����5t�e��'��$��'_�'&�S)e�*����ibҐ'﶐06CO��֠I�I
�M���?a��?	�\���'i"<Oʬqui\����&AY�<vt��K�0��o��D�O����O,E�%�l`"�5��@��OR���O^<�'��͟0$��r��B�mt΁8�n�	qg�D�s)�Qy��Q�>$�b�y��'���'��S)o�D=� ���%p$��1'ԻG�T�DC}rQ���IR�	蟨�	nkD��(H72ז����p� � �DP���؄�v�p����0�	w�S��MG��"�	���H���ȟ4�')�|r�'(b��:["��('�萋�.ϐW9@��U�r��}��'��'�r��m�~�j*��jT��3|Jf�Idc߬1����?�N>����?�	\Ř'�b�kQɔ�nM������(|�;��?���@�Beϓ�?)fY?�	ԟ��I�nչ���"
��!Ǌ��'����ʟ H�N�\���t
�����YF, |�1j��*�?IFa�<��I��f�'���'��ſ>A��[:8�t��uJD�oO|��	��?����?�$�o�'��!,���L������קs��XP�N�ϟ���Ms��?���?QtS�\�'E"q��a_��������M��'��@r��d�|2n�<	�#��i�׆%�Ҝ��m۔B6��Ըi]��'rR�'V����O��I9$l 9�*J�(����`nM�N��⟜�A؟$���j���Iӟ��\e,��,%d�a;F�:8�L������	��S�4�|bK�T��y�� ��60r4�+(�' r(ɔ�y��'"B�'y��?�I!������K1�d��FT�	ן���M�IWyR��a��u�ݡ{��)Z6��#f���'5 �A�O��'�B,O��SCp6��5�	$�x����[ws��$�O���/�Iҟ�'&t�y`
S��%�u/ʪFV4�[�e�\��Ob�d�O����<(����1v�T�QA��!��!QD��&(��d=������'7n�YL� S�"J�4��"Ōg��İc��O��O�1��<�-�����O��݉?{t)P�"X�YzF b'��9WJ�OD��<)R��t�'�����)֢<������Д0�`Ѫ5�'a��1D_���I������d�Iy�̜y�fŢTޙi�t�8�
>3"�'���U�#<�'f�1��F	���ђȍ�_"��͗����O
�D�O0���O,�S���xD�K]�kZҬB��F�	o剓
*P"<ͧR���͓�?�����(?d|�s�E4�Θ�'��YI�6�'r��'��E)�?e͓1L�x�g�O�&kX O�t��̟�$���I�i ��?��w�*pZ��;lܔ��MI45~u����?�����|ډ�bӌ~JdIk��4>@A���#�'���@���y��'��'J��l(����9�F��)Df��[B��ϟ��Iw�Oy�-
f7�%�V�E��Ic� P���'w�)�O��$�O�i�<�O�b�JB�����e�+;L�����?)���'r]�,*�L��!"���
5СI$ ��3J���Mu���I˟���V� ��I�O�у��o�nUaD�Ŷ���jD��O ��6���<�'�?�ʟ�ꚨqR\�!��fv��D�'�2�'��-��'E��~���?)�w����PJ�<ݮ%�v*׹D�:$S)O��Ļ<I���?�J~Γ#T��e��}���pG N�y�(��/�X���?������'���'��T8�x�Y�d�%�۾+��æ�O���?����'��Iޕc��� ���DHAf�����,��8�`H��'�rg|�>���O����O>�'����@��y�G퓻D��ұ�ܶe2����Ob��OʓO�I��b���O����\�c����oPD[�����A�������\�Oʓ�?!�'Մ�J��,J<xDpv��D�~�A+O*�e����K^t4ͧ�?���?A�C �VU�נ9y���熠�?	���?Q�Y���'��Q��̻yع`v�
/�"�8��'j�D��'[`��'bV���'��'���y��I*t4�䂅)^� �k#hĪLW�>a(Ol��<i���?���-ެ9#��V3	I�͂ᕷF*(�A,�<Qg�<���?����n��T(����(�t�^\T� �gi�?�)O���<���?��~�<���}�0'Â[���C�$�g#������?q��?����(�@$�O,�Δ���ɻeLց���g,U�[��'�����I� ��h`��O�� �gb�'0�d��Z�҅��'��'��1Z�'���~��?I�T E+S���7^����g�rTQ/O|�d�O��Н%��D�OB˓��DOF�e�b��
ץ����ׯ�?���<���&�'=b�'Vb-�>�!�E�'�y�ޢ�5�p���?1���?I�g��<aO>�)�(4����H���j�.�j �UK�>t�D�O�]m�ǟD��Ο�����D�<Yr��6^zAz�*_�>�P$c�N��?1�˂s~�Z���O��\��O"҉��8���3GH���U7��6��O6�D�O"�$ Q}2Q�����<Ib��$m�b�G*I 
�+֨��L�	ay�Ȍ��yҦ�����'�=��9K5��L�^1����/|�`�W�'���'�����D�O4��y��6Z��E�$?G��9��Ҏ�?��?4hΓH��ϓ�?I��?y+� �3v���(O�q�G�-b����O(��'�����'�R�'�R�L�q"9�"Ċ$f����	Ñ��	�'�R�9�'���'8r��� ��B�{N ��1`T7`�Q�',�؟��'-��'cҁ��y�"I�v,���Ț1�dZ��G��l9���'�"�'!B�O.哅����O^�)�(\�gJ���Ǜ0T�dtH�(�O �Ķ<���?	�`)28�'�$���}�QD�)26r�b�S�d1��'r��ؖ�y��'H��'�?���?����$���S�Qm�)r�d�����OD���O:�11����'���I�*p6�P�hK0�<�@T�)Li�ܷ�y��'s�6��O���O��dT}�ș�$�6�4%��#s�
(@�FB��'Rb�Y=�O�ʧ^12�Z�
ҪQp�����2P{�#߼�?1���V�'n"�'��/5�ɩM�̑`P�1G�������ɠd����	o�II�D�]��y�'1r<��.�y������2&���DCg�z�$�Ox���O���>9���yR≋�t��#�΋nnx���ͻ�?1I>�pd�<і���<����?����@��
k��i��[�Y�QC��?���j�'�r�'��'�(���&W��l���@�>e�|!pS�<s�f�0	r���������l�t H�q4&I�AG�{�)���?�p���O�O����O�T�ǈϮMJڼ"�
:l=NXQLA�=���MV�D�O���Oܒ������9=ą!��A#�Z��C�4�ؓO��d"���O��Ӫ�������<��l8nb�9u�R Z��} �2O��d�O~��&�)K[�T�'x��ۇ'ڑ?]��r抏X���j0�'|"�'R�I�Q�����v�G�	��H��˳-b�ͱ�H�O\��OB� �9O^���H��'���',H�86�L�4��f�@�6<td�0�|r�'=b�~�"�|"1�j8��\�1t��R�$�5^P,��'U0��'J�ne�Z���O��D�O*��'��B�R��Ȼ+V�}P�����?��Z>H|������IX:VO���PB��7ٚ�r�mޏS�&x����Ox�$�����ğ�	ןĩM<1����Y�1ò�c�����
�O��H�%�O��O�˧!�1��?ه����t�2��4L|��d٨���'^��'��1�$�O:�Dy�4���F�6�d�Hr�K�4�����Ob�O.��r5O����5O��D�O���3)��i�m->Y�Q)"�$���O��P�����}�0{�pĊdD�2���Je(�8h�'�L(��'��[�'���'���?�S5+@"jx T�.�e�D�!��O�)&�(��՟�'�,��՟\��`
��z���n�ujᣚ]�,��8n�	ꟸ�	�� &?Y���E%Dpt��AI��,
8��<���hO>ʓ�?�R,NrtG!�8����!=:�Γ�?����?!L~��[?1�I9/X4A%4_�dYQB�G�_!��	˟�'r�'-�`���y��'e��T�܌$�W����ǀer�'B���y��'4�ꧯ?i���?aḟc�x�8��P�o�	�2�L5����Ot�D�Od-�є��'M�S?`���vk�=��h0��ɦp7�I֡�y��'I�6��O*���O��$�S}�i^1/��3V�d�@��i@�4��'�^����<),��1����DY3�ؓ&cp��4HN�A�b�d�O0mZ���	̟��ɾ��D�<��(��#��e#g�ς6��#�JW/�?i7��<QK>!*�$]��3O���Z�����kp�J6���l��p�	����	����<����y2�G4|�0��I�(*&Z��H�?q����DǴ]���`��	�O,�$�O�� N�;Eˇ���:��-`����'���'x.듰��O���y��]�kd�1��c-�d-8@-B���!]\��
wf����O��$�O�9O�5)� ?�$�*5��+���"�O��'��	���'�2�'�R�F).����&��)q��x0%bE�J�T<�'E�d�P�'G�'��[>�	�ܓ��0cC��C�ꆹZ�R9�v���$������g����'H���샎0F��u�\�i}N4B�+��kz�S�'B�'�B��T��~*�R%2�U,g�d��C�ƕ(�$�����?�N>����OdM��|�$Q��	��al�pc�'�2�'a����'��f�~���?i�H�6�8��PO�|��A�/��qN>��0=��['��� iEsWP��C��B��s� �	��M3���?���?a"W�XH`D;>P�2��t�4���OD�$�Oqy��Q�4$�"@�Y��M2Gr���pg�5W�����'�hx�`�d�O\���O� '���I-9 D���5G�^,S�n�1����ɥ2�#<�*�hT�@1O����1X ) �	�ZcT�����<�����O���?a/O�ʓ�?�'����T ��h]��4L٢0�|#�G`�'[�TF�=�yr�'N��'��pQŹG9t]�!��7AX�L�0�'!��'��OHʧ�?�*OJ�!���,��p�-�)t����"�<��h��<ՁP�<����?A���B�OV���g`J�!R�<�dA�6,\!P����d�O��d�O�O��Di�0��%��}���	�`��\s���c��O��!0Ć'_����O����O���^=�@�@y8S@�(�OG(&T��?���䓰?��#q.���gi~ų�O~�$pTh�r��a	h���IΟ|�	G�S�����O��Z��xtΙ�p@��>:�('��O���>���O����(`gqO��i'�9Ea�E3g�W*��$��'B�'x�X�'����~����?	�e��14�R�G��y��	�AД�H>����?���^���TbW�|���lQ�jRE��$�?9Γ�<���4H�v�'"�'�i�<�%=@�I�$ݚc�A��I�ğ��I۟t��5��򩝠W�aȄƀ��(��F0<�@�	�O����O����O&���On�����s�$٠HNs�zlatM_�r�^ʓF�2�Ex�O�H�A�'RC��0*
-"%����O�n��6m�OD�$�O~�d�Z�	I��'Z��Ȅ��3T�}r��#$E�(`�$D����Nx���O���Oy�!��h/��9�$_�`,����O����O�˓����O��O�y���Ap�Y��Õ�1n�:�.�$JN�H�Q���w�ˎ*t4Y�G�	�<�ءB�Ǫ,Ę�"��
,p�+D�#�X�:ҁN<\5v'a��?I��?�����&����!$C��:�{v��x?��P��M��y���'R�'�'��	`�,�#��>�85�p,�/1�@̠�H?\�t�A�V��
)�b��t�|!c�"�H�J�.�%%�l�GM7v��R�9ㆰƈKU�,!�n�.{ը̣��0w�Д�4H=b�^9��7��P�G�NA�|��Z�z�Ǩ�ar:82��G�X���ؗ,�k�����$�,YL��	�w�
9PF��uZj���L�t�(�*�_ET�R�"j,�*�%4a�j���� !/o��Baעhl�s�(�c}$@2(~^��5 ܣM�ؼ�%`AR��9�b*��H���:�E�yh�Q4��%��̟T��gy��'"R;�X�oR8c��їM)������z�m�4m�n��(wx�,�w#�Z�Rl�!�̦DY�T��g�|�24�H?��+#]Ax��*4�lӎ@Q �	.�tH�fG܄Yɦ ��؟4D{��	0 {�9���+�ƬQ���5��C�ɾa�FM�7�_�0��h޺.kz�'ABꓢ�Y�s{���'qr�i�  ��K�4Av�9��Z�DTVq#Eɣ<Q���?Y�P�0�!�@"�� ��\�R�Zw�@�7Sje��E�Df��(����:�8 ���
�ΐ{``�?A�2�װK(�Eq��@85����.�"����	��X$>1 hX�3�b1ϛ�]a y�k0}��'� ��$U ^GZ�[�H��Tg�X��P)�� 	�~��I��{F��� c^�na�'e�9`�k�>����䧨?�ܴo��
�]g�4I'���\���'p�Ѕ�ދd�@q�bv}*�f�8:Pa�9p��#�5}_��#P�����CV�vq�����0|2�/�Q?�5�2	:i��QW�\F}���?�������4S�dj��_�~��E97	˅[��A� #D����%�?M���r�˦�F��0�	Ш��u��-"5 �e��s����R�O(��O�����M��U����PyB�i��	Di�Pj0C�n�	rᔌCS������9O2�(
V�R�3�	�.�8����
�b�piÑn���q��>�-Y|u��ǒ��}®A0l8��j�vܞ��o��~�0︡�I�,D{��'�Y)U��h���j����wt��ȓs��@�H�|��P�R/�}�L��:ő��'��L3��T90��&��mc6�Z8^�xQWH��1������	kyr�'��8�&5J�iP@�EG;`�*\R!��U������xmڱ'��s���yK0t�ã�!���$A�cK�� �i�$ꁰ��x��*)���X�KDH<y&�d�֐AW%#��p�e%^q�<�WeΑy)�����'�b�`uL�b�$�`�=^��#�i���'�f�U%T &�x%�K�+�*�1���	8�~��?���?y%���?��yZw��RS�`:�pR��Z?*r����DX�t!�>ӳ�A3@���CN�Y�2�2�c �6	���[�P�, c���
C��<����'�R��ȓj/T��2�X��L�A�޲` �i���7�~bf��e�� ��n� C����X���	�Q�Sݴ�?�����?q۴3�tqЀ��;t�t4�wF��Xؑ:s�'ȸ:t�I;\	��O�Y�S	b���a�,1���W.�;5f�LqV�qo%��S�O�B3��6(	�QI�d�D����O�EIp�'���' ��S���p��Ϩ^+�(9č3K�:�'���'2��r!':oHXYf�߉[l��@��$�W�O������ u�V�АɑFl�0��OT���O~dڔ ������,��Ky�iY�I�g�2Oz����HM_Ɣ
O<i���H؞�3p�B�r'�=y���g�n4am:��=�a{B���zm�׬�u=B�P�ȋ��&�z��ISX���&+��M��
�e�U�P���6D�����??�y���O*q�7���l����X9���tH�9�jyX���4�f��g�K��M����?�������O��n>�J�y�LM� �ʅ�9\�����$�a�����M� >K�b���W[.����Ey؟���a�쉚V��)wd��@�Ô�M>N�cc��kH<I�jô ��g@׉,�8����v�<�g�S�o��8��� {b�"�
�v���X�[���b#�ip�'ߛV��0T+:=�Nܙsu���	��g�˓�?I��?�G�ؑ�?A�yZw���2h]�W��M�����4bl���d��w��>5�ץ!b�鶪ڦ��z�	:�-����v�~*N!h䋁�+�d8k�Μ�[w��ȓY��țS-ҷ[<
좑i�4������~"D�%R���\�Iʞ����,b T1޴�?����'�?�ߴC�҉H��A	���F� �I:4�'��H���'`1O�3�$Y�zVn�;'����
�a�aܲ"'�	�c>#<E�@]��~�c�^2DsPHd�����3�r��M��y�^�H��Q8��K4�B��,8���v�J!Zk�U��(]I��>y�SF0�E͛�p������ZX�C䉾\4ls�JQ�{t>Tr�ŝ�CӦC��9xlz���j���+sʡ�7FF�xf��IQ��O����q���C9xq�͜%*{D] P�;D��:�O�.D9�!�<r<�i�D9D���M�Rl�$�p�U�����7D�d c��,T�����*��DE��2A)D�@Rs�۩=�X@ ���z�tep�'D��e��.0VQ ��J*u�8��6D����݅]��(�&�"��J5D��+��C�|�f]��&��R�qu�3D��#�"OT�qt���D�ǃ0D�ðț�X��J4�Z$�T
@b/D�Xk6��P\0ʇ>p���!&1D�IF�K�_V�`�dÛ,A�V�+'C:D�l���
��4m���b�Q��;D���5�:e�:�w��Hv� �#D��4i�4��Ed��6�V<��'D�$�$�=�Q��,.�ĚE�%D��1+Gt�⡈��������a'D�Xr�"\,[�@ԀEcBW��pl$D� St�%��U����V�ɉ!�D�i�~��%IE=l�0����!�d	PzeR'��Is����E�O�!�$I�m],�KM,	o`�l�ݏFe!�$��&��}#�O��y���2sG�?�!�Z{��p����0��[�E�}h!��  X'm)
c�Xŋ�X��S "O<�YV득~,�)�����3"O�ɢ�&�ihv�8.�Zo&�h�*O���� D�VӼ\�A'N�<cj]�'�J�9�� )/�A*�'F	1C̩��'�T՛���hmR��$��<:*�b�'��	Q�#N$Q��ptL��8�(�'�`Qf�$����&��C]J
�'?����͙�4�q	v���8��'zLPp���*"�̛%O�)�:R�'��!O�� �őt��j�|Uz�'7nQx�c�RЙ;�� |� �z�'�j�P�(X�*�0���I��,$�R�'g@!(W�V�K"L�����9q$ҁ��'��9����#���G���;�8�`�'0$)�1ԁU��ZټL^��''��2W�'5'\�BՈ�:^U�5�'�����~��DO�(�@�ȓ_ʴ-�q�[�~���X��r^��ȓ`�X1�G��-=���I�
vo����4%�]�g��<9i�ݩw�Z�"����ȓjJ��d��w���rB�S}�d��U��m#����<�´��:�مȓi�ޱPƍ�,���2wE�v'H��5�yv�ǔ���G�ۉ�$��+���&�#!��s�*UPT���ȓ6j��t�3@�*u��'�W�m��3�)
c+F!t���gVQv�,�ȓ\[�	�G��9L�J��e�R�GU�<I�&�d]p��qC��K��<�6 �U�<ѲC�c\-�Vʘ:,���)�K�<���R�w�\���F�b49x�_�<I��ܤ�p(2�
������Y�<�$��#�r�����a.��t��T�<1R�"H��#�X�ZN�:�\�<����Ji�u#��G�2[$(c�dZ�<��f� �*��t����:`Xs�<�%�D{��!W�ĬIe�Ā��Ei�<�!�}V�<3�n�+`G�<����k�<Fg�'$"��w� &^�I��ٟdsR��qO?aׯ�
pS`�r�&.�8�z�E�S�<هK
���x��! ��*E��W?	�gY��v4LOF�B񤞄@�xZؔ�f�K��'a�E��ƻf�N�Z���\	���5�
+
j����S����ē�Ќ��f�%uOx�R��Ť7_���>y��b�(DjcJ��g��5��4�vD���ģ:eV�#a��y�k��DwT���S�?��d�$��i�,x��;4��-Ɵ����Y�<j��B�N��xq"�
%a��\���/lOP�L��۱3;��E��!$5^}��9��+��^�H<��#�$�� �'����tԉ,NL�`2𠈑�{��zU�ز�]��2a��l�iA���U�n��T�1����瀌,G�U��J�IG!�dš:��	9񎏚d���q��Вn�X ��-�?A�/�G.9�)#?��-y�Nϛe���a\SI�aλV�VrreO�P�b@%�
=J|����P�r!�W83�L�Ч�̤tΐдb�%k�v�K��~��t�'LO(�Q���W90�X��'J̥���]�Tk3��,V�=�`jؖM�,�kG�&�jo�`�� 
2eB%�r)�z����t��#ѯG�^���ς�n��1Q':�lԃA�u�<�,��5Eb	�&���;Ћ�),��h���!�y�.���l����K�S��(B�Tf��CT�WR�27&#M�"��$��'+*Mi@��8\ܨC�j��J�0�s
�/�Y����h��l���2QTR%�Ra��q��JM����2)�m�`�5j��Hx`
�RR\ϻk�ά����& �јf��j�^M���5P�2l��&$0ꔅI"`�yjh�k��W��E�N�'�h ��%�^bu��%4����`H{�i�<yV�T.d���a�h��x��o�r�'�@��ET�:k �C��ݎ?��	��Sb�m30F^�I��x�A�\z�-#ƛ7 d��ʤ+M����g�3��O`�E��b�`�H13�`��>O�H�f�4T1�<S�耴i�d��O�B�(2,�#Ҽ�˥��V�? �ѫ�̈́�^F,���hZxd�5��?	�H��ɷg
xh�2$B%VnA�T�]w��TC���O \J��5L0� '	ȵch@��C'Wd]�4c� q���˒�<P�A'�kL� +��D�~�oQ�-N4:��'T�h�ڔ�]�8�H��A�"�L"e�F�O�ȍ�sOT�`H�	NA%Q�d��L?�|^B�BEDW�Az��� N�c��G~"�*#�.��ǔu^9�O��4SG��J�ڀ%B�K����i3tת}��,@ ].��D�-�џ,��j^g�xlQ�N�	�(����)�d\	�"����)�	� ���@�#��y��cE�"#��c`o�<N&�3�	�&>TB�	wN�h�,��Iv�3EGC�R�ba���Z�!�
��6���	�S�f�]�z f��BL�%IX���7�Y�2C�ɧ<���b�	�j%�-!�e ��t��J/3� ��v�>E��'�&9�� Ю��DR��� b<�=K�'.��y�E��(|��M�Z^�-3�'Z���� Ô�ּ��ɉ��X1pd�.��u�𫉷�D���\G�Yh���Mk�"��W�6���,p|��`#D�<�ב^ɚ1b `��K�ި�s.<�tz��Ĥ�- ���|*�NT3Q��!���Q����dCs�<9#GS�!������rX�tk#,�2v8�I�!;H��ҧ���� p����F�*
�t���MC=�!�D߫ ��)5�H,�t�
U�,��D�P���� ���p=�SJՔ���:�AI�f%B����Mt8���#�5��n�c�~��2A4�uH�� ��C�	8?r|д&�& �I�pI��ud�"=)�E;<�}���T�K}�����,i��q2�I�'O�2oYi�O-����2�"�%�$@t���'����EC����`k��uP�mhsKI�[1�3H>a���OZ���σC�L"	��H�2�*T"O��`*�|ꭉ��ψ
��m�X/� �"%�ym���1��4�%eۧ��yræ�@]����	7MhȜ(����`�b��D��uX"m�:g6	�a�����dZ<{w�d
ד*'V,8���C_���`M߇Me4��>����f��`�4��C�0�@�BK�����~l�p����sBB�	I��C'ܥn}��"#ĳU9�����>s�U�Ot�KA	��wq⌳L�쀟w��� �i�1V!�l�,X�A�'$���*��z*��3��-��p����a���H��ē2N퓒τ�{��Ov���dA4"��*�0,u�����'�h�P&�O�Z����</��T����aH	�1+N�%���F[n�h���Zt���V�Kv01 ��'ᠩ�� �/k�Oj8��!�Y�$�I��H���2�6)p�ě����hd,�	uZh,ۀ�)M���5>h�у��w7 0�j$��� C��<�'�@��!�h:p�%>��;C&ht{Ɗ@�H����8[�`0�ȓ/��� E�}r)�r���aq:�l>�Hc5��/g_�Ӻ� ��p���&�Ǉ���R�_5Cw������y��۲f}�Y�qe��V{`��a�\k�)�ɥR�R��֩�Ƚ𩟑��CE�9�t���4��&�"�O��(v B8V�t4@奖�~�h����-#  )���V[`���� �O�ib4�ٴ0PwD�aw��h���:~�Yk�cG�/
�9q�X��)�8��-���'H@;�l���Py&D�n�8X�g�2D1r����+�M���@����b��F�S���@eN,���rFe��]2t�wh��,������8D��9B+�J�ǈ��P)����LU�&����)�t�l�X5"(J�L�g�'��b�銺h�.M��W'Z��l ӓh��dh��S,UV. "��	m�d1	�g.f�#!b-$��%��א&u��	�Zy��L�lT���-Q�~7�%����&|2聡!T�.��9���
9�a�/���U�q��L�r�ό�Ԓ�"O�a#�Q�T��abQ�(�D��'���5)�%�0�؂��~��>E�vj���yG�ݱ~\q0���e�4�h�,ظΐxR,�/.`I�Ql*.W,�8� W�^7N��W6�ֹ�҅��b]�+$taG{R�w+nTHz$c 
TH �u��ذ<���F�� �Ԡ����K�}�Q#��:0�D�#u�-�n���4#pa~Bh�;_f�*'L�&FU�)�U�K$��L��03v+הN��Q�C�Y�a���
���S s@�+�H�%ZD8�)��<X�C䉂. ���M�:;n�b@��*wư�2G�� �����(6R�"��:�3�$��mͦ9����H���E'�6�!�$[r�? J<��S(5�|1� �{Ja�b�!z*����p>�V�T�NX��PfG�<fE����i�KX�<a�N7z˄�C��V?qw HY �ċ��̸:��ԑ@�E�<�sm��V�@���;��� �AF�;���(��A�?֑?�b���i���{��؊M�`��3J/D�p`,U�5Lz���B�m ���'<���-����&>�X���a��&q��aC�ƶ}^��ȓg�����V��Թ��f�u��l#l�JaN	-/��@I�W)��%�ȓF�� �!���^�x9��ˈ,�~���1� (K���d��ظ@g3	���ȓ0r�8��9<�^�@��H�Q����#R爭h7�8�Ȗ^�t�ȓA�h[޻E�>�rA�մ&�\,�� 'x#sFZ%��Qb�-̳]J�=��L�8ܨ�m��q,�1
Ƣ�>�U��%�rt�HE�xY�I� +�.\�ȓm�6�ړ�`hpL��Xu���� $,s�]�A@��Ѵ{^2��ȓ/����kU'z�X=��Iֱ@h���w-n�bѡ�t��x�f� 
ۂĆȓh��*%���jV�	��A�J�}��~�=�Ek��.�$ �%�9PՐ�ȓ�B��"
P�y�U+����[�&=��.nD������X����;���Y]b�q���	6F����֘)�ȓX�.4�(0K���҄��
#*=�ȓq>��JQN��	���0ҏS�>)���3*8�"���%��m.m&���F%����F�
L���x3���NU�1�ȓ gΝBB��)���(r��D7�ȓ!W��B��#?T����H�L܇ȓ	<��y�]���
�B,Ն�>�0"
��4@�&@�l�ȓ.֐e���A.b�6	>J-���*\�Q�C�%/rhqq�L`��h�\���[�Ҁ�oB�
0��w���a�R;�ѳ��ȥdN@�ȓ��i��٩VeN"��ݮ*l$����LBVF̟yD
�� `<B ���ȓw�������>gb��� o���r�<�2���7ެ��'e��j�p$Gm�<�fJq�0�J�(��Y���\�<��S'j3��1!�ri�y�����I� I�ƣL̽Rߓv��Z0��
2&�����)��ff���ğ\"`ƭ��i�����|�%9��Q�����Z:����g�t���L��mzj�I��[�K�D-�ȓ~���c�M�7%򹘂 3�ؐ��8�DI�B��8�`E��±a8`��ȓ\)�� �ƛ=l�v��GhA,-"�̆��xL�*ϹX�����(RYf��ȓ:{cl�� ��Ŭf�p|��gA�(�U���Atj@�DS4}	�A��}r|�cG�X����ڱc��(w긄ȓ|Nt4 5���J	b�i����U�܇��l����O�T��b�m�Խ�ȓDL�m)��	�q{�E1�,��j���ȓJ%Q�'喉�F�P��\���q�ȓn\l�rI%>�(#
G�E[� �ȓ%mh�A�V+	���p�o�h�\�ȓNx�$�敲p������Ll3������E��	��H ,��CF��ȓea��Ek
�RNFq�0
P�u�Jԇ�S�? ʙj�F�o�hIcKp]#g"O�!� I�J "ԣvfJj�j}�"O�\�GP��Z�{���%=��� ""O*x{$2X�&�2�a�(���"O�@	�D�� �e��ْZS�%��"O^+tiJ�\^�j�n��:L �8"O��)u��-!�MY�M�"q�����"O�����ުl�̰���U��	Xs"O��PQ��.\�6��2���,e�"ON �	$[s�`K7o@-L"J���"Oz��.��X�vN�1o9��]�<�w$_���Yj����=��0V�<a�C:=���`(�
P.`h��G�<�2ꇣaИ�P�K��z"`SE�<�CΏhj��1�n������K�<�E�7b�x�*�Ǖ�4�j���G�<�%	@��:�#�,�p���E�<is�*M'��`�Z�{������<���3kN�PwD�;bT��B��z�<!��	t8��j�l̴(@�:5g�w�<y��0T����%.�����Kt�<	�hÒC��E��\1��p��L�r�<a&-�m�*���4(�j<ZWj�w�<1������5��#@���x�<�OU�Z�V��!D� )��ٰx�<!Q&�"y���k��
̙��o�H�<A���-0����Oӈr5��C�~�<I��S�u�x���z͠ �Sy�<�"�G4�`���އWp���Xv�<a�-ϭ<�UG<5P>]`pn�H�<!�吺qè�Ҵ*�9-��0��L�<�Я�!>)P����/ &|\�6��@�<aa��H:S`㙢i$J�J%lW�<�v�C9"G��A����`�"��桀y�<�c�:j4���yR|:���P~��#�0>�#)G7qD4���҅z�Ir��v�����jZܟ�V �L�d�éD�`pkg:D���ը>M� I�p���J#��
����)��}$2m����:^�`�o*!�̦b�����HW�c ���'�[�h�d^��d�"~J�	
�0��ι/���rhZ�y�%�_���AG-E�>�4�J�(���[�u0���	b��`x���1.h�X�gʠ �a~�eQ�HGR�Ǭ#t���a��/��a����yr�C�tFX��H�O����i#��O*$��ӭg<� ���M�z�0Hgɾv�B�	���Q�$m�1e��Q�@B�	�-@������r�|�򈚲2��B�	�"B�C��M�����ؑ`N�B�ɀT� i�q�^�hnH�qD�2~�B�I�Q��x@
G�_���� oN�l�B�<(p
��¯ֈU$�P��!t�C�#z_�89fm�(o���J()�B�I�|�dh�@.R$@�w�G
N�����FJ���I�o��0�o�"-�8 3ӣ^0|B䉝o�UB���i*�y����vH��=9���r��Q�[�ys2$�A!Sqp�)"�"OSeC`q��	��f| �u�ij�A� �T�\�c�_�"~n�}��}+��QO�0Z��{��B䉛|�D�� H�.	J)���Y>T�ΓoB�X���
��@�-�[�'�^���d�Uk��|0����X��!F�Ɠ7ި��(��v�)�����n���8 L�yh��'W\��ǩ�p�b=3�cE�s�`�;��N��ܤ����#�<0՟�$��dM  숉sH��뚨�y
� ���&��T�,���%���	�,����K���/`nPAAv�"~�I4S�eI�hSKX�U8S�ݵ<�C�1e��!P��b] `Q"j^;p��	)b��+�	&Ebf� Ab"O� ��M�N�֝pu����،"��'n����L	�1�^B"-�0!�D-�1h[I��ZE� @h��D,��q!��F�,+�m"dt^�b�*�	�~�@�T˝&ؚ(�v��Fܧ~�b
.3�&�)� �Q�$�ȓ2��9��^������ր@��*ń�\.hd�6��!
^��Q��~�J�D�n�BQÙ�}Ha�"��?�yc�2G<�{�(C�pR6d٢��<����'�2���-�&��<�߶]Z��$�ӄO�����a8�����G�6D����a4oXq��I�Nڼ=Z�fN�=hVC�	0LvL�cf�.c��"e�56ʞ"=Q�(F��}�O�(D	W+X�@���ru�'R����'\��9��©d�iH6��Hq����'ި�yF���YR�{��W�;E���N��C��$5]��:�-CVD��TnљB3C�I�l�r������9Q�,HŠ��-�C�5V���ʗ�M�59��s��N�BΰB�ɗ=�(�2�Y%��k�kL�E��B�	fD�)�3� (
�:�J-e��C�	bL�݈�(n%�#�f�ڐ�R��Oh<�C�X9-� p�dDV�yo�1S�Z�H����d��(Za��U�T�$�;1n�@0��ȓ5G}�u ��ֱ����m�,�'/ʍ#���S�d���Eb��P[�9�A��3"7(C�I�$<��!V�yEte��L�	��c�D���M[x�8�*�eT�1����a�h�@t8�,x*�0<l�	���K�
!0� *I����ƓA���@:40������u��ȓ\�dA����V*�����I�l�:���Mt��ZC��0q"	�F Jf��ȓe9�M�ad�f� ٴ��h���ɤY`S��ٰ�M�fMǦHw��:�ℒP��{B��p�<�È���"	I�/@>��dIe�'1��d�3;z#}��gSm� 'ɔ�(�҉�f&�[�<iPa�8r�nq)@�F$��5��G��֭c���������ە'�F���̼kSL�:V+�'�!��O�~��؉�k�$��4�jחF��č�L�v�2OLq؞H!�߀o�<�ɓ�10�z�r��7�O��iV˔�C�4�l��[��!��I4' ��u#˯u�B�P*�#��	���BqΈ~X�"<C
)�tr��Ә!X�L�Ș%q|rᓭ�W�B�6�<q��?'{:�H��#��H����'��3J<E��'q� �#��+ 6�S�/@M��
�'�������7Vn��#iZ2L��`ʙ'x(8��?����� �:��!1u�ԐTP0Ȁ�( '{"�|�w��O�ß J�N���R%h!i�61LY[��5D���U��(ul�Xp|�Ո%	(D�l��&K�94�E��M�6˨�!N&D�t"�핀�ȵɌ!rl��E�<��۾X�&%�0ˈ����Հ~�<��,�W�j��S�:�;W��^�<�����K`����%�|u�3-�\�<9'��
А��̚7"�Ę0&�CW�<����(�1��ݵm�^D�K�<9�Ė�y�*�k��BH��]1VB��4k,P��h�#+��ؙqŁ#F�R"?ぃC+>yr$*R����+�@�U�����?D��*7�I�]�E� �CK�V��C�>��.]�O�>�B"�����qd����t�2D���%�Ӑ0����R�Qwg�U1��0��&�ތ��I!d�n����S,�1pJ[>x����F���(�MK�6z�e �ꅸI"\<;�IƆ��x
� ���fBs9�pɀ�U��Vt�R��Ǧ���n�%4j�����3=M±S4�u�Fa���%�!�dwUlhIԏǘ�~�1��"A�6�8�Ň�@�h�	�^�(��Y�l�KN5wb� �l�I��4lO�mc���~�"��ZY���Z�Z�&���M���T)OhT��K�&1Kaz���	B@a2���L�<\�qoZ��'_|���I@��F�G2�'<\0r BvuJ c5�0J��,ZF�<��N���"L3r@p�:@�x2�K�	�q�Z�M#����a�� ��_.{̺]�Ï	;V}�b2D��I��̶`L�LA2��+�F�h��s�
����H���>F��/.l�		�� ��G��n��0��
��$^�u�X|�@bբ<3��`!Ɛ?B�!��<'u���u�C�N&��2'�9�!�$��y�0�+VS��x���-�
F�!�d�Z��+�̍u�6p��V�!��\�v��ѸCÝ	��Y k+w�!�6�.�����n��)ɟ6�!��|�&���Ԡ|�`�AAC�G�!�$~LlPS�%C�J�s���)L�!�d3 bлP�٫=����EJ�!!���Q:�A�䋯t	z��)S$g!�$V�/�ft
�mS�Z�3��͡XX!�D�t֖�:%L<�*�#�JY~�!��(>�H�'�Wf�\�j�)�!�Djq��[i�4�k���4�!��ьk$�8YE䒷�8�z�n&�!�DD#�,yaAʱ��@�CQU:!�I�m�ޅ��ș�jw
��@�ת0!�$�%OX䉡0�>e�v8�F*��	!�yh`�u��y������̘wgPB�	��Ș�I�N0�q"�)`�:B�I�d&,�#o<�����@��PC䉟�AC��%Kʐ�1ӅӏW�*C�I�.�:x@����Zm��K^�r�C�-m�bP��� (Dta[�n]�ZuC��,p�Dzv �%��Ӣ�/��B������ۃ'�����*o��C�	 U�mb�ʟ=.�2��(�#�$C�	�b���Xl�V.A9�,�C䉔����(W��A���R���B�	6Fk�����v��m(�A�H��B�%G�Y�a�
$�X�yp�I�B�I
[��Cl�A�m��iٖ_��C�IZ$�	c悱2 ���`x�)Z�'ɪpoP T�� q����_�X��'��%�dn؏"{����ķH5�M��'7�ZOܘk��%�dEN/��!�'���Rh˟x
Z5yׯݷ!���'��D8��J6�^t�aA0b ��'�:��"��A��8k!A�o�x9�'���q�I9����h��y��T��'ѢYSA�Kܵpg�Ms�p��
�'uX�YrJ� zG�	�'�ܣ8�Q+�'�� R��e|T2�6H��P�'��u���H��1i�c�'��I��'�4�T&�7��Y�o�D��'�d-�a�L/^�X�R3N��t-	�'��Y*R+R>>Y�A3>�$Y��'�ƤK�Qr 5�G��5F�5�
�'>]�#��/�.�����,]�6��'�FQ ��#���䘪S��H��'��E���?����M@Gې��	�'� q�iC�H٘���ዸ>�.�)	�'1ZD���K�CW��*� Ǖ)p������ VD�� e������><�a�"O��G#�)p��ha�$N9&�x�"Obt��N�9E���0D"^`""O�@����Q"t C�w�(�"O�lR���K�Q��OS=P��2*O��`aW�(�×�s}Bu��'If�k�nˤ/T8U��Ț�o`0E��'{�h�wS	E�E��@͕3Y��	�'�P�����
x������'�H�a	�'���z��Cc�>��T`߮�Ν��'�m�׎Y���4I{���'�($��]t���y����>jJ���'�<)c���*zh�p���ny�$y�'���sI�Z�2�.e�,��	�'2F Y����!{ć(a�4��	�'x��CÊ0U�L��n��%��'h��/YO��0��U�l$�'��p�c�R&��(�n��&���'1� `(I5j<���C�nb��'�q������bN�\�{�'-�DzQ�X�A��}���+\�n���'��!�"ƈ*�D���OS3 �����'�ЛA� �9��ɳ�H�aD��@�'^d��+���L	V�"���'Ji�m� <��p�B�<I7iS�'@�(ۢQq�q�Q$��F��X��'�!�˃0mk4U�WhT-<����'�"�H2 M�Ln�Hw/>:/R��'����
�m	�ٶč�ϒeh�'�p���*&�&���`A����	�'r�|T���>�l(z ΍7�u�
�'���pL��R�:4q�T��C
�'t�P�W΃�B9(�a�jT*�H}��'�y9 ��O�ި.�! R�M��y�B#�Mʶ�ɠJz`��U��y�ӵ���`$g߷|ˀ�b郟�yB�����C�˪v���
�<�yR��2xU�
3�V�9�^m��˟��y�(M�V�^k�Û�fL���'�yB�M9]U�|!���4�`]PWJ�y"�W3�p�u��.�I o҇�yBI��m�@����#�إۀ�ʨ�y,�(�
M���Y��V��aP�y���t��*��̕�^�X6��&�y�����As�$���i�U�%�yr��cj�QED�(}�`��ƥ�yү I� �;!��n�4@��y"�E>�$H�Rnѿr���a���y"m�$ހ���L�n����p�M�yr�ߕ%�v��" �2]�5{��@$�y�@b{ ���&v�����yҍ� �����N�R�O�H-���]F��rMآg��%���-�ޝ��K���z3�#<���+��u��}�ȓx�m�t䙥^;���b��l����~IP�
V/ɢ)���Q�Y���ȓx ��:E���1����'�|��%��`��8G�Ǝ|�	�a�4e�	��$A��F�ܫ)dx��Ȇ6.��ȅ��XH�r�C/Zb���!�T�C�|<�ȓkv��KȦN�e��&��ȓ2r��Kp�M`�v|�&ᑈ:,t��}�t���5+t@��&�zB4q��=�`�P�"q"�R���|_lB�)� x8�ԃ�<M�.=�b���50a�''�DK�}��	6oЍPa�� �u!�Q�>j�Ȩ2\�|��5!���喁B����VT�jVX��!�d_�f��U�_T�����Ԯ�!��P����5j���!K��~�!�&I"`<� @�4R� 4/�!i!��Ֆ��փЁ_G��آ��#F!�D�#Xh�����5�(@"S�țH�!��{��P��C��D6�P��"O�E��3|Rrd� ~44X�"O8���5d��	y�Q�Yx�Y"O�ə�H��	�s �.��,�V"O���s$�
#0fCwES���a �"OV��u�G7Y�b����P�7���7"O����%�&x@rL+��V�,��X�"O�P��ÂM��8����,�`!�f"O��PG�X[r�A�A ��q�"O¡�G�@�|�Q�Q���t��p�B"O�P%g��~�`�*��$���3v"O�Ia�
�P��L��O�X�\i�A"O.���mCl,B �U8`axl�G"Ot��vA�'n����b��u&�D��"O>�DK�G���d�=jnUR�"O6���S9�$�['���>�4��"O�
�R(��!`�����E�!�$Mc�ܗ*m����׌̃l��`�'�P�3a�J�:%Zy3Fn�&o����'u�1��n&+ L���?7k�'TL�YoJ+
�Z���)���@�'K���A"h����(�h�0I[�'��!,�Jm�!�^����,D���BNY��Q��B��	�,|a�O D���`^*_�|#��F�V�Ju ��?D�82� ��\$Q*b�ɻy��q��M=D����b��,\t�#�`�����<D�4�H��3����&:��]�:D�d����&�n�*fcC�[Rl��-D��b�[�l����j�-��s%l-D�\`�y@�4����6|]<��2l,D��r�݆#��h��(~��(R�e>D�(H�O�~Δ�[3��J<�0HĦ:D�( F���E�9f|x�	-D��p��{����h	l\0Q*D����gD�r{R���OȔ_�����=D�` QJ�,��p���Ə_OؑA��;D��K��܍n`0ä���!�����7D�����~�Ju�֍n4n��ԫ"D�|zU�Y&�N)@�֦#�b�2� D�(�BG�Y �;�Ӷ}�t\��k D�(�5�xAz�AR42��:��+D�X���
�pV��� �e���0T�+D�(8�⋤1l�i����+ �����*O����oL*�}��9z'֌i�"O�!b�:@�L3&ّ[���("Or80�	����s�� ��(��"O�1��U�S�P�B���,�d=�D"O�HvY/{{p�3��)$iQa�"O��فL�
��y�� a"O�T����0��]S&׍Wӂ�j�"O0�p��F�1����ƞ�ĚI0"O��F�ق	��H��e��c���T"O�z��%& �16�_&[\���"O���M�� V	S��=�b"O� F���$��W;8z���9?�0�#r"O~��dL����ɧn݇j�t�Ҷ"O��[(��������Řq.	�"O`邒���fD������u��i"O�����v���C��rL��"O̱JB��i$�sgN%S�ą�W"O��G�"\kGX;(����"O�I����2v������=w��A"OR	�R�@��I�aȠN�\5	�"O��Q�
+�x쁢/�c{�e
"OzT�!�	p�^����\�?P`tI�"O��apdHu�#хL�Q��"O�9�K�0Vc:�s���\�t�"O�����r~<���7Vp�a
d"O�P�@���d0�E�f\a��"O*Ia���-&�� b�!���w"O��7�ߋF�!8��\).�̈0�"On�S��Rq>`ڦn�:�1K6"O��rj�d�X��lʟ18�Z$"O6P
�-�J���!��ɤ%4�	��"OZ j '�l���	�u����q"O�|4��v�J�瓔C�"Y"�"O0 S�͘ ��b6���s"O8G��]����s�M�&�8"O:�h�L�6:��aš ����"O�xK��-(��P&f��Xs�A×"O�L�w���L�`xc6NX�PUj`��"Of�ӵb�[�tA�T,�(	��0bB"O�嫥�_�������ŉ.!�!��		���8bcڷ�h�T��1"!�[0z1��ʳΐ6@ P�����B!�ٴn�BE�"j!�!`$�A�!�d]�Y&b�!�(�>	bE36���!�,4l|)��΂z��D�#cE�!�D�[�h	��-�f�ȉ����'�!�dBz���	7K�>p�phk+h�!�dώ����d�$aj�u��$A�<�!�$�z�����,�Y���N�Py"')%���h&b�)]md4c�P��y"��mVb�!E�K�I4
���啲�y���j��0*�lL?�L��Fˁ��yb���\v���%�%E B��K��y��]�]�n�r��Ik��;&&��y�žv�^=p&�JD�4����L��y�=gȵA�Kޤk*8I���&�yr�Ζq0U�`	]K�P�B���y��8����2�h�@���(3�y�ҍy��B��W
�Qr��K#�y�(I7`Y�Go�P����0�̶�y���NK$�"�a�25u(@K ,��y�JW=H�\	@��Ͼ,6���2(H�yrE8>�p訑%�2�i�qD	�y�� �o���K�OA�9�0�*+�yr��,��H�v�J�5N��g����yBѨ'�6Lk��Z���X�n�5�yB�AV�2ɂ�/]�Y���l��y2M� ``�h:�	���Ь��`V
�y�m�NJ��㫕�F�S�$��y2��?6�|b:.�aC�y�'Y2T��sC���H�*�E��y"��Z@��A��m��A���y���gy.��l�!;]H�	 �y�BT阝�B9Hք�DfĜ�yB�:I�I��Λ�G�ȕiW�D+�y
� ��S�JF�!)�Ѫa
�#�h��t"O&8C%ҭ'���{ei�O����a"O>��pA�%A� H����#@�v]`"O����]�B��I"�W�\����"O���n�=bF��!�%�#E��� t*O�2� ��K�0�*��9br=H�'i���D�V�Fw4<
r�O	i-���'����pDQʅ�˨0��+�y���*,��4�F з�f��GȚ�y�ťg�>�{���w}�x"��Q�y���@���u�ϏY8���@���ybD��n䰱�X�[�z����/�yi��g� e���(\�� ���ա�y�J0�L�� ��=<Nlh����y¦A��e%�-v��bɼ�yb��7 p�IV��(R>����yBm0
��تW�F��BQ���y��� �)�G�&����D7�y��S�7��:�*ǃ/m�sB���y"��fc�L���݆*��!"E��y��ܶ4���Q3C�,*����I��y�J�dP\-�#f]�s{p#F@ �y��
�u'��sgir�!�\��y��װ^�	eX17EJx̙�y�*�g@r�
�$C2X�
	㥋��yr-��3�X�+��[�G^|@5m��ybD� d4<�an�72�l��&Գ�y��D�� �$�R&�oc����'�n���M�6S�LPw�A����
�'�
!SR�B	?j1\	uF��'�����E�/O��Tf;�"(�ʓY��9�̀�,�*U2��P�=3"��ȓ�90��8RP�Yg �?h�N���DīG�Ղ55�|�gKX<����ȓ1(��ek7v�)�NS�_�8ل�(t��3צ"�x�I�i :m���1G�Taw�$_��5QU9ZT���x��$ڣ+t<E��I@�N��مȓ{�)["�:�He;So�'w��T��F�R=�� ��OvA�Cf�IA`M��j9�)J6�Z�\O�@E獬sk��ȓ)7����疹 �$(��A�0=<��{�:����ϩ �y���R�4q�ԇ�-[h�"�n�:#n�qc�ҟo�6�����=A�fĆT\��LO�v̈́ȓES�`c� p�> zt����D�ȓ	�@�3e⇑q������ռt38y��*C���q�Z�B@�3D�N�"	��x,-J�@��o�#�!�8���ȓeI,I�ƅ
;^��I"�ӟx�zH�ȓ2j̫��D�#<̤ao�nav��ʓ!/:q���*wY�h@�c؁GxjB䉭wr�k��"h{nl2&!�*
B䉅"�t�.֒0}�d�	 ��C�I�hK8��v�?;����$8kC��4��M�r�O$5�j]�1�Ȁp��B��-46d�3��.l��P��G�B�	�==���w�͓$� �X��W�C�IW���M+
��%Q�([��B䉜=�İZ�eBn�~�ڀ����B�Ƀ4Rr��4,�v|&�Y�� C��<X���j��'v��"B��|Q!�d�S��Tд��4pA2AA8!��O�ȴ-h�j��{�\�W��?8 !�� @�3�IO�[A�u�s�L� �0�U"O����� �vT�K��fŶ5J�"O��ɀ�6vl���i�@�<�I�"O�p��f2,f�f���w��!�"O��p5a0j?��(�?v���k@"O
�{�Ȁ�ܨ���B�J��`""Oڬ���H�%9�����PI���Ǟ>����A�g�^H*����7���@�c�/0��O~�=��|�a¯��������!'j�a4"OI�P-;4rp�K�d�6��""O�XZ�B�X y����c(=J7"Onp	��� 4Z�1�"�"O���ǁ�~�]�!f8=î�b�"O��J�,�`ؑ�e�*U�R5�V"O�qR��U��#��5��E�$"O�@����%,��m`���<����'"O 2���,���ܹ̺E8�"O
�bC@Q�J0�`m�0
�`�;�"O���1����,zQ�ú|�(7"O�Xc7ŗN`����,Ϭ+X�w"O�U*T"�>|�V|ᤋ��&D� �"O�5r��T%^���#��̣#��S5"O�89�c�(.b�(�d�X$3���J�"O()����56AZA	N�`"O���¡�?;&ERPO�~�h�c7"O�5A�[V�P���Uz���"O0�î�2)�dRP	p�ӗ"O��4�/-��SC�ݑcUzS"O�i��jĒe��%r��()�y�"O&��ä	4ݜe�1C\;I@D���"O���­�0T"Ɖ����w8,�bq"O�\�s㗑��"�F^�d��d��"O�)S���Daab+��ˊ��"OtuhC-�	������=��{"O"8'o�4z��Y��j��2d��"O��VBH�*� �����"O����� u�R��p�t����'"O~]�`�߶6 i�� ^0�1�"Oʐ����=@�u�H�)A��RE"Oȉ��.�*�*�۳u(��C��'Aw� ����$���t,= M�C�ɦʖ=��e� *`�`WM�.�C䉑�t�(�@Lly��bƻ8q���d�>YtȚk��T�2�C��\�2e��<�$�km�@�`�XEe��#��A�<q���V\���l˥e�F�S,�z�<I�	gN��2!��M����E��r�<aPh�Iz�2��Ł����nr�<т�M��y+�R�K~�1���Cj�<����>՞��RKؠ)�(D��*Vf�<YF�ΕL��p�c�^�F��Ad�<!k�.g��8�U��hS��R1H�f�<�ц��5+�U��֒p�b��W�e�<A�g_�B�<��͙=<N!I��d�<!r�Y� 5-C�!�: i�B��]�<I���\G�7�L91��dkEC�y�eV�{{�� ���$��5�s�6�y��Y�Y�vE���b|3kؚ�y��P:�̘7�P����R���>��O~��b��s���b�U�`x���"O���"��@D�����7YVp�BT"O��!�eK �
�Ӛ9,�"O&�s��%N�x���i�6���"Op5���g!�����/ `�`"O� Xq
�$��X�ThY��9R�:�aT"O!dƄD�|�&��"�"OP����	��t�[ �w����"O��`'�	��Bf%N�#���#"O-�v�8�`!H�AX;r¹�"O |��l��(�q�L�;H�4c�"O>}�GMY�~�*]��GֽZFnh�$"O�!�gG%hs��Yc�Ԉh;2��"O��7��~:r�(  �{2Z0BU"O2�g�tؚ����"|���"On��N\A\�Ȓ�`�	�E`"O4ٵ��\��@��Z����R�'��)&�HJc��\�.�ucFl@�($D��SW��dѢ}ô��o��+E� b��<�O{��ЀgOL]@�p�#�"W48$��'���@���)3͈�ە�G"V�Z�C�/�S��?�t͗�`�,-�`�ޒ]��Pj�C�<�"
R���g�*(���Lx�<��L�m�@"�S/j�r2E�Gq�<1խ05i��z��X?s�|�yᩔW�<!��Zqݺ��!�7nr��qAGR�<	�@�<o'6�p*DP��@��SR�<!�F�$��=k�!�a�x��M�<��ǄW�b]9�o[i`�����F�<�����`���TmL5��EL�<YP�
7U������}�N�U�WE�<Q��K!&Ёf�ܷx|�'EK�<! �S�W4dd2�L���Ͳ��En�<14 L3f��s����l��-i��Uj�<���Pe��0A�@)0��� �L�<!P@�/IVe+���1w�EF�<��],1Ƣ9ۗ�
�:�lZ�C�<��o�\�6��-�+"�x��!{�<��Τ(�h��j��&��9 �@x�<�G��O��"beKQ�0q�O�<�,Ŧ&�rQۇ_*i��	A@�C�<9�#R��Z�[�f���Q$�\'�y�l�=}"T@a#��-ݶ��6�Z�yb�
�u��L�d��h�Ʈ���yr'�0r�~03��OE~�8�霾�ybƀ4.�bQ !��U�hu� B���y�%PT�D�p�ۦ�qI+	�y2�Ml���w��!
Į-bpD8�y�j�m�@�X�P�@T�2F��y�k��m`����2��EZ�R��y2�	+g���@v��
��A4���yBkK�J1���������]*�y"H�5����X������y�O�����˴8͞0{���6�y��@-vb�UO�#2|���n��y�gA)yئ�SE�6j�:�������y� 
���(�hW�8�8��%I���yb��3k���n�
1`�4�L<�yR+ �sPL2|�r���y��	w��`� Ӻ�h8��T��y�,��^^(��R��ŨcK��y�j� �x	��"��<�m��� �y2��]�LY�`�G�n$��G����yBd˲����Ph/m�VT�7d׊�yƣW���ɓg��*8��I�y���:m�Dm�5�B m��aFF��y�ϓ\Hl�:(�/���2�C��yb��?�[s.�����ª�y���崡K�&�� p$���D[,�y
� �� 4*WTM Hƭ�0�$"OjU��,�N��`p�S�9g���"O�l�uo���
��Dc�?U��x"O�D��#�6zCP�;ޤ=2��"O��I���ίX&
�A�"O��(���J/:����2m
]q�"O앒`˛�<��Pxʌ���"O&]���P�	�P�q��k9v(��"O��z� .J��(U(G���e"O������8r͉i��'��pa"O
��u`�JL����[;aT���"O��hϞQ�\=Zd��
<La�"O�Y V�R�S��p���U��Z�"O����"�M(X����9����W"Of�����M�S�@ 0�5Q%"O��)ׁY������ڱy�<���"OnE!,߭
"XA!��ʒB�ؘ�yR�m��1�W�s��q��畜�y��]�H�ڱ呖]Y�\����y$�Wmf� r�>!/j]%bX��y��U��:W"!A´ӃhA��y«K�'�(��E� 1��83�B8�yb%C�*��5q�E��x�v�GP�y���<���[QZ<`z���]��yr��MǸ,k��9n�����i�<�y"J�cB��i٢�:�O��y�DˊaΤ�!��N�9�K�0�yR�+3^�ԛ��^�(lx�º�y�I�*�<��f��\X�+�E��y"�U�hR�;��ÉTҼ���+��yr�Jg��S��KlRyȣ�0�y��Y i��(���W������y�C�%! ��qĐ CI$�f �!�y�!)�ޝ��� ����+L��yr C#k��QaAB	�v��p ����yJ� �8�o��f/�aV#Ր�yƞ+����T(��1���O��yB��
.���݉!�d����ߒ�y�愋vȾ��fL	�Ⱥt&��y���2�D%�7�rt+N'�y�I?.H`�'�­���A��y�ϋ��	���o��۵ K��y�Ƌ���zP�E	���ar��"�y�4-YLq���N>��`\2�y�˟g�Z`ɗ�F�F�J��"�yrL�n4��"�B,o��0a4l��y��nv��C�eM� l��C�
��y�I��[D �0Cӆ�t��@V��y"�͙��GI������(��yX0+BuaW�J8$�p��V ��y�U�(BR�q�f��&lܨ�y�	 �3_L��dL�&a�@Q�%ϓ/�y2m�3
�HQ��	U��X�6l?�y�ê�2�1х��If�	ض'N%�y��ѷ$4��j:*~�#��yRc]/4C� sdՕ˪q#R�X��ym�,08�Cu��2��*6���y'�8lT)3q�Q�ta�qv%���y�CH:�4)RqEΏ!�Xd��a�)�yr�
Q�m��B׷�с)U��yE�6���Y��K����O͌�y��)/�j������ l�yr=n��]
W	�YC�$K@�U��y�!PI��I���S`:�ŊX��y
� LШ��4�m��F���5(f"Ol�*�@N+GT@bǦ�,u��Ӕ"O����D�4��Is�C_,,s�sV"O 0���0":P�K���[��8�"Od�kB���[�GR<ST��J"O��B�(��"��܀Q�Q�X_.\ʡ"O��`��R�2�dā�+^S��s "O}�E-އ�, S%D�p�P"OJ�Sթ"I.r����M�;�� 9�"ON��&�O @�!kUD�$5���[C"Oʀ��B�b6���碘�`�Y"Of!�Fo� m�8y��M&f��@p!"O(D)�� (6� �ύ"k�L(�"O(9�%���eX���nV�4j  �2"O�H(gI�I0\�!cV�:��ey�"O�4)�;JÌ���Ώk��U�U"O��K�OՀWҤ�@�(����A"On����Md{1C�fP1�"O�k!eʔY`��!�!��l��"O@h+�MN�b�A�5"����"O����F��d�T�`�~�<E��"O�)W�P<{A�͚��̱s"O�����	��*�M�sĹ��4�(�x�eA"�J$�B)�-1���T��M) 嘪W	���,�h4�ȓ[i���%A���Խj��|"��ȓZ�r�
��G���ԩ��U� $JՆȓI�a%N[�����21@b=��#߈�jQ%�0 T.q��O�=�,Ʉ�D=��8�`P�-�.���e�8���OZ���D��-mˢ���
���3a�?,��k�L�9��	��VT�]�դW�5�������.���ȓ|Ɖ`�l͹o�)����̈́ȓ����a["m�6���PǺ���7Z�@�f�*ʪy��NA�Aڜ��ȓS���S&�0��柖>����h,�*�PH�])&��2'nu�ȓiJ+�Bԓy$u�'5��h�ȓ+� �4-W�'X��ui
�5��-�ȓZB"��K�;W�<PG��7�y�ȓJ��9��bLy{��'�'22��ȓXɌ�;&i�:8�<��$U=/U Ą�558(t��\�k�Q�Z���ȓtBr��V �&�T�+m�5g�9�ȓJ�"�9�f�4`@�k����Bżȇ�5e�౔�å6/�m�/ה#���Ҳ�A�#Z&V��z�O5y"̇�]� �IW �|Y��*b:e뎀��a��,�K�D:�O��`�ȓR���恌.o�f����M �~A��oUb	 �G-<�!��o�6؈�ȓKV��vOȣ�XP�%F�\�$$��.�ށ��Q3����&¢yk 1�ȓy�LhB��+�Y�ӊߠ*D>��8���a�ѣ(��i�;�~��ȓ)���0��)}a�(ك��u�T���k��\9$��)Ԥ���YU�ņ���;�	� ������"����ȓd�X�"4�o����5���Ȕ��
S̙��Ib���Rɘ�.���hآ�ɕA�"(�2*N�\@��ȓT]0�"eeY/ �T���+$%����\/��!�*:.S���BW�9��S�? \a2�H�!+`�եE;/�p�"O�pK�/K#.�µ�Aō�+��BA"O�� V˝&�,�$�eb-��"O}s��E�F�,N�>��;$"O<�KV〸X����d�{��"O$����x��'�W~r�"O��Y�F��0����aE�_2d"O|�':��y�dF�MNp���"O�� ��|r�HA���0d}�`"OD��P<yD�i�㏈-�"O҉�2�N-���U�V-G����"O��%@'!�:E�0�F�#/V�@f"O�aja\�aڸj�o,4��"O���Fe�jlz�;a��P��h�"O6,!��	�����'�1D8�Ä"O������&hej�"(�&�<x�3"O�ث�⅓<��s��I��]I�"O<��&�>U��
E�Ҳ3{J%a�"O��Y���
��9b�;�|�A"O~�(R�h��e0K�;o�$�"O������p�9�gׁw^�AZU"Oz�)�`�qipA�Y'c��!)�"O�uз	�:���y[؉3a�E�o�!�צ|��8��Spd���[�Q�!�͂Iڴ�C#A�6~|0����V�!�$@�x��bs�$J[`��fb
�5�!���n|�R�^�7^ʵh�L�!��Κ้ŋ	!�G��4�!�d�rZ`�oYԜ���Q�r�!�ح/��t�a�*I_6�@��<�!򤃛�$W��(��W�X�S�b��r�~$�W�D�GW�5�ƥ�	\e�ȓ~ڜa@��0[3&���W��݅ȓ1�vI	jۯ7�:�б������i� E��OD3lv4���[�zU�ȓVV��:c�ϫ"�J�R�Bي$�r��ȓk� |�pO��c��}z�U6��$�ȓ/H
U"Ga4�����ܭh0T���o$�A�@��0f(�2�ω#����hʶ-H�R?O��%Bg�Xc�؅�B����p�W,����K:]�vB��+:������$a4ř�O�#|�pB�	 F1`eLC0�����H�;ΨC�	7Z��<ٔ��%A�B�T�G�GP�B䉫�l�)��^[D��BB�M{�C�I�)d�&e*�,R�a
�i��C�	
$t�{"CD�"\�׀�;^/@B䉶'(�y�N�A�41'ҧ'�RB䉳�0 ��^XT,��AQ}�B�ɐ<��H��҇g��]�7��&RB䉻r�t�5�ܴa�>%��&<��C��c��yzU��  �9i����b�>C���<hQ���h.R��v���PB�	R���A�ʟE�Y��bB�ɀs��h
�͙e:�0��-�C�Ir��\����	f�����.�B��*�����c�2j8���F_�^B�	�1��#@�����F�%�TB�<;p~�s�o���cs�D8&B䉠0~8e�g'/#���F�f�C��$���I�ҷ�\XA�W4=��C�	:Z�D�pa��&ߘ�x6n�>��C�I'0oPM�G�FUO�!��/��X~B�	G�~d�7JTm)�(�� ,(�|B�)� &�qDo��$E�U�c�T�wE�Tj�"O (�� �@�p�b�
9V� "OE�Lv�~\�R�V.�U	�"O�@X H�?���
ƠVE��L�0"O`�K�b�-{��R��
�$��)��',�Od��B���o���M^�I�dpQ "O� K6��'#d��+��ɞ�6	�'"O̠yhG<-�(��M�`
<i3�"O�ݳ%D�3v�!àF�hPJ Ip"O�!:D��N����MΒs�tm��"Oމ��=�JX���0�`�U"OjLQ�T:q�`X��
��OC��"O����aTlF��6��2B
;�"O�TP��E�myfL��J���;"O����D�g�d����	����5D�h�ǈ%?n2��F��4!~���2D��r���L��`�C.]�!�5��A/D��ˆ�ǁF0ԝ8����.@�s�1D����}If!��Z�M�،)Q�/D�t�U�#����3GԤ����Eo/D��[���*4�Z	 �źfuV(i�%/D�L��S޾��@�C\���Sv/D�L��l�BY��&�S��'8D��iq�&#�f䅧o�.��'4D�TC��}��Y�+��vt�x׍=D��;�E�vY�MB��45i��sg��s��ryʟ4�����;�'�� v�3&��C�!�$V�qr��X\@��Z��1�!�Ɔz�z�{����!*��G�	�{L!�ԊU�H3�R�,~��!�!�ƕO["��L�^��{�O�6Q�!����)�KÔr��Vo�9g+!��n��EJ�NN!4�(���̂l
!�D�#?A�iA��?R��l�l�g!���g�A�um�9(��hՂe3!��	��T#�/c!����(!�ы.l���X5,B��Rh	�]t!�DQm.L����ׇRF:�1-ΪAb!��nLRc��'$�QA�T;QP!���K�lA�
Б4�`b NC�]�!�� �R$��-�jal�K7_a�!�$M��I���EB ���lʦ4�!��:G���w�J�'�Q���'!�$�p�<h�J�5Rm3��ǐ!�!򤘭P�{�#�6+<չԋH
�!�$�7`�2�(�	�R�[PJA�;�!��߬/�m���ΩOxv�W�V�fL�:�S�O�x�rf'XS�"tEʩ9� 8�
�'�rLbB��s0��p��U\]X��
�'�nQ"�h�t�	� P�v�	�'�Ĉ
Ո�u�^]*�B�4Xs���'�i�� ̈́))|���gB��qb�'�<��F.�JY�až=�s�'��Y����/9%���u�X?°is�'��8�A�G�4�hH��J��R�	�'t8��$.e|���bsȋ�"OR��B�(�HSd�;T��)�"O��h�3�(!�FJ4��"O^�X��jU�P�Y�R�V%A.!�ڛ������)VD-���.!�P�7�(�y虻,6��W��i%ax��'��O��A���y��a �J�ʌ2�'��O�����7s�������U!���"O�)��j�?)%����F�?�]�U"O� <�z&�ɮ02n��1%S�I�"OT�A c?�:<k��VQJx��"O�0b���\i�]P4?JYB	�4"O�X"3�M��iaRC̿��@V�-�Ş(��ݺ�Cү=��a�+H�F|����9r�� ��Y"�,��#��3�C䉮1�htu�V�C�$`R#oܯwG�B������U�)>���i��B�ɴ|�(�:R&�>p���d��8��B�ɦ
�L����юѢ灇U��B��j��%�a��찤)��3�"<����?�AФH�R�V��v��O����7�"LO⟼�Tmr���AӠȿCGpL���<D����!� n�8�b�@UJ؂�:D�����P�{���E�< I��%D�6�کO(���#�&���3b�^�<)�(�0jcg[�h'���q�<Y�o̳{�ZIwl�;S|�2D�R�<Q3��6Q|9��3��Ҷ��Q�<!����^D8p���f��+OI�<�d_<,�48'"Lg�� (a�Nk�<�����!��!펏C�R��5iGk�<	�E�h�m�m�ʒ3'��DC�� �2�$cׁ{�Th�UG�2�B��o��[+�o�,�R�a�i�hC�9p�]
��ܮN
���e��w,2C�		��;5FK�	·e�J7�B�/�y[ǉ�.Ajޜ��=P�|C�@X*DP��]�T"
m�q��tUvC�I"?�����aڅhr�LYd� ^C�	�d��1J�W[�)Ec�)y�LC�-u���r�M��Uܩ�č�9��#<9ϓ%fpɢ��#';���*ƹ,�$��,LPG�ʘBt�av	�_ND�ȓ~�b��I��N�0EI�JR�FZцȓpM◂�9�� u"N���\��1�V@�te���� wo���jņȓvEp� ч!�x��	,�ʽ�ȓIp^�� l̇7��p"W�g4^��ȓ'0��R!�{��A:6Fšc�Gx��)Z�(�,HoT���n��\�=�p�Om�<�S��C�^4���υܔ�*&ng�<i@��*��U�[ބ:Q	~�<!Nܢ:R���G�0u;NZS��R�<�d$̼s�0y�H,*��pá�Q�<1A!��@tvm��L�G����,�N�<1��6�Tp������thr��R�<��Z�cPF0{U%�@��mPr�<��Ε/�Ⰲ��4�Z	�s�LW�<i�M�H^������a�eS�ɀj�<�OҤP�d��ƪh�jl9�#�o�<1�a��bܾ4��)��%6.HQ�
�o��$�'�H�@u�� �Ht�J\2p��+�'Z��h�
0�Z<hBe��h�1�'��p��LM=������?rs~���'�t)����8�Q)��ӱ_�@`��'[�8�aʲ0!��K��l=}3q�<D��¤�k���@�Bw��}�0�-D��s�gS�{ì����N�ڀ馅1��hO���l�� A��[ p������n{�C�IH%\<�`�I Z@5��5N@B䉁f����)�5H��T��\�4B�I�o�$M	�鄩jv��AT�[�N1�C�	.:� UX�̡MX�(�EY
��C�)�  XZ�b�j��`
��1|���"O���oM�(�)#g� D(S��Q�O�,��ukD'��)�e�zG����'��w��Q}|��%H�u:����'��0`X,J�6ii�o48=:�p�'��x)�PGw"��#@�5�J\�':R��Ԣ�Q_��#sE��,�f��	�'��B��E�)RII���	�<m+
�'6R�j�Ւwb\|/L�x��I���'ўb>�v��R����B�^�bD(�r��t���I� ��C�_/�ƍ�j�3�RC�Ɏ+��	S��C;V�q��M�Yk���d^���'�84��s�0��J���<��'��v6Yo�AB,8Aӎ؂�'��KއFXn ���UlP�����y2j���$Pq�E��(�!���_���M�)§��Ӏ>��-(7���/�
U�׫ ���HE{ʟ��*#萰_-|�+�L�75R����"O ��4�#�6�Q�N@���')�O��@��i;4d�P�O�B$�A�"O0�S�h�=)$Tݢ&
E�d�е�V"Oj���(ьx�t5٤HA8ʪ鱶"O.Q���[��}����"y�a"OL��	X)FԠ��fƷL�F�A"O8�Ra������|�~4z1"Ot"fB�	X���V��=ps�7�Ş	U�� ݏ&��+�9zx�ȓi�$�S4(
�h�r���%�XA�ȓD���[��Y_c#
6�E�ȓV  ��J�!��
"��e�	�ȓ:}B�ʓ΋+TC�8
���=�p�ȓ��{f�ԁol��I���u�x�ȓ72�
� O�$����Ń�GfՅȓ8 �P7 �>�� ¨<(�4�ȓ9b0�����0���ĊL�o��Ňȓz�tze�;P�X< W�� 7�FP�ȓ ���`�AH���a��I��l�ȓY�p
�e�.tW�y�A	N�0,�Gx��'9d����ZB��e�^� �Ρ��'�NL��%�*w�8;���%O��[�'�X�&U�"��X�3� E-<�C�'>��������M:g�a�'���� $�H�vn�/,��'�0��i��N���+�`G�.� �I�'8����/���Ҽ��cH�"82q�
�'�ʘ�W#�Lt��uDU!����	�'��Iբ��[_�يŬՐ�,4��'�����.W+N����� jyt$X�'/���Á2OEԽ�*�f�F��'ƒ8R�!�m�YY1��[����'0�!c�:�j]ȁ/��LPЉ�	�'��d�$AI�}&,(qa�@�=b���'x6mhfW4 ��Z�' �<��5�'
���T1R���oH�!!6=(�'� $�V���?g�Ē���fF*L�'�݋P�����$��d���'��HdC�&�T�K�$�R���',��y�K)U��!���X M�T��'n��V�S�kC��RjF2X���O��d?|Ore�SB�+��D󪀹\'x��e"O:�ٓKSp��YtHCW/4��w"O*����YJ����@�q��"O�UzU�>s����GgP�1��"O,����('i�X��ŋ�'y����"O� ��L�Gb��
� qH�ѻ�"O:������/C.�� Ȟ -\<;�"O���P,P7GL�����+h��P"O�`�e`�z�B�[e�W)0ғ�|F{���Zh6��QV��`Wz쫳cU�6�!�M6 ���������8Rc�y�!���i��tsc��8�T���D�	{�!�d�!*�DɂE��5���:!#����'ўb>��PKи3nq�� HK4[A�3���<�'�,h��26"� J X�S-NZ�<1U�/,,��s�3!�ѓ`�T�<��A�W݆QK� �z�nQK��O�<�(L�g���,�w]b�
��I�<����W��[5ÍvG��Q�^�<�P�Y�n[�@�E.��sv��<����ӵ���{g���>s4�r�
=A�B�ɝu��j���9iء��`��B�	�X�f,x�N&D�҅�Z�T��B�	�7ȑ��O�hӰ�j���'	DpB�	=$,\ !�N���wA�~��C�	:*� F��_5��@���3��B�	�/�8"��ӥHtU��j��9��B��ퟠ��A��ଃVo��J��A�#D���խ�z��U��W0\  M��"&D�4�&g�/-�a�� �+X���:D��2�%4�8їm�.�
���-D��Ԅ��h�l ���J���H��y"iD5���� ��8#�$~��
�'��9Ђ�\1
~�I#��3=P ��
�'�Dh�RЋ��L# �+b`�O�%	�`�7�
���N �1�"O A���� ��� ��B���"O�a��	��)�֩���֧*ǆ�+F"O&�P���ھ�;��,I�>���"Ov�br�G-@��(C��jB�"O�%���� .����ϋ��4@"O�ᢅ�0u�<�1p.ƒ|���3"O���i�4����K Z�*�"O�1�䨊T���ѐ(�9���JV"O,�S��?N,��$�3��e"OnH���L�u�8cǓo�Di��"O����=찊�#C�&��)�"O~�p4��1#�aMַ�X�0�"O��[��%;�3�E�4���pQ"O>]Y���R�$���0A�h���"O�A��/K�Bd���D_&Z�����"Ol�1́	c���P�F3Bx��"ObU!��߀s�rɲ�#�	o�p)�"O�}�'�)�!p���9e�]!�"ON	�	ՈwhPa4@A�G
�  �7��|���ȯ"��H9͂�dtѲ�C,6B�8��	�DUP��@#�����Y/A�B��#B2�0�ѪSQ��}�#�lB�ɑW�"���y��1)���2�RB�	�A7T<r��:�����ę�
� B�ɫZ���e��h�>`C�-�0T8PC�	�K�r���( ��Iؕi�BC���,*pL�)�D��ӎx?
y��2D�\������+� i�L��-D� @u��U�(�Æ(O�9Y�D���+D�0��/��^��݀�(ʱ@}�$*R�(�O��c"��`k�,p�Y�h�cѼ��ȓy���[�#VA�ą6�p@��E�|����	5����D]?=X��D|��'$�>� H�yv'H�F"b����{�<`�"OH����o�4I���u��iR&"ONY#s�L>m:~d�@�� �~��q"O���#��>����)X�����O��$ɸ;����
�c���r�!򄃏k&�!��Ðk�:���#�9%�!�䚏n<p;S-Z7�P��L�����6s>Y�D
gG(�E����yBH�K��#�隲aZ��I�m��y"��5�=s�Kӭa���h
1�y��2\9��{T�Y�^�����y�%���,�C8"�� &�
�y��G7iü�����'��Q���
�y��=�*d��;i�4kGƸ�y2K2%�� �̆7Y}���mޙ�y��tW����'<�L�����y�b�z����D�:��#�Ƀ���'>ўb>! G�Bz���1(��Z�ցp��=D�0!��6kne�NZ8F�`�)!�7D� ���VVpƮV��8��5D�����ǫy�4�S�T',fXhB.�O�ʓ��	
&ğ�#��ٗA\�em,���!Iz!�3�!l������YL���#���!��@���
�ҨK�>��ȓ���'��� |1J��rx ��~n�1I�H�V�<MIq� �fX ��%eI�0R��D�7
� ����<uɺ��8}��h��A6fL��	Ay"�'<����ߩ}����(0Kq�	�'��������"s@�q$Y$��y�'�ȅ��b�~�:�7o ����'#���L�"�Ղ���~9~k�'~D|��@Lzcډ����w����'|1����0|4��rF�v�j�'{R@چ#�Jt��yv�M�C�h�H��?���?AƁ�7p�0�H���"8����UC�'rў�'Z0�Ĥ�|���娄d�Ja�ȓ1����B�Z�k��
-� Ex��i>��	�S�"x i�!QtPջ�ðj��B�Iw6V��q͑�9z:q!dݏϞC�	j����g��R�����Y��C�I�4���P2���wZΈ�E&:`H�C�v5T@�l�d�h��jC䉮:i�7ߵ �P����8opz����4��P�mX6�j�dI���)�.*�O��/���3U�2D��m�%:��܄�*���H�ˆ2Xz���CdM$O�x�ȓ_@�Җ�� ଜ �bG7���������΀1+����F�t��4��e�Z�p�@ ��dc���/ly�؇�C�wS�d#`�q��Հ��
�o���qbH�[�F9]��$mĺN��T�<	���i��A�B��S�9XE��I��LZ�!�D
/D(䅲��?BT��U�51!���Y��}I�D(=̱1рl�!��G�18P2#Ι�V9|esR��jU!�P�f\� Bw���0|���EB�p�!�!��m�ቁ~fЬ��o�!�_Jl�(��-|֜�$M1}�!���+\ɪ��p#ބ8_|�%�6!�ć)pJ�����hFr03���N�!�DB!+\�H����I?��:eo�9s�!��J<uܝ����:"h1@��_ ,~!�DI-d@N}:����*H�u��O�� Hp��.�/5x�	��1w����"O*�	�,Φ:t�KW�� o�U"O`����S,Zq�GJ];���"OƸ "��-�Hx��ȩ
�?�y"�$F*D�R	���7���y�I�!��us��=X��)R'���yr�R*!�>9X��-�
��q�"�0=����6}l���4�M�zT�j�@��y���+>� ��qO���c���$ �O���#Δu�}����JOf�h"O6����v��q����_F�)�"O�v��C�d"d
�Pa� ��"O�����C�؍�F`�0oX���"O8s� {Rn���
D��ȳ�"O"(��ŷ9�=d�ͨn��`#F( ��|�����'����Q�'b�t��GC_dTI
Ó�hO�i���o���(nK�6�x-@d"O���2�V�D�\��CGW8	VH�e"O�ق��RDfᘄ��5T�u{�"O��%�.t<aw�X[��88�"Ob%�3D�s�����3pZr� "O��2Q	�H�`����RK�}ʅ�'T�O��	DƎ�vX��D55��5"O�`ș�>�*b���/&}#��"|O"yy�d$f�qC/�;t�=��"O(-���'IZ,�t�#D��y��"O��*�E@�j�T����+n�>I;7��l�'��	
9�0�B�Чh��횄�\�0	�pD{�T�8�ʄ/�v���A֮�2��iu@��<9���ӶQ
<�IqO��W�f�����C�`"<a���?��7 �Gy|����������b�!D��`��<���!�O��ԡ#	!D���ЌD"'�Z���^1��=D� �@F؊G�H+�&2uR i>���	�mb�m��Ym�����O8i�����(�I+9�i�
YzР˷kL�0nC�	�p���d���:���g	�bP��	~��xxr(;������	�0�p�W x����	;{���#�kR:`�jL��Gů&�C�ɺeoV��g�!��*Ŗ7P��B��(W�@0KDbC:r���k��S���B������˃�*�5��<v��	{����N���F\c ���Ḳ��!a0"O>��de||4�P�&ɬ�r�"O��6`L�|T�j�b� zR?O���DB"
>��"JӠD��$�����
�'>��"1b�X��@q��ܧre }�	�',f���@K��9t���V��	�'�xz��65o��ul@�JJ��'�,-h'�o����t�	��)!�'<h��A��%Pb�,\*p%�L��y��)�S�08˕�R9$�K"l�?�2��e�I_y���YV$���0�>f܍�����!�T�6"&�#38��W*��!�DZ����x��P��	gK�!���l�4}�s��	./��2��`�!�[R����v��/Q#��[U�^(�f�=E��'Ɍ-�@95-�<��M�.5>�`
�'z���R�K� �Ѝ���F.�0�K��d3<OZ$r���_,X���k6ʥ"O��ѓj�1jJ���ᘍM�2r�"O��r̞�[tL���MؙSs����	x�'~:M �Ϝz� �4㏣%u>	�'��3ǁM�I��U���ߕ ���y�y��� �Tb&	�Nl�X�!A�3$�PК�ć��P�0Z���!=F�0�� v FC��"h��O-�XA�[y�NE+�'Bb���>+�@m�$	��_ ��'��x&��/���ιd � @�'�r�8#�Z�c.���I
��!�'�����12�Z��@���8M���)��<���<q�`�R4NօrE�0Çi�R��F{b�L7.�*��Ȗ�0݀�P��6�x�'D�$xQ�C+x��%- XJ���'����M�$%�T�WQ@H��'��d�Bb�X@�$fܹҒ�I�'��jF
�/w�ȃ3��3	}�3	���xU��J�C��h qf�P*l"Vчȓ+�tX�l��LIj��Z'e߆��'�}���??kt4�Tm�R@���4�yB��R�� V*�-b+�I��bG�y�!�*+Wl� o�Tu]A�$��y���<1gDTZ�G�H�F�ϵ�y�nR���5)��-S2d���^�0>9I>	0�'��@s `-"����<�I>�
�Mм
4jGF���mН>!v���h�r��Cl�1�����O�t`��ȓvk�ȵG%Lkr/	�~����.`8���"]�D�Z�h��U;1��]ʕ:e��&��##��p؈���V��$0򏝛\$���陨����	s��UU�Wꛌ_X61KǤT�O�x��y�IXLD�3�O_���`[2a�#q���d'��(_�R8�A�z;�xYg��w���|�IE����'>�A��,_0�j�seZ�!�䀣�'MD<�	Y+ z��F�|��Z�'�H���C�W�v��D	W�El��
�'a\U�GX��i��K%U �(z
�'66�J�%t�T�b�c�4#9�M��� �S���FiN5x����.ǚ���,�y�DiJ)`S�1+�z�[�%�3��'��{�kQ�;0ܡjP�M�BM D���yR�F	sԢp�gL�y�D��)S��y��S�t��5J%�p��q����1�0>iO>�r&Œ-���8sO�6�d��B��q�<�H�	?�]{uI�3yj
�Pҋ�n̓�hO�����)uf��֮B\�Ċ5��<	�*��+��-�d��:��P𒀘n�<��%҉2���e�z�.̓��o�<1��* �`�,����A��h�<�tI�mx��cCg�|*��d�<��Ӛk ��5M�|��u1Q��b�<aЩ��ؤ0b �0��y���d�<�Sd�{�Ġ���Zc��p�����x�jѓ�N�"f����(!��yB�6�d�qG�s�x=�ߔt�!���Z�aZ4�	�%��d�sυ�e�!�D[�u\�����Al ���4|�!�''�S�K��p��h�v�9!�$��PCr�\ ej����wa~�X���T�C�2u�s��,�"�;D��)���) ���\r� ��F/��蟾���e^�� �W� ��=(R"O�8{cT	fv���a��j�j�"OH�``�3f�89��K�/1�%��"O��ف�
���Nk&��"O��4��8����'
՝iall"""OR�1t����P�I%Y�f���"O� h8E�Y��p`�=��!�"O��xP&��}R�}�R�E3��dh�"O��3�OD�5��Rc��%S�F���"O�-�CcRh�p@I���C�|�@"OJ0e)��k����Ά��8p"O��XD��V]z���õ���a�"O|ȣU�ͭQV�(�L�.ϰ)*�"O\�G	?aL
7�OeHX*�"O�j"�.U�B�A�Z2����"O�	pѤ4QOY��蚀v�TU�S"O(-�@�T4�9#��W�3�v� �"O��%��8Խ�F���*�pȀ	�'��D���@W�ܫ���S3���' �\+�	'5�Ȅ�b�	���QJ�'	,�1�����X��=B02�'��Y�SH�?x9r��q��Ezhh�
�'i, KRhl�(\ ah�+f�l�3
�'D.a��g��7�^�S@�;d�.�a	�'E��
7�*Q���b
!+)�r�'�<t�P-�.
	;��_O���'���
J99�u��fR,І�rd̜§�#ɢY2B�ɱxS(���l��<��O�U�0�"�� vF4��E�Da�o�D.H�"�!u^���D�N �A�a�Д�4���_M�x��S��=qW�_5���k�G����Fj����*Ǯ!:�(����NU�Ѕ�zl��*����C�n% ��K�ͅ�=Ɯ����\��ѻ��t����"' �3�M�	D�,i��
mD�D��\����ʀ>2u�����np>���8�^�!�S2����HR= �ȓ*��Y�F�O$&�t��c�'\�=��N�P�;�V	3���t
S%Z�>��v�����L74O�)����9T�����	�ȁ��S�k^r�瘹v�����2�����Ͽ.Ѷ��1��6���ȓu�@�� �L����'�.����)&�x����${#�t���t䄇��b4R��c��̀�S�s>�ȓ؂ThFX�4"���D�h�����{�ܣ`�HL���M &���$�0��*�UCj-�.	;Lp��?�@x���Ch��b@�J�4L����0�le�3ǄN�^U��똀y@6a�ȓ P��䃝�4��Q�$й�^T�ȓP�^]��K�+>���Q��4cT`���9�8h�c��T��)��b�,g��؇ȓ_h�L�m�[ߚ����HEg����2p`t��%K�)����
��%��1��F=��37�4$��)���΁#10��	�=cc�K�b��B!�:M�i�ȓf8
U@@���k�<�4A3����}8ȵ�b��2�A��'M�BJ�`����"0&��eJ�#ѵdC���rV��!��oi�8ZR&�o��ՇȓE����D
$H�y�Ŏ1T ��T��L��ǟ5j���!� �-c��L���>q�Θ	���%�G�q<�=�ȓ?DAD�ћT�r��� �V���W.����]�d�!+W��J�dl�ȓwgl �p)��'���R�/]�Ml}��}pE��J���V ��<����ȓuB���7�WtjZq��R+JR���S�? �)feB"TDy@!�л��1ʅ"O�(�V��dl�d�ցYh/� a�"OZ��E�:���@@�K��('"O*x��ѡJ�E/��
�d���"O,E�e��4	��{�B�\0B�"Od$���Y�b4d�����V���U"OA�D�J&a2l��)��i�"O�5@啯/��(���O:���P�"O��0 ĉ$�^9SU'�M�|P7"O�	�%o�;�J�jBGB�A~�-p�"Oh��Ӄ�^�V�i 畼3����"O��x#
T���Cf]��F��"O�z?B���0�]k^��"O����d�t�\�T�I��txJ�"O�Xӕ��S�� �5�ߩh�h��"O�<���B2u	�`9 @�F�He�3"O,�ZaдJ��!��,�&ɲ"O�R����6���0��1�0���"O���t� �$#l)�CF6�Qt"O��C"�c܂���OT86�޹��"O �*��-EwP�y�(�1*�8@q�"O*� �o�!���!���R.p"�"O0ɐG���]����
��@ʡ"O��x�Č9�`�3�>v��`W"O|hQ2H��G���������5[%"O�h�&�#Y

Q�B��6��i�"O�����C�{ t}������jL�w"ONY�,Z<O��	���P�n4~��@"O���$%]r����fN�cN��u"O��@F�V�DT��o,3��[�"O�X�Ɂ�_�l��ՌO0�{T"O�h���ƬR��x��p�	>�y���S��ŀ%ʦW�xBwgI�yb�F9x:��`�RI���c"��yr(�ppi���#=� �"&��ybNY�LG,8�iǽ_i���f˒�y�HI#@O^�*��X�mI�]� �M��y"ċO����̅hUΝ����yRd�m�|�{�l�x�����ۋ�y"� |^�TP��N:WBl"�lX?�y��Ƙ_�(���9���J�I��y�NX�~$�Q[��E&*�(ɡ�c���y2`�  �l�a𠁡$5��26J[�yRD�2T���A��jY%CO��yb/��;�(��3V�Xg� DmG?�yR �,��	'�A^<p,�sc
�yR#$��I�d�ԛT���q�B��y¨�+$�8��DN�LҜds"���y"�� 8D�S&��
Bz�������yRW��a�@�R�L�:���y�+B�tQ��"��3G0@и֠�$�y�(A�f�m)�g��:/����A�!�y��ؗV�p�I��Ո/Vޠ:��V/�yblZ�L�aqFAT�HBg�^�<ye��>��0�f]�Z9^a��k�<A�`��/1 �`� ��'��;V�Q�<�r냘��	8�"�-cqJ�O�<w�)p�j(p��G�����O�<q� ����B�`
 ="��6��H�<9B�]|��`�cK� Ә(C@��K�<�TC�Y���Y�[�4�j��I�<ٰH�I�d� G������H�Y�<��GQ!j��p3���c�H0� R�<t�Q15M|�{d,#�6�Ham\O�<� �A���� ��*G�D9Yo$� �"O��@�	C�D���V�.0Te��"OVI$�J�=�$ �gF.#8��Q"O�U@`���$����%�Z>3E{�"O>����<wLE�'Ś(p�C "O�ٲI �%�� �#�ޫXmNYqR"Op�kI�c�>��v˘g�E�F"O8�'��?)�H���	d|I�"O�Py��޴�BC�4n��u�"O���''G��a�Ί-���!�"O����1R���%#��~��`U"O"�C%�҉@Ш	�A@�S���"O���%F�.�xq�g���z�c"O�m#w�	6J��t07 H/M�0dA"O��Yҁ	$� VL�Q|���p"O�����X�71��zV��c�Q�"O�E˂����U��;
c�ș#"OtX�SLײn��Ѷҩ
V$Y07"O.0*&(D$U���!�VN�qF"O�9�����8�OF�v���JE"O��p�� C�R�r�@ˣS�ĜS�"O❰���$Z^���s�x-��"O"XS�
) ��@���{[��'"O^��2A�:Q'��QEL]Oyp"OVdB�tA�4�!��*=�E�"O�y���=?�a��
�6��H�"O�9s��q���riA^'јv"O\�{����&5���!Q�5��8'"O�`
s�÷]0bw!YZ�9"O*=��蝲�(��Q�B�%�T�"�"O6y
��ʙ���#!��ڈq�"O���%P�-�z�rGk��Z�6`s"O��C1����U�7A�9K�05��"Oz��g�T ���h&��u�d0�E"O�<�SlI�*���)�߱���r�"O^E��:&��1��k�@��"O<T҆ŶQ|�(���Ů�3q"O��Mƞ%O�u���E��p��G"O�0��O�)���6�� Q�5�"O�E��mV�4�e��-H6��Q"O���t�^%V"�A���: G�<��"O*�#��L g��TP���,��Kw"O��0�'�kD<� !U�4)SE"O�Y�4��<-���B�o�H���s"O�qC�NQ�>���R�k@�Q�,iJ�"O�p�DƑ%��(8���?ofX��"O^q��Csm���D�U)P�,s�"Oܱ[U��	n���IG]0���b"O � ��A�МYR�^ \{$"O�$��T6tI���(����"O�Y ���wP��Pl�8D���""O�����A'$�ZdQFM�;Anfšs"O�������~�4�1Ё�.lf\��""O Y�ъ����-!�� |U��"O摲E��>)�� ��C���D"O ���"�0lL�9Z�f�q��B�"O��xB&V�=�����-d��{�"O��A"휛I
�"���6E� "OU��F�XИ��зv�B$�4"O��A��^cl0�[����B��x�"O���&�;%Ά����Z��m��"O���ȟ�7�z�!@;*��Q{�"O�M�pe�	(`D���	�/��EYd"O�17'~��r����I�F$s�"O� �	�O�_M�չG�ܫN�ܡ�"OV �g�(j���l�x�� �R"OT�a��,8�KA�R�`{�"O��ƀ�V�96�ՎdD���"O~y��a��kݠ��`�<v��� �"O& W��n�2�p�e�T�b�1�"Ovx�S=���0D�2ҲQb�"Oz����2=ެ�2���b`x�5"OЈ�獺P"$pu�P�M��"O
��䟓�4i@iG?f�K�"O�wOب=�T��'VVyp�"OQɷo)nx(��i��[R�y��"O��briJ')e(�&Jh[��+�"O���a�Ĥ|����P5$��&"Oq嬓��is���j��S"O>)c!�B�|���JO����B�"O���Ő)�(��7�Șxj`{ "O�]Y7-�)( ǈ�z[�`��"O~�sp"T�U�(`*U�W}V6�i�"ON�a�ق?�-��kN�:��@""O��`-ݞ+4xc� ݆%&b�C�"O�y��	�0P6E�ůBE�P�r"O��f�A5o��j7��U;&��q"O��	6��l�tUz�M�&,$�,��"O��q��OQHE��#�� "Or�@��,f�VIB�j�/d^ZEx"OH�٧.D0mmVM��^-\Ndܻ�"O6��U��r	�)HB�Fg����t"OV,��KY�Np6���f��
�"OF(�i?7~6�a�Ȑ07E D�'"Ox�!�T�*�"wN�\�2t�v"O�m�����r�tMQSσ1��)�v"O��	��D�[1.����U�<�.�r"O:��TGI5l4��"�
�6~8$��"O�̨VDS�q�]��Ƙ3z6�1�"Ol�0�k��=�d��Y{� Q�"Ox�yg�M�\��kRD�Eu��"�"O(Xzr�۟�Hi���̎tYZLx"OLh���ݏ:�|���!�{FT��"O��#_$��DPӂ�G\b���"O�ً�˃"~�2�k���+3cJ��V"O�T��+ �(D:�ŗrIx<("O��0���:=(���nQ�JLr��B"O��/����"��ía=�`�"OVX:4���f^Q�f�ƅ(�}@�"O� ���d��'W�"+^h��"Od��S�6��#�#�.E���H"OB�
�"�<(��(ǂJ7��I)`"O�ARu�E�B�QH0t��p*@"O�1 E�y�$XX��O�G��0�"OąA��W��a{�덬J?*=:�"O8��Ca�L�p媥
�'P��Y"OdPK�	ֿ?�� �
׍Bdz�"O�y�D��*�F�P�IڡZ�h���"O��	A8U�lp�Pg�;s��pju"O�#0���% E�y����"On��j̆�FuZS�T�ߒ�"O*��aP��V��1��U"O���U!r�`m���+}�
5�7"O^�Ԯ� N ��H|��S���y �&7+��8��ڐ9����'��yRF״��(#ԫ�24��Q�R��&�y�c���p�#���0p��e�R��y��E�kq�����U�"�� %E���y
� .yk �%0p0�t"J=��H��"OT9�S�=}��BQ�V[Q�`k�"O�H��L��]� ]8<̃V"O�0ٴ�W�mVf�Ή�}�F8��"Oy�!	�^$.q���/�F�0�"O<4��C�xE�I��4T��"O�����Ͱ4Q���ː2>���"OLE��ė��8H�)E/F����'"O$��<����G�@ؠ��"OT@Pbl�'{��Q��f�'��A"O4�F�|�v�k��
��%��"O��������VCQ��&��\Jd"OΡh�b�L<��޺p�4C"O��p��Ⱦw�1��� ��t�@"O��􏋨Y��X8q��"��Q�g"O���d�k��K�N%�ڡ�"O�X�V�X��y���F$C�j)3"O��KL�mw�l�បU#�q#R"O�a���D�gM�8�#D=pQ�"O�����ZB�|+&�N0_�ƨ� "OF��L�@���q�*ó?�ڵrD"O�1Btl��h��h��kӜ-R@"Oؘb�H	{��Uʱ�� +�m�A"Oh�@ <�D��o�a���"O��1��]�$�
A3�
�]�f�@B"O&,��)�*]�ځ���C�X���CW"O��CT'M�0�2��Dӕ*c��"O��x�G�_�j�9Q��{vr=��"O��9B��>
lP|2��+Z�P:#"O��
4^_��� r-R�q"OTQj���X�s���H�R`i�<�#"��`��	{�%"�����i�<�F�5t�H�e���,��Gc�o�<y7㕸i���b$�<���GPd�<i!�5q��lpE��b�X����k�<A�,ʂS�|�	B�B�&ƞd���j�<Q��O�h�Z����"���b�<q3D��*����<g�Ę��_�<%m�/R�p݃��@
9�v�PЈ�X�<�'⇠�j]�Rh�MA�Ux�SU�<Y����#$l<�)�N�<)�mʦ-PpS�M]N�]���d�<9���bΈ����D�D
<�"�_�<ie&�$�Ѡ5L�	k��$,]�<�B/ԘX+F=A*Ū	j]��$�X�<�a��iI�t��ҩ?�x!��k|�<�'ގ 8PHJ�k�$2R.�#S�M�<�&*�j�؇�_�E1����(Sd�<�`�"O�L]%���r��̐���d�<	���mV�I�7��wĀ��"	�`�<�B��<������9t�r���_�<9CDI.���:'n�Hȩ�#jI]�<!'o�=[�de�'�Q,��0�[�<I��B�nV$����h�V��K�m�<	� ��'�����Z��P	ԡBc�<A��"N�څڅ�9	��a�a�<Ip�������+- �M��R_�<���Ҍ1�`C�F�Rה�*�C�o�<!�" ���@*�Bɿ:����b�<q�%�������9d���+&�_�<�C��;R��t���ܵ;�@h�Du�<��iܟ:��t.E/x��|xLUX�<�U�P�f��x���M+y��T�]M�<ѳi�6=����]� �HIF�<� ����Ib5&X¥O&����"O�i:5�BI(�kH�r�0K"O��y���D�u��V9sё!"O`�H��)R[����Uw�5�`"O^�9f��&N��A��o4}�"O�%Ѡ�J!{+蔑���T�8�"OP�ks�V�)�e;Ge��EV,�v"O�����5siN������k�``�"O� �tIQ�DaPt�S�N�^���"Ox��的~��ePw���<�l("O�t:�.͜:��A۲A�oÎ	@�"O9��@�5:H���O���L�`"O.1�%��~>��O���N��6"O��u�ˋ:G�)�N��X�9�*Ot�A�'���)P)�-T��D;�'�"Q���h~���2�T�`$�t��'��Z��Սn7&e�3���D�����'�򱂇���c��Mj�T�/%8,��'t����A,u�1�2C�{0Tؠ
�'n�eCJ�����B��yL�h	
�'g�1IB0H��K�yqJ�	�'F�K�OF�Q����s���	�'2Hd���	][���-g$�9�'h"}�4�ݬE�T8�ph���!��'@���-�Z�2h���ϰ-��	�'dt�j�$�>sPR)0�Ω,����'`�,���<T^�����'A2���'p.�����L������<���A�'�m1��0{R�a
٭D���'�,�g \_<����&OM��pr	�'yV�󴊁g=���!�&JA��k	�'^�i1���)8rD�s�C!;�F���'��I ���?�>Z2��@�>�"�'-���0��a��)2��5���i�'6΍0d��-p������.��Mp
�'d�Dg�/:�t�`#]��z	�'><9a�B-p�~�y ˂�t��'�P�b�\YP�����i~^$y�'3:���\8Ŷc�'ج
%Ua�'�R����:% t���Lܨn�B��'G"ݒ��<@����7!�T�!
�'�T��R5f׊�`rAM�=�hl�	�'�l�8-ڭ&`8���-��&��
�'���JPN�� _�M��L�#9�1�'p.x��K���e����XJ
�'�P�viX�<�
���G� *�!	�'�z�V�J>HH�C��>T���''4`�4M������e� H��'�tY�1�>�5p��ΰ~�r�'+���i&�%���b,��'l����Ԓ�`+�B�X� �;
�'~���!�͓.���A7ȝ~��
�'i��;" �3'$N,ʁ��
yw~��	�'��$qR�W+_�j������nH�UJ	�'�<0�ηWڢ�js�C1s�P��'�:���k�s4La��7d��	�' 䜩�`�1/]�jE��s��+�'�*)e��Φ��Ĭ��rGdp��'�,���B�#&R�- �lڄm�$d�
�'�����G
N�K�R�h��P��i�<9�l@CD��o�a4@�Z��i�<�2��KT�Uv�;\؁�iHd�<�w������ɾp �U'�\�Ii���OyF=��딇.����?������ .�w�B �Z��FfQ�k[�j��	_��x�iV����L_�p�S ��y���>?�zMQ��߷% P�:��#2�X���'�a}2+'[����� �8�"��-�y��C����!�A	z� ��+L�y�cU�dT*!�X�1�
��TI��hO�'�"%��mh�H
A�3cU��0C�	K�"��Fk�����B��Q5n�,C�Ɋ\��2d��d�d(7aq�����n���J�$Bs��@�Ȕ�9^ �'�ld��	�/	BLse햓?�>ZƉ� �^��=}� (<�eK1��10W0qs5�е�yR�[a�|�fe�1sH�r$ݔ�y�ț�ڹ�v�K(m�x�X��E�yBJ��m&����`W�x�̈��y���L� ��E�"]ٰ�
�Bۆ��>O����	^L��4�Թa0=���+D�ԋ�
� �X�go�,����
*lO�����DW?8j�8�ͤ_ʥb�)'D�K5�Qsl�i�� wQ�rp'&�	J���'�^��U������OJ9��.�p���( ;�$) �M0u�h��ē�0=� �#������v�T=.԰���Cs �sG�������@\"!�X�ȓC�X1@X����E�S�|�Fx��)Z!aŎo:�	` Q�FJ���l�<I�OH�g��Lj�ɕ=M˾a�V%�M�<i��!E���I^e���3�E�<��@4:n�-�Ԏ�".��(���F�'Hў�'TZ�4��-3'6�j��hfC䉣8�R��E"υN;��30��@��hO�>2ɷ)Ӵ���mX��hQ �2��l�l�� �! E�/&`��˒�C7O���D��OIjty����XcdU=r!��@tL���󄒪`c�����]2W!�DU
 �1���؎CF��IW�בl��OȢ=�OP��[�o�:;�L�!���(	��:�"O���M	� wکq �(1CB�9�"O��AeYp>��V�6��p[r"O��u�5^�J� �+�9QdD,��"O���O�J�i�JL�M$�qC�-�S��y�-]'O��!�'b@'8RqR�Q?�yr�P�K�"���gR�^(���@/С�y2�.�Of�7cރu~�`Hr��F�6t��'��,�O|�
0ς
Z �U�F�\���ᕟ���)�O>��`"�O���q͘�.5���W�	`�'7��� �I���2X���A��oրB�ɜ{�xСE&�T��(��֌C�ɚv��Iqai��9Ӷ�p#�	6��B�I�f3����EU*��$1V/�L؆��ľ>���ҕJ	�l��ㅵ`��|�jLL�<E��6�HM�7%7e��b�F�<��iF�:��J�
Y2���f��wx��Dx"�ʚP�i.�
Ղ������*�S�O"d*�߀�&d�튞�t K>1����S�\=�s@�Ә*��bc��2��4}�΂`yJ|&���Ԭ�Ta�$ ��C��:$�̪�˪L�D�T &.Xv@���ѕo��$�,x��ᯙ)�L�b�|�Z�����#<��&��`Q�*�!��܃=�R�(�	�;*�� BV�	&�!�$�<`0�㊋S�~̈R@�k�!�D�"e���B�]�9�8�W�^�p�!�$ԙq���Ҁ�+����MT��Bx�� l�K6B�+U"��{׎hrD�'����<� hJ� �6o�Z)1� M d B�	�Y�$��s���5�*��I@�Qj�#=AQ.2}r��̞YJ6eB"G�!�h�26�9�!�d�tx��f�+� �Z�KL�0��)�'P��g��A@��c3e8�%�
�'ar	��G�q�c�5Y?|D�N��D{����ם+�B`ƄX�Qh�N���>��O�9���O�����-a�&0)�V�D��ڰ=����G�=����P�
E��jYx���I�<�2�ƹXO���1��9)�P� ��Q�<��lU�z�IDk�5�\=�O�H�<���5�ԑG��o����,�{�<�d����5�B,��"C*ࡓU~��(�S��G�0H���T?n�Ȑ1@��L�L��9���Y���/9)����ϝ�NlX!�=	ۓ��ٓV��w�*��kI�]Xj���x t�t�F3Ʀ��6i�����hO�>�ȇFEr<U( ��-O�L���J"������;��P3�@�@��Mˡ@������v�&�J���ȴ�ޖ&��i��h�,`��'a� �Crh�(�R��"O����G�zb���MU�^�
4�"O4h�Q�Y{��l,ƗY-�T�Q�$���F�D�B�9�"�a�04d�3we�-��D?��b8�;+:S�D�Ҋ��B��+b��O��d����OnU�,��'���f��7=�\`:�}4(@��TX�ܳ"�X2c�mp�K�'0*���'�:D�� ���6n,�@�'�"i�4�:S!8D�����֠:�9{6�^�\Y��1��Y��(O�b��bǡ��4����܇N���0�O��'q�)Cv*���P����Dwf�2��)�t`����2�%ׇ\����C�\���'K�M���"}:��	aK�x�!�@j�BD�gg�<�g�O	f�HU
F�T��*$��Y}2�'����,	)  �,ɶ��
&u���
�'H���b_�eeF�!(��K�١	�'�(�� ��/����-�.�d1��'=�dI�.ˆ.����k߆r��1�'������8t�4�
���WO�@��'8���g�ə*E�`9����M���:�'}@8qP*��J�RI��9S"�@�'&�
��G 5XPcs�&z�(�'���Faԥd�t�ӥNH�8���'�8�i�W $ɤ0�b3h��q��'Ųx����+|��rS�O���i�'~(��F�
I2 l�wjK�~�M��'���Kb�6'i��kB�Ӽw��d��'�6��@ګ*IB�����)w��}��'N��ه�ӭhɖ�CZ>|�l��'Sح�W!�&z.��0u����x��'����s�4-T�7��-P�-@�'�Ԅ���	;�X�@�/luP$��'�-r1'ڞl�X����f�n��',���D�
���4D߇J���'�Z�q�m��Kv��>�-H�'�BU9�'�oc�S�� +���A�'��ذ��O�x��е�'D|E�'k�	9�C�3��hҴ�P��fԘ�'s��qB��|�%����8Ċh��'���	1�8i�]A����e+�y8�'J`� 6L뺅ؓmD�]lhe�
�'��Y�&T�k�V0VB��&����	�'9�`9҅�r�'B�,�e�	��� 4u@��T�jSj�3���Qt�"�"O ���\*Q�XC[�ud���3"O��Xe����p�� >4���R"O������U�.`�F�2 FԹd"O�р&$ީ�JUb��X���"O�pK�8g<8�篅+lL�T"O����IC5D� 1�2-� k�"OFX(4���C���D��%g��C"O� ·O�"[)��)*�xl�Q"Of)J!��HА�1I�T+�"O�(���Ƚ\ľdc��=	f�h�"OZ躒�N�)/R�Jp��Н(�"Od���V
y�P۵���S�"O����=R��(wX&�Q�"O�50c FY��Q��T�^�Ҕ`�"O��˒���;� эQ���s��^?+��!��? ��d��"L�%ҷ�)b�庆�F0$(!�[�n�LI�-��j��M���� !�D�9�ݡ@eD��M��gд^!�D�;��ce��@h�I�� �!�$ݥ!IP�u���mW�����@�	K!�dЧ�Bh���ԬDQ�b�\!�$��8!�G�<i����E�>!�$W�*��l(��@�3i�CPo($U!�DS�&�BXi�F̯TB �5�+=N!�dO�:v8z���s�rd�����!��)I��rG�L�A!TS����!�$�?gDQI�hL�g0k7���!�D٭B�<��ә8&�Ȫ*�>5�!��1o8eY�DT+xG���*�
9J!�d��j>jeh j�<*(�&H��24!򤗉�U�ь��|?"ŋ�B��~'!���3L��#��O ��2��
=�!�d(-�P#���Z��y��@i�!�DO�q�j��T�j6���8�!���\J��Q�A 2�6ܺ�ڌU�!�DU������-��tp����ю;!�dʎ,G
�U&׷xd�VG�<<!�D�+�2���懆Fd��a��b*!�=yS ���A��1&���M58!�䊚F�|Y��Y�l�	���T!�[#��e�ૃ�#� ]�a"��8�!��84�q��G|�
��RI�!�ć1uY"�����&���×.M�!�DK�Vw>@� #��C�d�1EL�<�!�$K�YҊy11
�����RA�3X�!��8�[e].k~���ҫ�\p!�ʔ,��HȤ������7z!�dϳG�5�uc�7���'#�PZ!�$�����1׉]�$���aDۉp�!��		�0�p���h�<,ä%���!�$�/.:�x��dΆb��]��d
�E�!�$�o7����	j!NMZU Q!�DM:Fh�l2���&G�X1E ]=No!�D۠@�4X�SgDv�P�xw@\�FJ!��I�֦�Q5 V+v�!�/!�G�Pef<9ӳ9~`,*�+��<!��1�%��MIQ����&�!�DI	�
��@�Ή,Y�4XF�^;}!�ĎO�@�*WN�P z4��J�H!�F�B��ӅkYDF�[�	Oj!�$.U��B��ɩ^9�"g� !�dZ+7���R�(He�,�e��i!���6*���+��LS�(j
�HZ!�� T*S$�++ [��h�Tt1�"OD�ڄgM�^�:aZ�C�G�j�{�"Oz��q�Z3W�<�ib��8v�(��"O�9�3c�-_��]� 	P)n
"O=�a�E�`���j`� ��RQ�"O4�6O��^h���؍v� ��"O���E��l��
����t%��"O,`�X�_�T���&�'Ws���"O:a["�$BA�W�>s��{u"O��㌎�$���w���[���V"O��QKi�kq!Y;iQpՃ"O����Ʌ�x��&�ZK  �D"O�Y!傲` ����+���"O���B�,Xyz��"%lPD�"O�����S	p�ң����S"O�pXf�ۃ*��6m@w���J�%�O�}s@�֞�����������U�������.D�xAb U&�f�
�qz�y֬������BV>�k��'tѻ7��l����	�������$��N}rݫ7�D�b���b�b��})�iJ [�LB�2.�Dq� ���Sw7t�Tc���m��Wϲ�:�M�=%jh�}R�e�t� �*6�8. $����g�<�� F�c�4:"���x9�&��hƪ� �T�H���O�uF��O�a��çBŎ���ǣs���*��'�D�hT��~y��L����3����Eb�E�d��B�?ۨ ��-ޥT\"�I��"�`"ˉ�aS($�($]4��=Q4�ү�(�.O�\hp��)L�|�s@��+z��gF��:G�ԧF�xU3�"	�x�X�024O��_u���&H�>��}��eK���eg�l�.i�c��R�
T��_v���6��y�V@��|�0%N>N�<���-�'�p?��� 	YL%�VD������@�@�,�f]�mJ��
p�@�>�I"�̒<d�-�6D�����П��aPj!qL�ǵ6�TI<�C ��0)���0vf�"oMR�
��=q
�i%*�ZYz0!�+;���T垽	J�\�RO��J��bC��L]�ͻ�D.�!�J�8��.@�Y8�T��̓RL��R�o�� :�I��Ş�"�N�S�x�& �qn
-�T8���E !Y���D/N�ԕ�d�4B6:ҥ�K����@HF+v��	�%�FU:dȀh��px�BR]�%�EB���Ђ��G�.|���[�@Y.x��(m޵PU	>rJ�W�<�h1�Ot�;(D�L~���Ύ)�.�"fJ��Z�:DƇ�i����rM�/f�0�����Aap��KO�,�"�2�O|�I)	�q��
�/�����r�#>�p�A=h0�t�cD�9��(�`n�?�Ѥ�!Q=PQΰМ̊TCL)b	*��Q��$k�MȯM2�E�홇H��%� ��x2J�;"�ȥ�y��3��W�=$ޘ@��͹|�֤ލQ��lc��
�b<�1f��<�m�s)��!�"�"�cf����I�p	�G`J8%0�0����`3F%������CR��z�@y�U�`)ʇ�;!2�$��oe?^�W�"}
1iZ�9�n<�D�!D�"��$Q�JV}��H�Ѻ};����k����N�3{�|]y�M�7r{���v�
�d=��H��۪eח~�'W��	2�g
JT�6�Q�5�䠢��$ΐx��4{0B�7:���-��kS�T6� 	!s�ӱJ@~(;�O:6�Ji��Б0R4�t3q��?fÃZ7l��D��(N�\1�Do�ɔ)J�H�Do�(L�LѤD�c26���Y�m�,�8�b�U0Iaᆞ<u�1���(F:}j��� &raM؏�
��B�3�� 4V�hʄ]� N�(���ͻKF�j7i��X���	�̉�=�(Q�ȓSS12a�/r��a�$��$�P�(ue1%��ba�9}��9O��Ą՟4��{`ń�}Զ���"O�젤�V�i���b�*� )�=Oj���� X��דA��g��%�� �	W��@)��)N�6=x�
!d��(T �Lϸ�fσjR��� )D�D�0�� $ �S��6B`0R�&�G�L���IL�|j2`ފ}%���iY:+4$Z�D`�<�V��l����`S;%��YDc�4h1`���n�>	2ӧ����	`��t�Í�B�D���FԋX�!�dE6�X��ԾiN|�RQ�:���S-D�d���=�
R:b���wu�T��K?�O���i�./:7m�?H)�%0�˧,>�e��f��b�!�$�C�vɸ�`�@?�9�Ȭӑ�p��!a��>���#�kP<�
�g�-/���y� $9m����'�g�? Q�(�~�^�2s$�5n�r0��"Ol	R�gQ�b8�i�P��w�<!����w|�9��|��d8�# DO*� �'�3V�bM)n5D�T9�`�!EXq�4�� ep�DdA��(��I(ߓgS��[s�l�����L�Z�6���i�b��_�:�i��`Jl�c//X���{1&Йz�5�'�����"`��,���@L�\�V�x�+R�?�	��d�w��9M�O=����)v��V��&�;�G^&i��г"O@��ǟ�~�Z�GIW�ʼ���T:\~���gA>}�'[�r���Ç/B|�D���;bą�R�nHI0 hL��t��N�<�`V�]z���Κ�xh��"��Ɵ`#�e=��&���&�J,p�E�5�|"a�7G�`�c�gɊ$Lh��#з��=I�D	^�f$�6�O�� ��ޛL�4Qz��d<�S�lR��Ӱ&s����'�ZQ�GN�� ��� XY���}2@t�6-Z�^U�@-/�`MtjB<m%8��HC�'J�`p&�~����'�<#4���&�����W���P�O�@V�bJ<��n�f�� ��8�i}޹�W(_�x��)�1��;t�|ա�f'D�`�GHq�Cw��.��d�i���� ��g��m�K��s�Sg���4 ���"��67��)ӪZK��ȓ%I�Ui���ũ��ۧj3�5K��O2���O�i�u���s����H�O��A���jX����/7��}�F�5��$�4 :[��GC�cC��EL$����eP�Pya~B��KB��x�JH�d����hO�ѥbґt:ֽ"bb3�4��O6D)�ݖ!]4���Nw���'z�y���g�|x�I��D�\\���, ��a��
�4V���r	/�禅�C�FS�X[׃����h`e�4D��8pd� R�1d����k'�Ԉ@l U@�"E\�kA�ͼs�T�g�'Y��i��&�>�Q�ā^��	�A�� iH.U湨"��!T6ˀ�H� Tr������s��+�h٤��ex��j��[�a��� �/��Y.�����#� �[+��˱kïS���cj[
�ɕ"Jz����-50> ���,s=��R�N�y�i�00-yDU�jNrp@7-WF�xE0scБLL��$�p�nay����:k��,�;Z`dH��(��l��4��2'Y0���`�P�m��QC��pe#�T]����'V�B��pI�$R<��UEZ(|l� --�s��aD� o^xM�#��)�>L��I�B٨���ǉ�Vba�n�=5���(�E�T[��@�Y�AB
��#� \,�C��. 2��H	`���l!�:�%�$�gؿE<4EC�BC2		!l^"x��ɧ���N̢g[��k7��k~�4��"O���P��$9(��}U��x�c�<o�1[���B��)�E�!3���'|�X�پ��l2�K"/��'(�]��
<Uو�:b@�w$x"�)Z$��5�Y�!�|�^7V���`�H��C��+9�ay��#~�Hy��^�Vs���m^�I��ILoDB���7�!�M4qr��B$N����A�b]M��'���i���O��@G��)
��u�DH��`�^��y��Ù@z���EӫN7��נ[q�8���|�������3J^8%`�(sP|�'�vB�	�b�"\��玦L~l�D$ֆ h�C�	�p�(���\�0*�Ԫ�B�vB䉡�쨒w픈��QW"!.TB��:>�\h�7�_>o�d�	�%�*kxC�	�g�tV�u��@�Q�^�J���"ObQA��	�U[KL�T�D�P����yr���
� Ѐ�m>L��2�6�yBʄ_VR:��$ip�:�&�%�y���5]�8�`��7�H����y��C.Vu�X7!BY�]XT��(�yr�X'8
��Qe��\�8#c��y���F�N�b��*��Â��y2fP4.u�D�a��l�b4`i��y��Ǔ&s ��'�X�0Z�JԘ�y��>�,�{���X��[B�"�yb�ڊD�P�1�C��i6�U�p����y�{`%{!kP3eqę{U�:�y
� ���ٚ�he�R�^(�(��"O`�c��ԟ5�xaF�P�6����"O�(��h
#�T���N�=���"O|�:���Q8���FW��MP"O�`fW�=�*L/k8|)v��)�y�_55`�P���pgH�[f�L=�y��0Iq�ͳ$�=v�FC�ؚ�yR	�N���wk�;��[a�=�yB@L	!�� G�sFM��V#�y��+�=����o2��cn$�y�ɏ/�% �G��g�Rx9S%-�y!�M��J�>G{X8���y�o.n�YZT��;rPhj�MA��yB`�>��Y9�jNXh��k��0�yr	FO4����#"5� �V��y2a�	Q�B��!�y5.!2A��:�yR�,"|�h��vY0){T�ϵ�y#� ~T�A��.e��!�����Py� �%`�ڨR G��3��+�^m�<���(,���T�Q�J�V�ȀB�<���U�F!��aN��|X�[U�<9hT�W�d]zQ �f�>�
fM�Q�<9t@�n������ĹGٛ#��P�<Y����6�>�L\h(Fe�<���)\nP�q�\�4�@4�1l�j�<�R+p4�􎒣~Z4�c�[f�<����/R�@X�vE�99ʨs�![E�<��eYUt2��%�ސ@�l-Z�Ė@�<1�dݧNa�FXǰ�9�nGC�<��#��V�Τ؇䖵�L��B�x�<�7��[�V0`s慩?^hVOw�<1WO�M��@�K,tW���l�<I���c���
�H0,��C`�LR�<���V�x��ʐ:J�3a�L�<є�Z;�]��H�=�|�#���r�<QaC,)��O= ���R�$�:�'�f�
C N�}XK�n4��]�	�'�T��7���Kͼh�àԼ [�4!	�'����LM1M��!�C'L9
_`=��'��)Y�J�0:�� �be�+*0y��'fn�q�Ϳ;�x��FS�D٠�'/4���a�G_���r.�8���q�'8���$�V�w�ɂ�)�5(�|���'c���֤	O�`b@�Qq�81��'� ��g�Z��e�gm�&n�a �'B�ѱ%���I���~l܉��'.Xat������9�hh"�'��u���X\mX`yƅ��3e����'H�Rn[�Q���ȅ5)����'�*�FH�Lۆ����=dH��'h�0�ᜏ�����Z�Y�*���'uf�y���:�2Q0���oJd(�'�D��a�1=��,��mg�M��'�� �텳0��1���Ax1�'�~My'��ayzi�w��T{�T��';^�(%��=�A#�)N$\���'� PhE�Y:RJ�2��-O�ʕ2�'VV@(���U6����C�8��Z�'�5��k��)c�*>�0�q�'$���2e@6J�BH�����`�'�\�Bu蔔�t��vA�y�y
�'���Fdά]�@ׁ}�"���'�dY��?~R�Z`$S waA)�'�"�K � �v����;1ޱ)
��� �%����8��J)�B��"O�UH��C�Z^ D��d� ��(�$"Op�e�J{����Ab�6H�9�""O�9)��D:J��<�����M>���6"O{a�H�d�du)�ؓs.���"O�C��XVfh�%�߷` �(�U"O�m@Fa
�,4�<(�J�Դ:�"OF!S�� _����Ɠ%�03�"Ox� u�Fki�骄f]�8?<���"O��IvdD}��-#d%Ю7�A�"On���)U ]��2 0e"�"O\��g��2K��80�"�$2Mu"O�dk3��&@䭺�AU>A�ذA"O�Jv�W6@�z�pǃ��N�qr"Ofs�����\��@��
`�0Ӂ"Of�'D��l����/֋fP&ى""O:�Y!�)^tk$�D�n�˦"O�;4�5�ؙ���	�^l` �"O�d�4�ҴVܢP��ҚFs2X��"O*I�뚑�θ�be )Kzn��"O�Y!��Y5b�HhÆ�?��I�"O��Q LϰU'>��M
�d٣t"O��6��$0\�-��a��"O"���n��_�H��q�p�H(�"O�(A�X"e�%
Hb�U"O>D�B��N�`
�W5l���"O�@ch�]b���a�'T��W"O\�;�J�=B���"�1+vhÐ�'T�&�Ny��7fd���ȃ%E�g���y"�
C��YZ���(F���L�޸'
vI,*(r�@��IȄ�4�iҤ%�z1��}�!� �-0��1���j@!��`���b���?�&As�\9)����}�A� ��%24�@���.�p?�KZ�cE�A��-=X���M��}�RaئkB6l��q�T�J��|R�U.e���J�C�A,��A��@��O��ŬלX�Va�>"� ��Op�����e��0#T�Q��NP�yB�ѩ�JT��I�D[�O$N������^� �ɴW��l�DH����0�%N��}>E��O�TM���T�8 ��2&���-h��Z<9���I�^��dS�/[�ݳ C�% t��D��.{H8�rX�6>���[�,B�+��L��ҧ5�n�
JD`�I�R"�%;��4�0?a���r\Lx��޶U�|�� #�Z@3�2��E�ˆ�	>�:�`5��	ql��}�&����b΅M�~��UJL�'�n	�C�^�P�։�cIV��D�'}�~�b ^
k8��y��M�����O�XA��ΘH1x��I|�>��jY!C�bL*�FD�*�!�cL��<!��Ʀ7eP���	ѡ<̺	���6!5JS�#�+&�	ംV|�p��ɉ-6���B�'ؚ�ٷ��2D�����F�\�e�@���͏:B]`8I��\��u���b�]��.�W��Ʈ�Ge'	�L4pt�}�s��'�h����*�V��!ɸ��g��՛B�
d���;̚�x.ԠAH�,��))�	:V���6!���EN }ꑟ�X�P��H�1�,��.s��`����P�B|�⢂)M\�+����7���TQ��ƹY�џL+s/!%h$hx� s8$A	0�3���q=.U)�3��9��0�)Zy,�y���1
�ld�5Z @6|��P*��<n!�����%*��BG^���R 6ܸ�rCƚU��u36
Ԁ|���� 4�n(8�x 2��#J�agf�|(!��H=��� 3���F6�ͻD[�8�����
7��yL�"~Γ���e��k
y���3IH�ȓ��m��#��c@B��@ǌ�j4`ϓ>�qZƤũq���D�{�Ġ�r��9�0䳷��a|��_�� �UJ=S�< ���5`���v��4H��`�']H��U$�n^��x���
A�����dH0��K'�(��m� �w�(դ�;q������u�<�D!S�!hd@�T�i�l�G�ƱJ>EH"�`Jӧ����w���B��Ƅ�� �/�y"�	w&|M뒪ط[,��憣�yr���-��a��A��� ���d/S���a��Z%ApdyP6�'� ѹ��٩'#�fŝ]T�|8��ْg6 � �$�y��P�Njڴ�!� �|H��#=1�hߡ�֢}j�-֚Y6���mү`�p4�][�'�>�{��l�O�<dAK fuJ�:ԩ��G8���'�VYq �LS�!�(֍<�H5�2�Քz�L>���O�d���2�Q�=&P)�b"OR��2�W����I$vKh�i��iX��:��6P��5��C]�M���+�p!;p��60�����/���44��Q�IT�(�s4�G��z���� B���:���	1\O�1��(Z�**�ɗ@�X*q��d�IV��g ���'��A�ADrl#Bj{�Fl�j�f���	-�yB��i��:��gČ�I����X������!aJ�~�b�#Q��8CŒ�'�h睻c�. ��1E@b-��@Ƙ|��B��&�"�+dس`�p���j�x�B�B�cG�%�-7��qϚ<��[/��_>�K�+�t �@	�)�z<��	B8) ��ݎ,҈��}xV����@8������.?u�T��"I���<���F��EM�]�RTvNQ����#��n��'+ k�G�<�2���T�g��1�0Ɂ5b�zR��hh<���G�nEi2 �94mv��'�	?{"$PT�T�	#{�` 0h,*O�O%��ʴ�@���-�vN�ӧl��EI!�dȜ�B�XC��,�@!*��J"�����c���%�H���@�Hc�I����E�qAW�m�vY7�&O�(��vK"D��HTǗm�VL2�ǫ��	[WLC�E��+�% �ȐJ��ݰt�0�g�'ӈ�(LϠ1<\� �M�7kc<E��ka4Q�g�c�R�1�>faс�^��G���Q��k�3��MQ6g�:T��Kϩ+jqG{ҭL�hV��q���%���Sʪ|��/K�Ly�$ڮ1t9k�r�<Y��H�T�)��R s,N�zD�L�9�
�s�]: �D�P�X�)��s�P��!��&.Q��/�9�D�b"O$Y�ō���AN@Z���U�s�yЕb�8L�!��K�8x�r�g�'��,"��6^�Sw��h��Pӓ����H�j�~kE䐳+l����@��9��Ԡ��O�'EXl�b�J}��cႭq���kF�5�QMM`p%�0���Ojd��и�Ƥ\ ���,�d�b3��556T!2�u�8#c"O���!�6P(�(P2 _7~�d�T�IcE�#	��(cǑ�{B��>��CHO<�y��ٷ��h`�	|�`yX�߬��x�mC�\ؼ�C��UU�1����P|йu�J:A#����1}r�ıp%ǜXҨ�G{�dغnqbh��B %,���-Қ��<���H�F�RhzGE�%6.�c�M�0O���&�!	0H��u�(��d��qla~��n�X�1��(fS/���Q7,�PV��	 ��)ؒMZ�;���cB���ӚeX�q�'���
�i�%�*h�2"O�49���"F�i�F��-V����&"H�e���0B��l�X�r���k.���'"�i^�8A�e�q��8��Аx"'�0Ġ��@.YF�: J��M>�K�L˹dd��E�'�X!U�� ��!3� �w��m�˓%B21�3���e����'�h���AɟaOةؒ̍�8v����'Œ�kw�"y^����=0��msO>��S�2��ySw9�,�z#V�5*�(P��$� �ȓ-�$pr4-)y�&�)ъ�
4 ���
����4��E��O�lUO�� ~�5�s��07X� "O��h��M���1J�
H�"O���ծ=7dm0��$E�:\Y�"O\hC��Gt�A" �@���"O�%��x���`�B�!��A��"O�=J�	ИNM�0�$
� �NUh�"O���t��
���K��h�����"OP�)oL:h��@&�B���]��"O�%!��q��s���i�d�w"O�l� ���iwp �箚4C��;�"O��2����k1.���M�;���$"Oi�E�J&>�� b B��bL�Yt"Ov�����u�\!r�V^�İp"O���H� 8��`����/K.吠"O� t������(J�L1�D@�@Ob���"Od���ճbFe�1!#�YE"O�P�w+[�&�y�ؘ����t"O���KV�n�DA3͞	���I�"OHmp�D�Mf�͙�K�:a��m��"O��X��Mv�h�p�Glp|,�u"O�LR� � �>��È�sq�f"OV)"��&x�$���gը4t���S"O�)
!���!�ѡP{0�X�"On�BA�<p��.�?J}|�"On�FA�4h�0��^�d�B"O��y���/D5re�ȫ���!"OF����F�Z��U�'m�����"OiaTm��cr1��+��qks"O��@���|0,XK�ˆ
!���U"O���5_4Dl�I�W�\�܁(B"O����Nۣ14�0��uu|i�"OaZ���=0���%�o�t�"O��c�O�|k�=��N��D��q�"O"R�9�P᠗�^ XD�ʵ"OH�m�xӂ|�+V�
��@v"O60�C�I��P��v��k�"O�U�5B��*b^�@�/���� "Oi����ކ͛p&9�|��u�P%����?h��$��b���c���@aVx��� W!�ĀI9�dY�לp�>��?oB!����eK��Y��0PD�C!��Y�
Z�+��A�gr"E�_�g!�ċ��@`�£� a^�t�D#K�|V!�d�%��<�G,ľ9R�MA!,�+kE!��J����7CC�c�\�ڑ�K�s�!򤚧�X� �^���y�c���'��#<�����i:��<�c���W�Δp��:)���P']�<Y�lL5F��J>E��bW�90Ԏ�q�8� 4W)~e��A�1O�?�pb�7xL�2��׏� A��Œ%��b�P��E2�'����	�ҹK ���O�i��̕J��b�p 3%2�S�S�f، �IچE:�H4�&���O���u�lzC��9Y)�ɳgƂy��B�	�.���,D& Z@�*E?)<�B�Ƀ˾q��	�,2�>���H0f
zB�D[�#p�1C$z�)��[jR�C��4���*J9,p&/^:�!�dLT�d��CZND�qKP,V5aB!��9�p�v'�0/�>��V*�+:!�dR�>�J�A`�I�y�i����1~!���W��0�N;w^�i� Ch!�IO�����׊Zm�m`� �n!��(3j�-�;:]D�s  �!�䓍^�T��m��sN�\(��#,�!�d7���c��6�T��3�]w�!�d��`R����M�N�i)���PW!򄐐x�]�W�Ңx�$$��XbT!�ܒm���7���D0A��:g!��З)_~�����3:�b�AЂ�g!���*4GN`3�D�"E�\pKs"8M!��߸gz^���G�S��d��"Ov ���q���q��(�tHh�"O����% L�yH�c�j�܀e"O�1��M Y�,��P�̌�"O����L/ �1���J�$�d*O��eO�c�PA�]9iP^���'C�i�sj� >*���u*�r���'6p}��'ZF�0� ��L�d�>�Z	�'<\��.ˣg�6��m�X��ؒ��� ��Y�mܲ\9�������jp"O�ZVė�gN^<3����G�����"OT�y�����,���-Ǽs��v"Oz�;`��:H���,P�#��="OLY������P�	.۬�c"O�0�N�C���w�]�-cyYW"O�Xp��ε+O���$'K> ^h5�V"O���"�[�q��,:q�ŗP&E٦"O�2睘�>Xx��W26�,Q�"O
D %,�N\�Voȟ� ��"O� P2�XZ�����+\�b(�'"O`Ԑ�I�x���`J�
��d
�"O���n�/O>�q�<�\!e"O���у-b� ��[6w��K3"O��ZUcV�]:���P��"hh�*�"O�A:ǣR�A@�@�E6��"O
%��oM1?c��z���#�l8��"O�,���Q�^ř5Q0ݢ	JE"O�Ѣ�n:[�ҤpաV	,��`�"O����D�9���v�1"B��"O,1�B,ٹ]nn)��˔/6d��"O�z�,R��q��к"�f	�T"Ox\�sǒ�~��C��(�(�"O��w�ƪU^谰��%���B"Oxu����Lr��R�

t�*�B�"O��4.\���\���
:	�N���"O�4I#(����ĥC ^"�D"O�xCZ-���IՆ�jLr �"OX�����Y�4ܚ��^�vg���"Oބk��Y"vE!#Q�_]�l��"OJ�2�	A�b+�(v�n��#"OZ ɴg9u��"�� ����"OxQ�@�l�>s� N��@|��"Or�aa�^u��)�Ԑoʈ#0"O �е��//��Q3�9R^E@�"O�Q�D��6�bQ+��	6� �"O d2b�&1|�IA��>��a`�'��@���	l�֭��@W0��'M�#�лf:Ik�d�<(p�(C�'W4���ƃY�[W��Wt}��'�>��g_�#(�y��AR�����'�@ 2�h�a�|Φ���'��|�b���~�QY�hI#n��'��A*��Vd�B���Ε;�'_jE�d&ك]�
 ��Jx L1�'=�\)����F�I*Kz�F��'˖TC��M��œ�������'�4�ŬI�G�x�����c�`���&\� r�d�[�ސ��,W�~��ȓ<�����
[na�Lv�ӨQ��h��S���`'	~�\A���0$8�T��yz|�gh��$>�Yqրű�vņ�"Aр��q���Ё�ȓ#���R�b��?;�I`��r�Z��ȓT&��q`ɶ#-�xa��<-4.��ȓm��K(g��)��Ҽ
�	�ȓ�d��d�ϷR���ٴ*�ܝ��/�`��Ġ�� �J��b��n4�)�ȓFd*T�_��DЄ�͢^�� �ȓ3+\� �!B
��b�R$�z��ȓNg@�T̼);�����P�hD:ԅ�&���(��_ct�)�G�ZI���ȓ.�|���h�z�J�3���T4��q��!H�M�����/�����S�? �i �N��h��!�L�&���"O�����`��ܶeڔ�Q"O"��q�2d��M�o�BEE�"Oj�2d�;M"���H�D[^ h�"Ofػ�X8Ȝ;f�y\�4��"O��Ҕ��Qz*ĻD`'��*�"O*�y��%^oĴkЀ��hzj�"�"O��7
L�Mq�P L�fhZd�a"O qň[�m��z�/ū���°"O ��o[�$+*��.	�K�y�"OY3� )Zv\-�LF+N� �q"OB�S��M�1���2`Ԓnل���"O�]��O�ut\�(w�]�r��tQ"O֑��7�8�3�ʚ/x��;s"Of�	S�S�`p>�Ai�!ib���"O��Ò/�7K����	4��"O���%T��p5��fZ�g ����"O����C	����S���r�j��Q"O8�p��@�K�����ρ�D�(�0"Or|@�ɑ�g"�Sb�O�N��Ek1"O|e@�"Y/H��Dȯ�<��"O�
�.@�T���i�ݱJ�t0��"O�)��-Q|�hR�e@:-Q4��"O�(�.�;z?��8��V�X:�H�r"O���$됈����S6D%@u"O�5��)��G�l��d�'��c"O���b�ܝvQ��"$��
����yBO��9����ꀈ9h�I�/�y҉�&Ȯe��OCD�����h���y���&�>$`������@��yR����x8Wb�?y-.��dh�y҉N���B���n�Ɓ��;�yb텩	c �Bw���^����`��yB�D�HX��#ސ)[VHĢF*�y��GZ�"��F-�V�L�v/߸�y���a.@ 0bӆB�Ե���y2��s�T�Ң7���R�y�� j`Y3�.�6���C��W��yb��1hp�8#%�+�8���J���y�D���� đ�5ĬY�0���y��8s�:H�C���7ϴ�1���:�yr�K�{��;�%Y2t��D���yB��${��$���+A�5� ��y҃��&�F1�M%pzZi.��yb"W�wS���`Ѵ�����y�	H'략y�f�2!���`�L��y���<W@ahv#܌Y<��CG,��yr�Ty�t:�O�d�!�y�ʈ9W�\a�AI�0�F1� ��y�X�k�T� �J�whuf͎�y��ݴ(9��QQ�=�\�[�!F�ym)W]0���E䤽�A\��y"�7'��$ǬH�1"��QW�	*�y2��6ut�ؑi�4�`���K!�yRڃ/C|�v ���"+^�yR�в)��|��"L�9t�B2�T=�yb �l��#��w=E�$C���yr�C߈�A�"ʫZ���Ɂ��y2�ѐJP��ӍDQ��y	5�yR(P-��H��;8^֕�!�Ǌ�yR�$`V�	k �0,�"T
1�͵�y�ݨ���C�
�T����#�y���$�0�I��޽N���R��K�y���W�>�6ѩJ��Ћ6�=�y
� �qH��;sFH�%�� �RQk"O�Ŋ��S?g��i�w��-�04�"O���	_�@2�͔*���"O���.��ԁ͂��<P�"OLU3v��)�.؈��O9�"B�"O\ȷŮa�$q�g�9m��ҷ"O�(��(+|(r��/s�9��"OpH�&�/~��qz���T����P"O���ؔA�`�#Ӆ[�3�2�"O���7�V�+A��I6�&e]AA"O4��&nɑS����/AS\[�"OD�:�l � ]<i���M6oZ�6"O���o�g%���r ��a��3&"O��)U.�)�r�����GV0C�"O8Ac��"C����	4-���W"O��ь�o����D�9R�@�"O0q;C�M�'�P��M�� ��̑�"O5�T�>lQ�8�bT���"O��MY�C��8)�?B� �� "O Ń�[�B�t���$��4�"O�7JI8y� ��be&�T��t"OYQ��Z.���`���x�{@"O�q*V ���r��o&E� T"O"�!H8.���t�\�6{�z1"O�Y���?=�>����6^��8�"O�ةV��
1b�� L"t�D!�"Op%)����o���� ����S�"O�=8�M�n�����N��Sy6|�"O�u�k*v�3N��:PQ�"O.�)4l�`���i��g}��9"O�j�fס&�����+j�SW"O
|����@�܄
��U�[c Lu"O:�����N��<;�I�>~S:��#"O�E�G��_�:U"��O�����"O�A�́/5��9w
��~�=�"O*��ٻH"V��צOMeБ�6"O\`�qJ����Q��eҙMOƙ�S"O�h��ɞ� �C�v8�$j�"O�����(@�Qz��j>�I��"Oҍ��lW�
�b)�&d�
C�.$Hc"OE1��E�L�硋6~��"O��[�i�&Nv��b���l��1"O�I��d�z���p�zxc�"O�i�����v�pQ��;I�R"O؉��,�p˾�k'#P�o���"On9��M�&^�����H�>7r="O����(BP`4�&˧X�UcT"O��4��j�YFߚ�4"O\�ha��BoA�5�Z�y�l	�A�!�dN�vR~ȁ�@͓-�n��h��t#!�D�sL*�JGAȫ|������T�!�$���4X5�N4_z��&��"�!��I+��d�uK\4Bu�5��AԆq5�������M��OH����O��$iӨ�{�n�+@|M����%ibX����g������|f��{rx{Aчf�r�U��dlI�U'ɮg���i�nB����ɰ��N� v�čz�؆=D-z ��?1��I剀MCt#|����u ѧ�!LLXC�k"�Ҁ�a��ğ,&���ID�'��-�d&M<	�̴�u癮Em���{�,u�����O��oY�D�'ٛ�%݌O��8*� �]&i8�Q��~�Mљ6`�6�O�$�O��O�	}�JY�$+��L,!�*��i�J���%cڜ����p>y�a v۬�]5���E���Xi:١aP*��u���ևIP�(ư���E|���~��R� En.��AOD�s�ֈ�Q/�O���轢��[y��'��'��ia-B-:!��c,��!@��)�{"�'� H���x�z��#nҰ(q�m�!	��q%��`ش�*)O)Z��A?� ���RmZ�~JZ1�Q��=J������	g�i>��I�:�������#c�Ηh�p�$�M:+qj�ӶH8lO�u0�c�o�ԕ���(���]-E��qAQ*]�lRe��ɳ.(,�D�O6˛*U��.Up<�rG��y���ĩ<�����S'X9�Q�S6J�h�x�oZ�w��C���v ��A��l�A�t��6L>�7�lӐ}lZnyr�Ԗ�6��O�c?��CC�dx���>T�q+�M����I쟴���5�	쟰%>�x'(^�)Ŝ���a�,nu�epT�:���Vi\�`�:J�j����)VHu�yՆ�<d�)������O$��7�'��5�I�~�&F�������.�@��e�X5n=�O���<QB��5d�z���X�|�浓�'x?q��I��M��i��4b�����ƛ�jg�}`Rə�u�MS� �;b�v�'|�)����?Y��M�㝿w�p��%Z�y�0�Se-I6ykE�>�*���>�O��)@�J%j���l�Q���iC
��8$(������D�Yv�i>�#}�'�X�i6⋿x�|E�B$�$?����DO�Ov���Ԧ���9��>��BJ��a����ү[�!��i��ub�	m�'�j̋u�Fl�8p���U��\я{�N`��Ym�M���rڴ'��b�ǒ��h8�E�Ȝd?,���+	��ĳi���'tr�|�O�fI[)A�8S��Ԅ)��-��Pv���7*�j��P#c 	45@�G�1A�����k`ӈ��E�N�N�J�u�'�^����*_PS��S�^h����T�
�����O�lZ퟼�'��Z��n��
����PJ�.I0��ќZ��B�ɲ �ޝQ��J�<$R��T�T�ls�,K���d���'B�'��;J�`�� @�?�   �  A  �  k  v)  �4  {?  	K  pV  �a  �k  �t  ={  ��  ��  ͓   �  ��  ˦  �  P�  ��  ��  V�  ��  (�  ��  �  V�  ��  ��  ��  G  � 5 � � ' �/ �6  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A��!'��E�L��OL����A�*C�DZ6:��ga�3�a~Rk�>rk�;]\M�`��]����aC`�<9,�mj�pV�L���0+t. _�'"�?�w�M3s�r�k�$ޘU><�E D�"C��	��9��]U8��<D��"E K�Q�R�S�]�kg�ݳ�N9D�$B�f�$^ʄ�@��:)�M�d�<���S�!���D���<J07F>|9B䉢.����+�A'� QȀ�x>�C�	<,|@��Y�{�T�s��/F�dC�	�epA�`OE�5��ē�T�C�I�G8aS��+s�Ԩ䎇�jـ"=��T?y��HP�.�k@MP� "D��2��^�&�|��GM�/b<�eA?D���kM�ai�A�$
�x�l�At0D�(�ꊝWf艫f�H3nj��V�0D��"t� .Ş�a �o�Ppp�0|Onc�,�%T�J|�u��-UN�zc�;D��*��ň^�X'MD
4D8��9D���$瞶#^=���>��}I`<D��Z�Q;�Αel�pJ���&D��s0lʚc�@�� /^Ҩ��"D�8�`�+sP���Q��!x�����L D��Xe���@P��XS@����9�g2D��s"�Ð^��lQ���\(�X��o-D��
��������7��k�`�'�)D���ӊG�h����#�(hP�|�g�)D�@�P�P��l��+Ԧ  �dS$d&D�d��*y9xi@o�alx�2u�6D���J�Y�J��5-2PJ��5A8D��� ��R���-\Hr6F(D�\�0,Ke���Rρ�V�ڱ�%�%D���s�:Uy3�_\H9�*���y��ԥM�쭰tgI�v�<l@T���y�����0��|l0�C�a],�Py2 ĂF2$�ʑI�<��[E�B�<p��)dJ���U�)�<4{��E�<Iv`@�{^̀�nM�L��q+��DC�<��b֢	�0<;�CO�1�V�ƨ�Y�<r�]C�����7�h�+c�}�<1����*:֭X1Q�ܡ�l�h7!���V`�wa�6K&-h�_;&!򄟫q@��Ч���%��.W�iI�':��"�*�?@	�!Iq�U=8�k�'4|EB�H�$*�2�ʀ%�9 �d�P�'9X���Ry��@(���	|��!3�'=�5R�m6y�xE�VM
>t�{�C�2n�0����-�-x�ڦs�(B�7qrBEF)�:�h�C��\�0^�C��7a�m�'3p�p����YxP�>Ɏ{Ғ?������P���>��MȦ=D�� Bi���C�[�ZP�!�G
_�*�X���F>"�d^6RyF���
�&0|A�P�7D��e��(�X`4N�q\1�lwӂ ��ڸ���	��8 �`���B�̜S3�I	�p��DvӠ����%�	Xp&lYW�!͆0��'�Ƀh?U��w�_�e��'k�s��.Z���+V��! ����'�5�GU�����ڿ&D�ڟ'��	o�S�O�L<�EAW7��ĪŋW>o�RJ�'1�U�b`J@�H2�D�8�0P��"�'��ubԕv->M��+L�q�=�
��ē���KR�.iX�f��"�F��ȓ9��b#�D�,�Ĝsf��2m�F��ȓv&��y�e�#p<��%�	���ȓi�d�����S`Tqs���
[:��=��'��>��.@�i�S6O��L�%�]�qN�C�I<0h�I�,�'K���!N����O�х�ICa��G�S~8٥��� /�B䉀a��)��:Мɐo��b 
�'�D����I�&�*0�V�YEኈ�4�/lA� �?���iG퓳Ķ܇�\Ğ|R`�z��@��c�ssṄ��Ҽ �&K$�&Ib��c
�ȓO�*�c&�%����Q�M<ޱ���	e����v�DO`l�!�:��s77�O��Ŧ1��H�q�&Ce�֧�xap�Vrh<��F �b-H��wS�*U&�<SC�Fa���,�$Ǭ)��gT�<1k�~�d���*ƋyW\y(r.Le�<��ӆX$��*d�MM�,l� _d�<)�D�� ����K
��qP���d�<�C`�aW�T�b�1/��r�E[U�<0��! 
P��&��Dfa4��Q�<Q'nץx�@�u(�K!�0��D�<y7�K�W�����J��^�Y�Mv�<��L�LLI����%����#K{�<���O�l6*�"q��CSZ�*e�u�<!t�TuB�HP$�S�;4VȪ��Y�<�����r�fx	��1q�,ʕ��U�<15�̯x��XtiB/Pz>܉P(�K�<R��.]V�3e ��$�e�BE�<a�	�����+N=JN�[����<!c�$)p�B�ٸL
AS�O]t�<��G���]Bi4B�.c&a�q�<ɒ!	�]�l�a���-#��ct�c�<�r��c~���5!�j���l�_�<�޿�d�c �WBdL��E�U�<�s�%�P�"!U�(����X�<���V�t%nP��G+'�ث��W�<Y����w~pb��^q�DX��h�L�<!�d�%rx��Ԓ.`���R
L�<V�Z�"�]��bGt�$��fL�<)�S�.�t�qo�K��ёp]�<a/��w��������h������X�<�nJA�|���LҨ4R5Z���_�<���5�����L2��B�<i�$N�yj}cP�ϐX
"q1SOIz�<��Z�C�B��ǩK�����U��o�<I�㈤Z���qP�;����En�<)�N�-5i��b�"��ԑ�$�ZP�<���ʬ68�F�U�L���R�O�<�b�_��e��F�?T�e"#��N�<a6.� y�\���Ž�¤*�/BN�<�%�Q6^( p3�ǻp�
�Pc Q�<� "�OWC��	9unŌ�b`�"OfyÀ��Uђu�Ҍ�;�b��2"O��sU�<���[�=w�<�P"O��ɠ8�`�Z��)X���W"O���cG��;�0ti��X�.�4 T�'#B�'���'b�'�r�'���'-��
���-=>�ӂ� ipIe�''��'�"�'�"�'(��'-"�')^����ϓghrQ��M�,W�X� �'`r�'�"�'SR�'^��'���'n�0s�DݭW�P�s�*��{r.y��'R�'�r�'0��'���'x��'�E[���3��IJT6>ޱR!�'m�'�2�'�2�'���'��'Ht��fB
ju�0q���? �%���'Y��'6R�'X��'H�'2�'b�����ixH����V	}Q��Ҡ�'�b�'���'y��'��'2�'�^��A�#~=D���
*LZ� v�'��'3��'���'d2�'Vr�'�.���̟s���qW*�(C
6�d�'���'^��'b�'c2�' ��'��%���G��!8��� z,`��'7��'p��'�"�'���'p��'9*�ʃ�]�*g	`�'@"Jr �F�'���'@r�'�"�'Q��'x��'��X�P ŎM�-6���A�9Eo��'�b�'��'*��';"�'e�ݠl���dj@6Y>
u����@���'�R�'YR�'���'�7��Of���Le���u��7`��,ڵ�8�@T�'��X�b>�r���mZ9�@@c�,�mQ�a�!�y�\���ߴ��'���?�Vh��h��Ti��\1PБ/�:�?!��WQX\��4��y>W�R�O�"y�E�֌�f B��԰)��y��'��I]�O<�b�iId�j�ڵK�3!A�����>.O���#�+�Mϻzav���@�{ʬ���MV���?�'��)�S�
�Xn�<�E�O@��auF\�� �H��<��'f����hO���O��ڤmݔ4v)#�($-,���;O����mm����D^���ⵄդtj�Rr$�U��㟰ȫO:���O@��^}�	\�w� &���$DفA퐗����O��QG#ۡ/k1���Y�/k:�D��>ʠ���4d(l}yp 3za�˓��$�O?�	�fH���@�a�BP�V	���L��	�����<i`�iQ�O��<0Z6�g�S������[b5�d�O���Oz��5'k�4���$����hi�M��h`Q�In���@��������@e2����@U,A�C�W��I ����Or���Ot�?=y1�B)�@�4AD� ���(����O�&���05���H�1[T(2S��+ip�
���+LT���I���O�0I>a)OX�e��0�,34�G�c: ,i�'��?��j�3~nJ�r��
z��M�H��?�P�i$�O��'�R�'<� ş; �"��W]eZ���[=
ǜ����i��I�o�(`P��O��@'?%�>J��P!V�}��*B�lb��Ij����rf�`�Q	�C�Nj4x&�ٟ��I֟��O�S.�MK>�/7+��s�M��v�����䓶?���|�c剨�M��O�n�WMp��d�)��q���������O��J>�-O����O���O��S�^4S}�P $�f�&DR��O��$�<�V�,�	ןt��F�$GX� �X�F��	+t�
��[��$�O}��'��|ʟ Cv�Tq\����� 
�T�sw 0DGp���!b�~����
�|?iH>	���A��9a�@I��`�?a��?����?�|�.O`m1q�<�e�ʒ.�Pt���+3�n�	Cy�ks�Z�D��O�䟘q	�S�I��y�t�6i�&~�d�O��ᱧmӦ�A�yj������O�6 �Wo?E�}Y�m�:B����'�����@�I����Iӟp��p��&ѐ�J�����3^�a��NZn��?����?IK~���%<��w<�:p�A5DM�8�G��-I��[D�'�R�|����9>+��4OzE9����8$�A��?����'8O�(q��~�|2Q���@{�	�f�vqJ�D���Dl�O���I럌�	kyk�>��?i��.�&�Ye��L]�A�"/A��������>Y��?�J>Aw�^�ZE���1��h�84i�d~c�$_�!��nR���OR�1�ɐ)����sHx��[&TN1�gD��'|�'VR�ៀѡ*Iր��1]��(i��	۟1�O��$�O�lS�ӼSub�7Fet���%D�?�9�0��<a���?��{�2���4����_N�	�O��
B�L�)�X ٖC��p�t�sӚ|�S���I�	ȟ��I�l��g���r��i�/�~�RՃOjy"��>�-O���=�i�Ov��B=�&�٢�\�������Y}2�'��|���K�6:��* ÖI��di$�9Qw�h�����dh��<�Y�b�O��/!�x�Uc��
 �h+1L!Hzp���?����?q��|�,O`4�'[��
�P��G(�h�6�!�N�����M�r�>!���?��?\Vt[3�0�R�y����W2�+�R��M�O\1�"OM��������� ʸ` �Ӳ��]���ږ.���>O8���O��Od���O@�?q�� Z>|
���������I֟x�Iɟ���O���M�M>����3|xX�e��O4��@n_����?���|�p�U	�M��O�zrF�iM:p�B�d�^)Y6��=H��'�'�ǟ���ޟt��-@ u�Zg���Ԡ�)PYD�����X�'�<��?����?-�z�(R�eަQj ��+���%>O����g}b�'���|ʟ�}s�h&���c�#��a6L�7j�U���ϻE�f��|�t�O��I>I&�V6&HU�1�9J>N�·C�.�?���?��?�|r,O�1n>G�1���.i�5%�[��	������M�I>�'5��	ޟ���ܱW?l�Zs"�*�
I`FGY�\��)��tlZ�<)�c��0�F��(On!��E�>�����3CG�a+5;O&˓�?����?���?�����)�m�XH���[�>��Xzm�9ME�T�'���'������'�7=�.1x�#/C�L����R��U�P��O��5��iY�y�
7�p�h0`�\/n�P]j��@"i�� ��fa����&_�$1��<ͧ�?q�D�9-D���E� �3,E=�?I���?�����D}2�'0"�'Ό9a�R�TX,צ^�0� ��$@}��'�|2�8,�fU
�(ϚY��M���җ���Q������Oh���'?]c��O��ʯtERAxgA�T��ɸ2�̝[s����O����O���,ڧ�?	�?:�$�h�i��gx��谏X$�?�_�,��ǟ0(ܴ���yG��<gH��e I�mF�}	�!�=�yr�'��I.n�@nZn~r�Y�`��S�<RЩZS�A?�U3���_�6����|�R�h��ǟ��	ܟ@�I���[2�'w�\jwjH;Hl����Bjybj�>1��?����'�?�Q�I�x��aPt�Y�M�4���ۂi���ʟ��?�|
��(>Z�Ct!ːxN�ٸ"#�9D������Ċ��}���V2�O˓{B��xs�Ǯ[�I��ˁ�޽���?!��?���|�+On �'��B�y�v�+���=�x�E@�#.�fӒ�۩O����OX�D�wT^K�b��de�A�`��u(��i�q���
7`�0� ��ơH~���V3�TR�C��\���K4n�(�N�̓�?��?Y��?����O�\��]&1���e�D�L����'���'�0��|z�vN�v�|r�[$5���ੂ�K{�Ta����';����m�$��v����VJ�K�ꐪ�~3�<� ��Qk. ���'��$������'�R�'L�8;F�=<f@ЊNg�D���'p�Q�XѪO����OL��|:�B�	�pq�V��<T*��H���\~�í>I���?qH>�OE�@�OQ�o�(���i�.Z�bBD� 4j*���i��i>����O4�O�EH!だ!#J�o3_w��C��O��D�Oz��O1��ʓq/�f�ʬ/KF���ѝs���@SS��y�T���4��'����?9�J	�j����!8u�x��FK��?��b��9K޴���:��q���Ԥ  d%�fW�`z�a5ɑ6�y2P���I���Iҟ��I̟P�O�^p�u�;
,��A�U���T/�>)���?�����'�?�u��y�ΜV2�`1*�%��h���Q�MPb��iҖ�K^��y��M"j'(� n,1�
�ж��yb�B������m�'��������9\?d05�ĭG�x�#F
X�T[\e�Iן ����0�'l:��?Y��?A �^��� ��fI������A*��'U���?�����r���
F=w�����	vuz��'�mca)��ܢÞ�tN����S�'�&a+��LAz@I�1����LT@��'�b�'���'��>E��&7b�3-�.e5t�/�D ]�I����O:��N٦��?�;4��]U��"��(C-�6u����?)���?� D��M��O�n�6��i�5c=��`A��Jm�a�[4c9��yN>�)O��D�O��D�O:��O�B���lM�"!Ν������<��[��I럨�IY�'e� ����*DZ��K�(K�l9Y� �I��`$�b>5�0K������-|�Pr��5���nZ'�򤒋?��-��'��'��Ip�� ��%�
j��|@�I����	ǟ�����$�i>a�'7lꓶyr�S%o��1�ui��8Hv�)����?i��i��'Z2M�>����?�;D3��auDK�
E�]{d��>��*��ی�M��O� �D�S����#�I��(љ4�Z�6�|��d��L����0O���O����OF�$�O�?�)�H!�^����ssm�ڟ��˟8��O�ʓgꛖ�|�2��P����Z���<i��'������-Ǭӛ�����Ã����+e<;���F%��y�l P�O�O��?����?���{d@q䁉!v���Y�����?�+Of��'8��ן�O�Y:�R�?3
U����0�����O�9�'w��'ɧ�)W�^O�c׊*�0��'M�pK���	�ܐ1�����- �B�]�I�Pi��;2n�1|����Y�)w�T�I�L���T�)��ky�sӤЁd (%���wcU�h�( �0O��d�O��nZD�S���������D���p��3�6(�e蟜�	��bLl�V~Zw���`��O�6%��� ��Y�AW!h���u&�i��\��<O~��?���?)���?�����i< ��"j�>f9=�3�0�$��'���'sR��4�'�v6=�r�����	0@����N<-B1#�O��D4��ݶ�7m~�TI�oںU��p���?g���dw�����f���A\��Oy�'O�Cܞh�n	
�f�5�Ą8� k����?	��?)O,%�'�B�'B�Q�e��d����T�����6U�O���'��'��'�ƨ���>\�h��<iغ��O��q��K��uY��I��?	��O@�.BmD�r���l_^�"�I��odR�'Cr�'���s�	
!��^P���N؆!,\��ƌ���O2���Oިl�N�Ӽ��I]=-�x��g�Mp��1�!��<���?!��
q6��ش���(C�\��'p�8yT���_=t��T���q�P@��#��<�'�?��?���?T�ںL̪يg�:�\m��a]6��n}�'�R�'��O���_�J��#ā��y�'%/5���?����Ş�v�x`�Ǩn�$�	!>:,�$�Fn��'.4YE	��Ý|BU�P��;�`=�ਜ਼�kL1��Tܟ��	ڟl�����Gy�.�>��bh��Q��їE�*�$�F�{u6�9�1����N}R�'WR�'�:PQu��e�����%D�,�h93�D_�L�����0�EɌ�S��k�c�S���Ö+Ű>�
$���ʎ9Bje���k�����������I�����%�	��K�CRc�������?���?�'_��ş��ٴ��=��A{7+8dB=���&*Ɔ��<����?A��Rh�ڴ�yB�'{�m�����	�x���L2���{Do�Pʌ��Z)�'�	ʟ���T��=p����ݣ*of��ơ�$�0���Οx�'[�ꓜ?���?+�b�a��Q�6]�'��y7��@����O��$�O�O�ӻ.n)��B��%���R�ƴ��ֵ�쌙��'?�'c������Yj��ԅp������$+z�!��?���?1�S�'��dզ�:f$�'�rx �b�<`fx=kQ�}�0�IǟLX޴��'����?Q�a��J��݁�cO,6�����,�?��O�8(�ڴ����`�!���R+Od�;�h�x����Ä5gÚ��9OD˓�?����?����?����I�D{ x��:V�:5+��/e��'���'R����'�z7=�LٲK�R�N1��,�/�2�b�%�O���5��	r�Z7�s���A�_��c�Y�TH
��Q�|�ܰGع6���'�D�<�'�?���T�j�������%�@M��?���?����d�n}r�'�B�'��u���( TT
5C!��\ƛ|��'#���?���'�*�	W�s�YĨ �?#ք�'�`��[�	F�	��������	�'���ufSN�!���g+Ɓ�6�'Yb�'���'��>�	2�B�
C4�dI�@l�1�I%��D�<i��i��O��N��[����
��Nې���O����O
M	�)n� ��,��&$�,˖,�:e3�eH4�B�G�L�q�G)����4�����O\�d�O����ܚQ��O]p��-{p���Pʓm�	ɟ����'?牘C�-�b�XZ�	e��"(=b�Ot�D�O��O1���JĨ.�专�ݍS����ѨͺJtt7�=?�"B�3�,�IT�Xy�냺Ta�,�7��N�d��D�0>�FW���I,��}�F옜�։���7U����/�MË"�>���?q��R_�ydD�6�� :�e�B��IPh��M��OBu&V����%���� �`kƼA�(�憲�F���5Od���O��O��$�O^�?�b���s�&-{0��2F���ڡ�
my�'�d��|�����|r�T75��΍~�|�T�pU�b����jy2ǅH�֚�X2�NF�DU$�+���*���o�|��XZ�'�@-%�L�'J��'��'�ر��#]7HY���A?v��L��'q�P�Ы�O���?A.��A0��.G��=�4�Yf�� ��D �O��d�O,�O�S�g���[��2n1���s���<���yV�L�jC���\y�OC��Iz�'���j�cI�or"����!>����'q��'�����O��ɬ�M+�H�]��qs�K��X	�j��<����?���ic�Oz��'�r�ЮR{���b�8-��kBb�6v7��'�t�ӳi��I��v��e�O��-�,J�̺`���f֏>�������O��D�O���O����|"�I�?��h���� E�� ����
��ϟ,�I⟠$?!�I��M�; z����
0�)��/L0x������?K>�|��P>�M˙'�<�[$�@�M�p"�"���\�A�'�L�$K�០{��|r[�������х��i�m� A����qiU͟��Iן���ny���>���?���X�(Pʷ�N��v�A���;-����r+�>����?QK>����u�d�{s�
zLs��Yb~��6ĠQ4�A�$��O
���ɳ$���@]���(M�}I~�ksm�I�2�'�r�'�R�s�u��"Н�N0a	��U
A�Nԟ<�Ov�$�O�yl�Q�	���F��i���S�.t��b ��qɮ�ޟ��	���x�f���̓�?ŀN��)�|�? 0Y�����ld���k� D�����#3��<ͧ�?���?���?1�-�-#hl�3Ƶ�r0���<VJHʓ{b�I��Iӟ4'?��Ɍ�敺�(�X����U�x��O��$6�)擧$n���,F.q�5f����	�S�ܿ!���'�R�b��ğ("�|�T��2VE/kPzС��P��BM�������x�	��S~y�>�� '��Di��o,8|Г�Z�R�X���;����De}��'���'�6�J�F�e�Ȱ� {���*��ß3.����̺v�1M�Q>9�ݜmƐ��3T7v��s��(`>��������I͟���f��g�:��I\�t��K%!O8#��Y���?!�O,�i>i���M�L>AR�\!!��`�� �p6��9�-�䓐?9��|��E��MC�O��W!@�r���8"ܨ0�t`�*�|q����O��kJ>�,O����O����O
�᠙�
��aE\�0&p}"���O����<IZ���	ɟ��	l��A9�����l�KF�2 �����N}�'�ҙ|ʟ>T�!�WE7h\)���k�����C�3�I;��Εx�i>��&�'�P$�t��A	
q$|x��O,\����ڟ���ʟ@�I؟b>9�'l6V�`U���w!L�qt$� ԋ�a��D�O���NͦQ�?��S���ɍ{	��Զ����E�{�~��IßC+����'D�E�eܧB0�!�ˈ�G\�	�f�6v�Γ��$�OT���O��d�O�$�|�4d��\9�i�(����R}��ß��I�L&?�ɗ�Mϻ�J�:<[j��P�"a�����?�K>�|r�a��M�'���i�"L��\�f�
�9���'-¬ʁ�[?9H>�-O���O�i
V!������3k�!���O��D�O��Ľ<Y"V��I����ɠ,��K��ՒS�h`�V�I�Q���?!�Z�����p'��i/߄�xG�$+���.I��ɏw��`�	�]��b>�hG�'����I�o��8��� +�͋��6��֟��	���Ib�O��«H����ι-�� j����S�h�>����?���i��O���(
7�a�CmM�a���>"��d�O0���O�4�|���{�R��<�J܈#[&D��J�&#�JQ D��&�䓣�4���D�O����O>���(z�8l�U�ܤQg�a�� �{�˓j���� ��ş�'?)���U��ۀ����T؇��M�On���O��O1�i�����6C��4�Z�����=�b6�.?aEg;Hm���`��dy�H��!���脔i�����4���'��',�O��I��D�O��ö!/�q��A�������O��m�U�Qp�	�ĕ'~��:�J]�x���)aADŲ��Wd����� u�
�f��At������!�l����Jպ0ZTe�p/m���	��H�Iß�Iٟ�R�1;���z��2:�1��Z�?���?ɒR��ܟ��4��R���h�f��d�`&[�F�:H>����?ͧ/A�0ݴ�������rL�Kt����HV��T ��i	�&���$�	������O����O��C�ԮE*bJ%�2�l"1?����O��q���dyb�'�响A�ڱ��A� ��h�@L9\��{�IџX�?�Oֶ�`����#KF���h��O��k�20Yv�Q�4F6�+)O�IX��?��%��@ �!4O�!ή\3�ط-D����O����O��i�<�1�ixXy-Õ-�B�T��*$)���'�r�'�6%������O�۵�B�e�ł��]�,<r3��<q�e��M[�Ox0�Aۖ��ȣ<QB���v(5�S�=���Sh��<y(O��d�O:���O��$�ONʧ%1�aB�C2��ze��|%"��P��'�2����'\6=�L!��aڽ82�`���đ+�.����O&��/��Ɇ���6-d���6��@X�(;E�9��c�z��	$@�W��A}�wyB�'f�%�~���Ga	rz(�W7e��'Q��'��:����O���O
���-"߾,y�b]�i�$ ��1��O�-�'X��'��'ɜ��vI@�dP$uɥ�G����O�HꐋG�:s�7MTp�.q��O�]Е��6q��C*�b�HJ���O��d�O��d�O��}���0� �9���,6��3⥛�#K9k�hF�Iџ�	#�M���w�;6�(O>�����x%��'���'�bf��J�v���C� ��/����X�
;��R�X2{�$�C��(J: %�����4�'���'�"�'Il��$nU/�~qTGB� V\C�P��
�O�ʓ�?�L~z������L@	�|Z$�L�C0	Z�H��B�Ş
"����5lb
�x%ҢD"�'�9�dQ�.OM8�B��?�E!;�$�<�Ԫ@1&�P�z4��"XV�`x��1�?���?���?�'��Z}��'f!��}U�+�͜�xx��'�x7M*�I���$�O��/_`���l)O��-:&A&oN��Я^�M#�O�9�A�J���F�2�	���)X��	�"R�\z\b�2O��D�O��d�O:�D�O�?���Ȃ�$ur���H�-e��D1�mCiyr�'����|�W�v�|B��J����Q��6�T1������'�����ԨD�F���zì2� �=)�/��A,T胶n<2������?I�b%��<�'�?I��?I4J	�*�"��9^|��ӓ-!�?I���d�y}��'�r�'�-V����@���!��R���b��	�`�?�O���a�)� Q[�M	T��8�� +B�MV�>�� �� m�i>E� �'S��%�d�&
"%԰H�MD #{� ;f�I̟ �	��$�	��b>��'(�7m���n}���V2u��e��gR��On��¦��?Q0P�,�	���*���!!�����:�̰�I�0ЫXʦ�'��m�CI�?ɤ��	��� �.I:���&����2O��?���?q��?!�����	>|5�`q7�Ʉm�-�g*Cu��'H��'����'��6=��[�a�8 �����H߼�����/�O���?��	��o�f6mg��9�-"9�p�D���'���pGr��"��
3N���&��<����?Q0�I}���Q'ʠ$�T�a���?����?1����PL}R�'j�'���
$oP�I��d�d 	�#\�U�$V|}"�'l�| ����2LH�<nȡRF
����D��8yjdp@-,�1�p`P�)� ���T6|��!�܃���KD.�	� �$�OP�d�O(�D3ڧ�?�F-��v���CēeX�a'2�?A _�8������޴���y�Y#��ғ��o',����y"�'�R�'M8L���i��		D��h�ݟP����J)�J��g	"r*-+�"4�$�<���?A��?����?��ׅe\�}���4����,��D]}b�';r�'U�O?��T:>l���
	*{h�b�;W�X��?�����S�'Q�\`��H<&��q #�HI�I����M�Q�DJBHB�Xl�$#�d�<��υ�3Ŭ����]�	x0�[���$�?���?1���?ͧ���Q}r�'�b�Y�ͭG�D �	��'k�@��'��6>�	���OV���O�c���!%�2����9d��y b�1h�L7-$?��#��	(���Q+u���b�M�4
A�Q���KC�~�,���@�	�$��؟8�"SA�9�t����P�8����� ��?i��?1�[���˟���4��B��t�g��2jp>���bY>I��bL>���?�'1�<kܴ���P?#��R�S�<��
*g?:�zf��nZ+m��'z�i>��	�H�I8+��Ĺ�l�g�`ӐΆ9/J�I֟`�'�ꓮ��O�˧2vi�fRH�����_�V(h��'I�ꓖ?����S����7���a7�[!x
���^�/o>�yC�E�mv�=��Q��S��R�D�	;
�Xhf�/��u��K$,��0�Iʟ���П��)�S_y�MeӜ8�)�u�U�Q���@D���5O����O�4oZh�H����ˠ#ˋ<�40d� �䕉Q������ɭ]��ul�L~Zw�d @�O�䵕'���CF��\$FQ �o� 6�Q�'��I�����럌��ڟ���[��!�,g��y���#=�10 ���/�듬?���?�H~Γ>���w��8�G��!Kµ�t�Q�s����v�'���|��D*H�Z���1O�\x�,ݫ
������R�u7Oнڣ����~��|"^�,�	ҟ :�o�&=�ŋfG�]�%Cd*���������IzyRD�>����?y�%�9�_*�! ��=B�
��DS�.��	֟���F�	^���v��e�F��+�ު�"�N�`�H�:�U�|���O�U���c":����%*K
eV�Fe�P�����?1��?���h���$��gL1�ġ$1�T; 
��	iJ�$�l}��'QB,p�.����@�C����r�d��k� �	ٟ��I�<Hq�ɦ��'�\l�d��?I��^,���V G�n�CġB|9�'��i>���ğ(�Iџ0�ɯd4����$��8����kѺ��'m���?9���?�J~2��X0�	ŀ4D !��%q��A�S���	�'�b>�S��@�`8B�Ȇ�#���Q��9�X�[��+?i�蕣sZ������d�!x��A!�ψr��E�@�������OR�D�Od�4�t˓Y���� �c уD�PEjջFyʭ�à�⟤�4��'듧?Y,O��X���!lމK$�?K�t}+"G#'�7�5?��m��{0\�����'������`�\ŋgH�"K���aen��<���?���?���?َ����#R/���9Bb8�
�O��X>p��O��d�g}�O*�}�Z�OXe`���A�(1�����L:Ӆ4���OL�4���*��V����"ܲ O�x ���=98���^V>��Q��ilFI����f�P@�&d�()X�9�熕g���W��u~n}R�aG$��a�ak)�����6ct���c*oe�����:y2�hʧDM�!�@QI7ET�_�2��+)�aR'��`*�������R��� {|�����I(����'�&�isE�r8d��P'<�B�*���[�@�+�ZN0t��ɵ��Pfi�z��&�N2 ղ,k ��o�np�1�h�� ��te�i�'昍t�@B&&ʗo�@�+�NҝM=n�t�N9_R�(E�ˠ]�R�vӀ��Oj���OZܚ�%��"md�b Hƃ23��p�
b��̟ ��7!�Ld��m��TrV�V�7DQ�%@����$�ߦ!� ������M���?���?�R�$���? zź���J���@Gϣ�M���?�2��?QL>�/��p���iD�-��`�q�މ��$ �}ڴ�?��i\b�'��'_����D�t8H�G�E�c4p��Am9s�ZXnZ,�6��?�(��h
�2O:��T�? ��zdK�^D�J�Ѳh͠����i���'��'W4����O��	%W�D\�l�52a20��!#b��q�Bǟ8��q�D��ȟ��	," ��Co*|X��\�,I��ش�?A�Ot�	Xy��'�ɧ5��"B�|��B�B/R�b������C��
��,yi�D�Ox��O\�O���4�D
��M��Z�)ߴ2��Ihy��'F�'���'�ٹ .�?���C��V�z0����+�b�B��y��'��'��O���S- vY�.�Wd�
1��<�7��<�����?����̙�'F�t킢BЄM3Fl|�����B8�y��'�R�'���v�O����8s	��b
�7Th�:��1;��6M�O�O��d�O��	�@*�	9L2u 2�Q��`�N�$�r6M�O��N�S!�D�OHi�Ot��'�&�M�v���Pz���"@��<O���O������c���
�2�r�ё�[J�r�;�KJĦ���in���ɲ�M��?����?�_����)Ůa�e맢޸5�$���%��M���?Q����'���(`�7��J�DҀ�ƅ3y�E��m����V�'$r�'���'%rP����ǟ�"� h><�cJ�7&l�*��	��M{������	Ĭp��$�OR@�ff����y&C�Z ��z��ݦ��	�l�	�<�K<�OL�D�?-f����<30F�{�+��H\�V�'B�'�H��yB�'f��'Z���G(�`	2 	�:,�fK��g�8��O�$���O=�� ��&�؀s��2��Ea֐x��'�ʼp�Obʧ�j�'nJ�Z�픷a�>�7NߎF0(Y�ش���OX��*�I˟X��<�t��/\�4Cd�R%eA�lZ)'��m4?i���?ͧ��?iw$h��8�#�jY$i��`�Z���O��|��xyB_.�MS��Wz�ɑ'HQ�<���$Z�z0��ݟ����u�S� �O4�C�.?��C��r�p�3gFX�>6�/������'��H<�!!�+3�yj�n��0��9z�̃Ϧm���0H��Nwy�T>Y����x�i���t ʷl�Զfi�4c"���#"���OF�|�@�DxZw���ц`:��xI$�Y:&�\��4G%�Q�(OH���O(���O<���<��g��[pB@�\�`4��{�NlZ���'"H%8��4��탑�i͂I�5g	A�:%3�O#VU���4�?��i���'�'?O�ӻ>=:E"�N[�yK�A����7��O����Oz�O�V�\��	�N���cI�D�U&�������ش�?*O���<�O��d.�	�σ|]��O�<��г�	��u�O�yb�'c��'���BŞ&�(}U��"�`Ӡ��Or�&��S����xyR�^�a������7969C�%�5ho 6��<���G�R���|����?��'�~���H6qh�bF�K��z��_��M�+O���O8㟰�Ig?�`Fo�H��3�Pq���	F��=���6 ���ӟ���矔$?a��OV��gӼ,4,��$��%���(�O����O2�O���|�����x�U�V��0XX�t���
�^�<a���?���O�Oc��'�?q���.2-Q��:s��]s��.z���'���˟ԗ����'�e� I��D� zB�큱�҅'\�1lZ��Bψ�I�����6�$�O
����@A��Zq���̵Y$<d�i���ȟ��	�����s�S��Xvi.8!�K�.}��ه���ֆ6��X[���Or0mZ��X�I���I���1l.ޔbū �F�����㔫	C��]�8�����J|r,������i�f�c��ݼ~�t���[��J�4�?a�i���'���'��듺��	w�!��^�O�� ���DEo�-%$����|�'��|��vl�(ya*D�aA��9rP�׵i�'�B�'�����O8�Ɂ
z����^p¨ѕ�=@��'/�	�/��I!z�D�Sҟ���ݟ�Y�F�'�1�gV5"����!ԙ�M[��?I�V���'��Y���i���ʽV����L�#u�A�Eκ>��E�<i��]�<����?�����Ӥ{\ ����O��l�a	�aPv7��`}�Y����my��'��'G�lʧ�`���j��/h(1�2��y�IP�p��'�R�'e��Z>-��O�$$eL>n�ؠ�%>J촸ڴ��d�O��?��?Ѥa��<2�܄��S�Y�u�����`T*u�0�s��?q���?���ʧ��ǟ��Y���w	�$M+F�jb%`�f6m�O˓�?)��?q7(I�<����~�̙�CB�)�d6���(�-%�Ms��?Q5�L�<i�Q�����I�v�v�����).PQ˳$��b��x�OL���OV��A�)�$4�D�?�`���b̤0Ӵ��,�R�s�!o�D	z�3O�Ăʦ�I�4�I���K�O�nC�bK��h _=K��i��8?o�F�'O����<�,�A"g��e��)~L,��K:w�\@b�i�"�oӜ���O�$�Ot��'��	*0G��6@3pHdT�ō�6H�8e�ߴTc8��?�.O��'HF��'�?���9���j&Fk��ĺ���$����'�b�'�˾>i.O,�D��\8�fL�)3r	r��<�İCm~��ʓ�?Ƀ)��<����<���?��5c�X�o�&}W`��,K�:���遾i��'l�듚�d�O���?��{d�;����I�Ȃ�^;����'D��Y�'$�K�'���'k�~� >���J� ���cF�@�)�:��g�i�\����O�˓�?���?!'$̑Z�戈U�H��[1m�[ ��%�p�����?����?��'�����|�"�ɱ�
��r
f�<#'F���'��P��	��@�ɞg	,������ҌG[�`P#��+Q3��C�d�OZ�$�O�D��.�8m�O""l�h������#�Ԑxt*���7��O���?���?�b�EY~��Me&�D�|�sr�(;8��&�����ID�R�x���I���)�O:���O�((w�[/��k��<Un�P5�%�������TbTK+�������� ���;�l5��)��M�f���<Q��x��V�'�2�'���6?�U#�L\Dx7B�5Md��U�⦡��˟T����ݟ�$�̗O�� Q޴6��PU��E-6�`ԣ(!�n�؟`�ߴ�?��?���O�Ԩ����\�C�}���xքȦ�p�et��&���OW� �'	BH�<M~�Q�Ѓ@*d�Gi���:6�O����O��D�G�IПT��R?���'��A ԵxS6l�(ڦ'��3���@�}����ݟ\���;B�r y@�e�U)V"@�
�4�?��0��O�.��Ǝ����،�%QŤL�Y�n fS���!Ee�8ق����Iʟ��	l�i�+T�������CJf	:��<&��7�IƟ%���	Ɵ(; 
	$�^�q���F����8�
��I�`�T������ß'?���O�v!#ܓ ���b'Bk��j�O����O8�O����O�3���O������%1��[���2�i 1��Q����O��$�O��'>]�����D�%�A��B)숀���*cr�o��$�����D�`��ݟ��O~�r�I&$�⹡Ga�(��1�ռiuR�'
�q[�'�b�~Z��?���T0���M��
t��L�wOB$�s�x��'��/�/��|�ן�9&�~�p�&S5(E��ҺiY>Y�'�B�h�:��O����O��'����C��4�� ��I!޴�?���5&��p�������5���FR�#Ur)aQ�.3(HP1��6�M���]/���'��'�2�%�D�O�	�]8�X�q0�ٙRR�!JΦ)p"�t�$'���O00ii�'EB*�(O@�`���*e���&%+�'�?Y���?���n)�'���'��d���(���%.D��+�0�V�|�_��y���>�yr�'?��'&x��_���}�����%�����	c�Z�d�O 1$������@&��X�,�֐�����n�=�w#�V*b�~�a���f~�H��?����?�I?�)_�e�6���έ S��{�Ec�p�'�H��G�'�dW�\Z
�P��<[cn`�'�"��v�'� k�'���'������u>E[��Ռ�����6�z����t��ʓ�?Q-O���O ���Z�$L�B���Ч���J?�]��+	#x�]�[�b�'��'7�֝T�䀪~���)*X,8�
*s�h�sv�թN�$�p�iFR_�p��Ɵ�I�_�H��|n��bGC��2e�c�	�:�I3�iK��'&�Q��'S��~j���?���;4������mR\ ��@�X��R�\�I����	�n�B����?�`���
Bʥ��%S7�,�(n�\�k�>O��D�ڦ���ɟ���(H�O뎈
L��\���%�F��eD� }���'���yr�|�T>���zӊ���!0[��4�o6+*I���i�R�w�����O*�d�O��'l剨���L�W�|��
�y
�iCڴx�`�ϓ�?I.O@�'��Χ�?a$��<�ʵ�U�i\��-ReX���'�2�'�"c�>�-O�$����E��1l�t{F��o�"��c�n�`�D�<ɒ���<Y�(��|���?)��t*�8䂄�N����A�0H%�Ӹi���'X�����O�ʓ�?��C@V��d�� ^H$���O�nyoZ�8���k�,��ퟠ�	՟��	m�\c۴�
e�F�j\�)�f��u��IPٴ�?���?i���?)M>a��~ �����c���4i0f���M�A�
���̓�?	���?YO~��<��c�l��0u��� "ɪ����T����ߟL$����_�.kBD�G%58t8r�Ů Z�E9O��$�O��d
d�4��I�ODDʔ��Bm~H�����7�n4 ���ܦ=��K�	�8E}��).jɨQ*�3-���T��/�M����?�QN��<�'_�S̟��������D��u��0SH�tA �q����ē�?������Fx2ݟ`�H*ݏNq��B��y��%˒�iw�X �'� p�<���O2���O��'�щ���=��T: �9?n���ݴ�?���)q|DxbY>}Q"oe��̀fo\�l�p�����v}p����i�R�'f�^����yy�^�@��cP���%����~xt�d�1����G;��S:���	���j ��/iWPI���ž}b"4��Z��M{���?����?i�x�_>u��;i�t#�!�͔Xyp��B�.IЎ}ڏ�y"b�9�yr�'P2�'�H舆a �P
b|��-A&u�2�P Iz�:�D�O��K���t'�d�F��U�&��/9��X� IP7�� �PJ��M�<i���?�������3�2)� D�&�ecZ_����i>4Ol��O\�On�$�O�(��Z�>ZF,#��Y no�iY� �(n������O���OD�����'Ĥ����R�zt|!���$P�e�'���'��'���'m�y��O*M3'��.lN���HۤmIH�IfF�<����?q����O��'�?)'� 2u҅"M4�F�HE'5��RƷi���|��'�b�>��'��x��� �*�y4�Օmʜp��4�?���^p�A��?��Q?��	՟����m��=d�V��N�2Ӛ,hK<����?�!N~���i]��6����|�ӄ��S- iT��'S"�'�r�'*T�@ (G7B�+!��	
�T���Z��M�����20+��.}�7�ܬ|�x�S#I\  �̑aw��Y��f�'�"7��O��$�OL���d�l��c�� ��pY���`Э��ᦽk梐[��|�-�~���?�&V�ahl���Bt/��R���t�f�']��'<2R�d�O]2�O�� 6�W�8\hy��3�t��o�u�'���n@���#c�0\���P{#��h���M��v
5*��d�Ѝ@ܲ9z5Ȇ�u{�P� ׄZz"������Y�D���<m��	�ݗt�b��Ɍ4{xBF�
B>�{��˙^���/J:D��Gm;3�� �dN�TN�y��8@��`q���"6fAT`lL��E�U��|p�J�4]tt�G0J���
�ۜ�rv�HT��`B�i���qL�.ic���B��'&�aIp�G�xmPPI�КK��آ��
�P���HQ��ypb��Of����&���0�*^#?P`!�W�>�ED �~<��д�����iy��'�b8���揳06�kf�L�I�6�+k:��qtBV�9.��gZ���x�"ܔm��d��D[��|�i��HQ�u/���(�3<n�q�ǓS�=�	�p�'xE��V�>l�1 !+ݟ1F�芈y�'�&�y�CR	?��P@Ā:AS��2�'R�6�C*���ƤŲwXXtBDiU\s�D�<��J�4U���럤%?=�	�������C�jͤ��vKC�G����	�d*$�ĦZ�t\H�D&"�j���S��W>U
,�4�F�;��������*}r��LBsB��x�X�U�S+�V�!F��/u�b4q��0���'���h��?�����O�\�J�e�,jG���?�8�P�"OZ�ڡH�x���5���V| T�'��#=9Q�T,x�Jӡ1XN����[+%��ٟ �I!�����	����'�b��1�ȴ���e�����g�8P��'3:�F	Q�̘��-�L��ႃ���I�  
d��Ǝ�/q��d���&7�3����0	0��;Qc燃�1�|�D5?����Ο�g�'樸��Q��i+G�H=F��y��'62���O��i��}p�`�>7�.	9�O�`Dzʟ�[�8jwm8q� ��w��(Y5R�iE<vW�&�'���'������I�|zF��25�P���]��\5�̪�*�~@a���'U��i�MH
-���Dc�}�6�R��	�X$�ǟ�|Z����֋�ʉ;pH@$#*&�C6��zu�V1a�R�'ў`�?Y���9W��m�1	��ɓ&_m�<��%�� r8�eœ-E ,s1'�h̓o��	ay�᜜y�v6��O��O0oXF�bR�ԧU�X�˦ML3���d�<9��?)�O�F����FB�(2,B�^�����v&I��	!4��8�"�-#���ԤY�R-�B�j0O��J�jӎ�OH�x��P.�z�Q�L�7�����"O��A,G�N�"��ĊI�llA`�O"mZ�b���d�U�=9�W���c�t�d��M���?iJ~��7��eSt���GC��!6f�"lˊ�#��?�D ��?Ɏy*��I;��ݠ��?A|����ǋ�[=��'�&����	ޅj�L�c�ԛ4����G��4m��	N�S��R�����ωW���1�I�6����@#JqȐL�)�bD�P�{�2��9�HO������ z�h� �=6d@���ئ��I���5A���؟P�	̟�'����f��"���C�w�䁣S�/�dI)@����|��	+Ip��AǄ@![�m���7p�O.͒�L
�����_�u��m)���y���W�B�'�B!�8���,OV�D�8tԌ�`l�%	��9¢E�G��B�	;��H�ï�2 "РbD�߶ys&�����'���M�8<��'��|��P����=&w��R��˦U��ܟ��sy��'x22���DN�w"�I�Ī�B��USA-�'8+!𤆓Ah��`a<)�S�J�<D\j4Ox���A�䁛A�'f���Y� <:��'��<��cR�2mH�ط| v0��'=�����L"���!$$��@��P�y��>��
p����4�?Q�E��H0�ɉ�y��ȑ��h����$�Od��{>u���O0�ON�[R�!R4q`w,��D�fe���'_Z����ߑ>X��cK�)��a�!K܇�p<Y��W͟l'�x�c��$f�������w,)�L,D�d!���M`�t�Sd�����i-����t�? ���Ơ�"�� [��P�)@���b�D�}A��n�՟���M��՟x���;=��Xe��S�
�����<�	vY���	L�S��O��AՉJ�'դ%&M=n�L��Ė>q�ʗE���O�
(0��$j]��yve�(T���J�h��l�O�b��?�e&C5W�VAbA�S�6��yQ�>D�@�s玊$��:�O�\���)>O��Fz��ƄKٶ��G��'��� HJ�l7M�O��$�O��">�����O��<AC.]�Xǆ	,�	R�����'k�s
ϓc�Fl2���9-u���i��
�@�=��@[\x�8it)�<k�%����Z�C�Q̓����)�3�$ ]tX]�QOU�p�m�ݶ!`!�F�<�tI�P�^P�Y�&돀vc�ɡ�HO>er��(i4	��-�L�F1�1i](t7n���4�?����?�-O��D�OB�Ӯ/ضp{�*���ܐ1G��C,ั�,����ɾ#�(a��c	: X��DK�f�Z��\H�����\��(�Ӟk���϶�����O��$�O��D�<Y����'m�]����� Y�P�]�{��0��'�0�pf�
Ʋɡ ��; �X�h�y�K{Ӓ��<q7 �^ۛ6�'�Bʅ~�(���ʎd67��]��\���I�ϧi�4a��[�I8[2�J�/3@ƈ�M�=KD����v�O��Y�^=zS��RCd�.�R��p�'��My���Cg�
��Gh^����N%C����2������Izvj!�҂
)��u���M�&]-ll��KZ�L�i3� Ѩ��'�M� q�����O��$JEX|��!kK�Y���x��)
-����O���/�Orc��g~�R�N[����]�DI�`pkD7��I*�Z"<��D���"κ�A
�T�8���F�dL������
H���ߋI�,��nC�L!�C�}*�Y�s��N{�
tO҉v�axB %�V���9��ؒ-U�IzGm�01��p%�i,B�'�F�8����'Q��'p�	�m��P�ц�:�T<�7��&m� ��<��c�x���!�
-R v���ޮV�x��'�,�:P���"'pT@����Z� �w�-D\c�<�w�Oq��'�d�k����]#Ɲ ��	s?���
�'��(�B��L� �c&��	�O��Gz���&j9����K������҃,T�-��ɦ���ϟ���~y��'3r<�0�`E\�B�8���c�y� MI#�D�N9e*�N_[X0ϜJX�t�wm��XF�B���V�T@7��"��X���7DFrh6GÜȰ<�bO,.���CL��|�n	�勨�����៼��Q���O��ܸ�B�1.� 1K���4+�y�
�'�l-z��L�#
����x<̺�y#�>�-O`��C;O��D�OV9�u��#t^"p���S?(�@���Ohʓ�?�����P�1(b�떂�V~"�B4}��t���\ �XpQV �p<�!�_�9��ݩAF)?��c�7lCUZ���Ҡ�І��M8�iTi�O��D�Oz�Ɏq�@M�U+E���2 �1-���?	���	�=B�`�@�S�%��av����!���-�F�R�*�PU���jm�[�	��P�'��	PMe� �d�O2ʧ�
�DHp���I�1��}	�g���T���?��Ԍ�?a�y*��I8"����`�0��(x����r�>1q��[���O� -O�p ��jю?5xia�~�dգ{���¾R��Z�:t3��
�:�!��W7|�A�C���ez�
G'��Y�ax��=���R�%Q%XJb1 6�Ґlr���i���'�������'��'��	�kW2a�4��(#h,{�Nˑ4�Ƶ�<As��Hx�@��Oۍq;hTbb�S�W��O;�	�4��F�L����gr��,�@C(�zb�09���Oq��'�A�F�@�L���Ps��w7�t��'��`�d�Y��f�m鎀H�O"�Fz��I��?J����NL:a�bl��T8c'!�ԖҢ����C;�H�8ĪܳY!�AT.���4@w�N:@!�D�[��s	����A��9�'$�M�'b�,�ڰ�u�\5IA���	�'���1����G����W>B<�S��� �PZ�K��f�Dh�C�ʾ�	K'"O��1&^l��y�D�$o�TAP"O�-�bOR�T��b����vKd$3�"O����(8�H�P7OPW�٠u"O�Ub�NH�:����^rt%3�'�H*tGּˠ����A�,�v%	�'X�;�iM	FPԳ5�U�#��	�'�6��a�VZ��B抑~����'�d]�4C�^���9G���X� 1��'w>��%nցbƜ�F̊�f�Xi8�'�`0�7o��{x5���0�r���'�T�v(�9�H��`�+>4,d��'�b��g�?oDt0�a�Z0����'Np���ESbdPE�bZ�\A�'LUJ��!hh�)�".�.\�'�Ɲ�rO�:�&ta��,n�F���'_��E��1�Z1��l��:�(�z�'��DRp�O� �
x0��Ɋ"�n]��'o�����^]y�"E�-�����'?0�c&g�(R���J��;�t���'��ӄ��q���jZ<� ���]u�<)���+
5c���|؞��Rq�<)�n�t�����ʊHÌ�Uh�k�<����+Lt܌I6�@��L��w��c�<�3gE�R�y0��& Z��rc�_�<I� ��EQ�_�CB�t��FU�<)��^�n0J�Т� :�!S�P�<	���3o��	����v�F�:Sa�P�<)rˎ�8Q�n��-2���!�c�<��ل'��\Lُ�
@ �a�<I	�2���@��"[�M	���b�<� MF�%E,�����B똧f*T���Z�a�Ҫ~�щ`N)�l���N�>�A��"�.,�&�C'yEf�ȓi
^��bm\;ot.���� '5A�,��4����LʥX�}�bY��t�ظ�ON�i� bl�N|$���^#R�S��Wi��1�N;)K����j�رB!`�PD�UI��I����ȓ�<�ye$ُ�A�+ާ) j��ȓT��h�@��
[T <�,
5��(�ȓi\�t�QJ�]~, !a ���Y�ȓM}�`xBWn�������d����ȓi	(q2��!3<��EP�(H�����a�B���H�D�̗k�"|�ȓ`�Z�(�(߁�����B��r��ȓ7�<����\,j�������\���?B�����
�i��s)�*�9��>D�};WFI<s��c��E��I:L�}�`瘐0e�9B����3L�U�<1�)��Hy�����x�7/�Q�'F2xd��6F�������T�͏{�~B�	��FiB��>Ǟ���CI$P�G(�<;���	�`����FUN2XJ�@[9U�!���o$�����*E
�ס���'M�YW�'��YZ�鐧LA�4*�fN��>���O��y5�@�=M2���ڂ��#��y�� C�rwH�[��\jCFݕ��O]8@˼�лЎ�Z�:.aj��$�� ��\�+3�ybF�%�D�S���9݀Y�3"ĭ��d^�w4�dT�c̩Z���Ǣ0�+�cM�R.L�GώVh!�d	E��U� ��F:er!a�(&W֐R��M5ȸ�����O!xV��@뛶5(:�ڵ`�0"G!��Y�ʹ��C�.t���y�󤌋
�$��S�? ���"ΒeW:q[d�m±9u�'���i��I?��	^�l'�xQ��>|�t���Z�<�[>:����A�����Aظ"<!& 7�e�S�֝S@�هqp�7@', rB��;K��ԌP�v�,���m�t�@��0gˋMqO�nߴS�����C[~`�ىM���a#�j0,B�!"j=�w����3I��r��Ƀ?oHA�P��+l�Z➨�C�A��a2��E�7�<�3��>O� ����V�ޭ�Ɣ7;j�Qa]^*�J�oܠ@�B �տ(�Y�O(�BH�?�:,��$�Qxj'L��mOl��N3ń��'[��$Ľn�5�m����Sn��U+�0�R�{p9�gY�D�
ң�"to D�o�3�0?�$�ψ8����!�>x~���
	r���G�=!������a^�Ao�U����'��4��]3t�i�l��c�� w��sWO�\1p@֜R�\�kf6[-��5��q�d�+���`����(�0,6Z	p�c*Oc��-&"dRp���{�I��'��5��4&4�y��A�'�05jf6O$<�vD9;���;g�	�q��,(Z��͓C�~�q�a��[�̀�m?Y�D8E|��i8HQwMI�-�q�p��/&��b���45W����)�M7���D�Sc���$O�Y��x3 ��\�D�;1.�?�p?��VQ�2Q���,e�ް�	� ��|� L�k�F�6�D����D�FM�hȷJ>(���I6 þT�E�_;G�"�įS(,�R��t$�(���Ue?ғj{b��!���y8��&T����'��u��.8��esP)�'&��쓋��O�=�Z$��Mx�6p��B���8{��A��40$�ق��{��7mߙ\��u1���r�0�g�1���(B�� y?�������ʰ����d��������i��JX����7e`����s�i��c�pQ�	&�Oj*�D/�N]�S��g'8k�ր�azr욓S�����w����)�	JH����^Nl�H�P.����ϡt*���'�A5����V�Cz�� �R ��'�$	����4���b��*�L�M<I���ץN4"#��i��p!  �I�w� J������(�F���*;}bI�S���:��Λ>kV�
/l�I2��S;��nňPp�y"�B-2d|Ȉ�O�r4��,Q�yb*� GΗ�}�m#�I��M��ɍ$L�*J�569�ai��		V�"B�e��9Z�$��H�q� l׷<��Sb�I�,",J�a�_V���;/J@����4�c�!�\�lk
�L�ج�lK3e��(*�Fo(]a�\>⬝r��@J~�*�l��X9��T@�b����OФ��ȗkk�|0u��5�Nii5�I��RqPc�ەq�.�xBʛ�'��yP`���#�^��ȁ)VsN���/�H�1�|�:VI
;��� aPc��EZ��W�#5�����8H��3�ND��:L���S��"Bn�W��L�R���MZa�<1C&"=��b3��'@��P��s� �G�>!�;��) v3�} �	O��XϓE�*��S�^�gp4� ���u������O*��A�U0�^4��&!��m�$�
^LL���Uza6�ζ"ay���;,] j@hO&Y�X,�󡈺�0<�!@!�"��jѼO��|���6\���'�;JT�\"!FM��P�O�2tHK�`�����
MN7n�[嘟LI��xn�³��h�Dcӱ�R/-1��q���Q��%�g)��yr�4�ص!���`�>8!��կyG�'>9#��ŏ9Ǟ(B�M;Rɨ`�yrII�-�N!�`D�L�ZlAƆ���hO�|d
�WN��(��Vې�c���eɶ��'  �=���d�0t$�����;� ��'i�>
��|@2�B�qF�S�50�u�3�]��?�1*Ec�.���I'zc��H^+B�sB�C�5��i>���CM�R��Y�EIu\�9`��h�<�ą]4a;�P@��8nMlpa%d����D��ELH��R���4��)`FJ�">��6Hrޕ��!W� Q�y�)�x��)A�.�O��i��O�]b�a����a��dM����|}RO(+�F��$c�el�@���L��(O�d1��Z�pO\�q.�h"8E��I�"Q@�V(�eF���)�(��k���\(�u�Tvp���eC��R�X�ʁ��.'N�cO9�Ok�$
3'@������,�� �'F�3�dO�eb��S��B�M i�,g������<ͻ�N��c%N&_
	!5C[���Ȅ�x����kF��@1@�F�-`Z�D����L<fe{5!P��@�O�.ˋQ�� #�mݢ�8yF8{�!8w�ܩ"��P�m�����Q�i�ӗa��=%�I��X�r����Ҁ�+�v��'evdSA��k�z�r���iz"�c 7�"���LP�V%��ѩ����OpLC`f_�מ(բ��q�:R �@��}sv��V"`D�&o\#-�������'��}b!
V)r���� ��6t#�
N�{f(T�ԧΏ�qO�p�W��!� 5�����b�1G���� �	��j�=l�B1�Gř9%fH�I�"O�����T�i{�C�?x(�q ,�B�	��������=Q��9�^��צ��&�U�� 1=��"��'���姝����isl��Zh5����n	��'5�h��׳o\	��2t��p�r�٢$�܅(�%��� ���'	���O$�&T1m�TDR`4}� ���ia�Ÿ�j�[��-RD ��L�QH�N�+/���c�����dϊ)Fd��$�D� ri��k��'��2E��CWB�[5͘�v$���{b$,hFAdf����T�!�D]�ݘ�x��Q�5� %ٵ�X�j���ԅ�g/�7C���S�iǎ#٪d̻dx�ء�ڻ���"$��,'���ēr�@��R���;b�A�ǉխE��D�Œ�����p�"�R��q�qO<� @!	W�;y�~Yz��E0���I�r���	���p)��d�%D(�Q8�Hߠ{=^���Ź*�����W ��ę?/t!�� �ʔ1��_��I;C�>	*W�X*>� �p��[G՘�s��B̧P��|q6&��C�l���<���ȓ�2e#��ׇ4��$�b� v��i%BF�n|HG�Yk.�S��yG]I��R��ńW7v�kq�6�y2b�QT�;#�CG��孊�yB-��wʮ�st�L�V�Y��ɽ{���Ц��r����q&ą�x�<�7�ƿ��4�ޥ�tg�;d4[��T�9y�H�)o �e�AFXB�I��I�� �T�a��.Kh4a h��5(0�'Ն�*ƸiR֡�d+Qn���BU�RoWy��# �=L�Ɓ��"OJ	�6C� $< �A������&�i�v�����Mӧ���I�Mcw���4�8�h���=h�T�� L�0�� ��4���b0O^ q$��K,h��@Q�P{xA��"On�Z��]�%�$L��˙Wdpy���J�L���i�:2���1��۩]s�m�O���!��ԓ)NlBB��Dd���׎��n!�d	� ���EЬRG���Q�B;=!�C:a#dlX��Y�CX;c!��>"P0͉&Ĥ^��$)�́�
�!��gBT)5l�:�:<KtO+a�!�\M��bf�G��s���]�!�Ĕ�P���z$#�&m�m���b�!��߷w�Xy��0l��@3G��4�!�DK48M��2���~��=�'�ՌK!��I-L���`��?e��È �T!�d[$�t5�f��F��K�ߗk!�^�l���r�̥-U t��>�!��*�iIb$T�P�1�O�^�!��^1:�4�3�Z3� a�5hA�`�!�D��t�Zw)A�`�8 �����+�!�Y�@�Ti���9��4@���4j�!�D�Q�@���LY��� K�5�!��|�h�e�ݐW��Yq	Y�)z!�L/�D��u��O��m���-$!���
D. A�"/����^�
�!��x�t{Pe�#v:�u�C�G�!�$��4�Ƥ�$���z=R�!�!�Ěi��ФdH0~�Z\(4�Ϩ�!�d�<�M!�*�{��)4�-�!�$[a �y'�Z�f���(���!��Z��A�iP�GGd(�4GX�s�!�ă�.�����X�fG�Li�� 5.�!�$K�^�����׊36=a�g�%�!�."M��'A��/�H��0G�Uz!�$�E�nM��X�d�*�Sg�.E!�D΀Dǆh����?z�Z�x��I�j�!�϶ L�bC1��}#�C�"n�!�ą�M	�:bd�$eM΅��/ޤL�!���Y�lq#���hR�(�I(G}!�dޑ��!�-42�|k�ǎ�^!�d.� �32
St�L��bx�!�y���#"6u<q� (�� �!�� ��o�k�Ќ��#R�Wjαi�"O���$��(q��v"^��-zT"Ot��ƱT4 B�NЛX��̓2"O� �D�5:����)(�d蓖"O�5�2�7b�Fi��dN8�ě4"O���Si�q ���m1�`�"O@x3�D8SnN��R#�	��p"Oh�(D�O�wII^��p=��"OhTɴ��W�,�)�׀�6);�"O�M� ��4Ӹ��R-�M��"O���G�@�Z¼ƠΨv��%�$"O!z�nؿR%�����7���g"O�+YukN�����<,P*'�Y�<�F([�4�ᵌI�)l2�IV�<Y���8��MAmʄr��1��S�<���7]��B@
%�Aq���u�<9$��3 zU;�C!�jd	�c	u�<����r,ъT�;s�49��^t�<IVK�:> z,��^�S�|m�sHHm�<�7��;J�"%Z7a��kp��Z��^�<� ��#Z|���	�]����gc�<Q�n�.|���D�wd��i�<A'����s��ʢ{f����B�d�<�S�ʮ4T<+)*~=! _�<�Ve�)�0����m��وRD�t�<I�bӷ_����&GJ�a_����BXt�<16�ғ�b�GG�M��D"AZX�<Q��;44�Qj�+ܾv�6�I�aQU�<1G"�X� �jCf�8/4�!�`�Q�<�ņ�#(�.�u�L6?#Z!� i�V�<����ߘI�SeM�!R� �M�<��h�r�)W�@ ��J�s�<��OZl�:�qV
���1�jr�<���2g�b]hF�< ��	iW͉d�<Y1jG�d��i�5��2mٴ�I�aAa�<����#@���G��\�!�R�d�<��.@#|c��K"*
�r A�tN�d�<!��́y�$I��ރk	� ����]�<��	YV�xq6�[�u� �~�<Yր6I
H������5���PCev�<����PH��^"!.��'��r�<qTDC�x�� ��R�Rl3F�l�<i���ݤ�2��)(���0�g�<YbOD?V3Ҁ����+
	�=;E�i�<�!�:`8�U�g%ѧ<^0mz6�Va�<ysMO�(
YC�� �D�]�<�C,�ʩs6��" 1h#�HW�<q3�	�qRx2č�c����Dd�k�<�ޅ]̀a�@m���2���Mf�<�U �?+��[FHC�\�8숷�`�<���'�80����+x�lYrvK�A�<�V�"
mЙ�7Ǟ%M�\k%�AV�<Q2��-[Հ�û6��	�e��R�<�F�Y�.!�`M�5X����LO�<A�+(8�0쫱��W����<T��q�ļ.�`�F�"=eTԊǂ(D�4��)A��i3/	�| ��Fe+D�H�V	5jr0�+$F�Mj�a�5D�(xb	9)��h�@��yjs/D��0�׈|�����>x�< �+D�$�5j��\f�tI�J>Z��h��E<D���4bߕw�@I���D�#�:D�0��A�{�"�(Ab�T���CQ�-D�@��F�v�3��O�	*���!)D�� ��*��uh��@5Gx�<�y�"Od��!����)Q��-S�8��E"O���ł���Lp��Ġ
�v���"OT�+���>�H�f�T#G�ؼ��"O2b���/X��`�$��3sH]��"Orh��]� ��äh�	$fiH�"O��h�&�'D�� �&ha:��"O������:
(`�R%9X��qU"O���G��b�N���-j>�d!P"O ms���.#���`�H EFJ���"O����7���r�9��1� "O`-z��[:(F�<{�d�!�R�;�"O�,ђ&�#;� �QS!�3l���x�"OL���lQ�R�a#fU�>0{���n�O`���iH�Pwf�K�e�4Z0����' V@�W�ܥ1hL�i�@�fy
�'�v�x`(�x��1��Ȝ�7���A�'��Y�g�8)X`���%������$5<O�ᠧI�,�Q7�o��͒&�i�ў"~n�<�ЂCo`}��̞1<B���j�K�ih ����3�VB�I�k
�R���"7 *YzC�I��z�;�Z���U��B�	�UP� ��"�?YݮM��cO�|	,B䉊Sz�j�B7J�9Q�LL"q��B��)� uh��Ǉp��\�$ V�>�B�	�4պ�N��j��u"�7]jB䉾Fy4=:B⑛.>u9v�ؒh�jB�	;vGB�)W�*a#&M��(��Q�DB��#+ 
�x�ۂ]�x���Դ@6B�ɿC�PQs��R�T �	P��c�tB��"
"h�סZ"]H:r�R9 �.C�I,=ג��e��Og�D[vio�C�)g����bU5]�����M�B�ɻ*Ӝ�d�4	�, !�-J1'W�B�
9L �a��j�.بW��"FXB��/#������Ϩwmލ9a�g�2B�ɓ)0ĵ�	��{]�Y�I	4]�B�ɲ'84��O�z��)�ƕ&�B䉠!�4t�a��!9a<@���@�C䉰���iP���`��
(��;��C�0f�d1��
W�Qp`n_N��C�I�4��C ��"w��E�"7��C�I�$FX���+�.w��w/ۤ&�nC�	�T� �� K�7[��!��&\\�C䉙>@H����;�q����C�<b�L��-� �FD�&HҿǰC��<L"�1�ݘq6Fp���Ny!tC�	0 �[4d?�~�����rC�ɼɺ���_4Y^=�U�)2Z�B�ɰx��܋A�!k�v%#t�J*ŘB䉩n
�hb�I�6|U���(7XB�	�x� P��G��eq.mY��S�zC�	�z���ǣH>Hh���X����6������a� e����᎐;т$�ȓ>2�K	"+��L�33p���S��)����;���Ə7LaL���:I85TbK�����K	V�`Є�� �΂�>E�ghZz0�Ʉȓ\��dX��\=�,�¡DZ�Pٖ���yGR�H�+��~W�Eq�R�\j�Q�ȓ_��1P��7�za�ɜ.�P�ȓ#8n�����qV�� �S�H����<�G��9�n)�"�ۧ'zu��S�? .�Ɂ"'ਙP�H0~�*��w8O�=E�4���"�  8�I&n�Vda���y���)+�iH�#��im:�C������"�O�m�'ʅ,y��|R3jW
c+��ʖ�'��#<��BU)#�-"D�'�H��1��a�<Qc�*M���bg���Ԍ����]�'{Q?�q�$ĚN����Ȕo��c��-D��P�ě"w��G,LI�YI� -D�2Fg��ɞ]bt�E�	���@GL%4�����S\]���3e��y��Om�<S+�k򼹤߈
W��
��]�<97�ĩ��͒���	*���bAS[�<�����^��`!� H�s�Z�	�F[Y�<�gI51�ʌ*B�� _�flyvKNV�<q�%
b�4S��:_>H1��n�<��,��h����(�F��@��g�<�p	_-E48=�c�M�P���GK��!��� .�x5Ȳ���+T���V&�!��,�eqW��Xp0xXČ�9s�!�дTQV-�f��%Z�43��,e���hO���4/έ82I%��)��y��"O�	�G�+^�ذ2bC��a"O�5�fD�v���*��ZĚ��$鉤e��?q�L#[�!��R�l�x�I�` D���vaY7h�vek�"��K�@�@��O�Y�����24a8U��[���)��OG�8?�y����@�G��_������;5����'��}�F�7^��ܣל����N��y�V!f��A�AcB�ېAsE��*�yR��!w�6���M8ŖX��Ǟ1�yb�#d�FI�`薱Z���yB07��d�D.M����L���y���a%6��b�{���eE�.�y�άn��Iʅ 7��|0&�&�y��Bۼ00p�2�.��d,��y҅S"~ִ,�gڽ1�&1r��P��y�m��k�dUٵ	�'���;�V��y^�H��yy�U�$��h� �y����_�_ .�q၇� ͚1[�'� �uE֥bT�E[��A4����'��E�7��0��]�dS�6(��Y�'�e���&(�4�q�65��U�	�'N��{B��*WD%g&A<KC��7�"  ���{�0)�6�نQ��B�I<HQ� 2�	
���"4��B䉉b��K���p$��0Y���B���εS�,d�]���A�;_�B�I
W���
'X�RM�,0���Z��B�I�|�}XA�t��P���A�*B�-	7�p�!!Uz
`����.O�B�	�v���iŬ	� ��qSaJ(nB�I&���QjG��� �4F̦B䉫ך�V��:J	��0�@V-l�,B�	�=o�]��N���m�JO��B�I9/��������T! ��C�;"غ���Ȃ�q����l���C�I>�|`�*K��K��3f~tC�GŐ離̍z���[Q��M�ZC�+$��QU�H�m	`=T�BNJC䉑q�>-�ѫ�/�`؀S��X C䉄����\
�s!�̰b��B�ɹ ����<"���5e�7)L�B�I�:)�AY!H͵R
��ҬɃ[|B�I�,:��%%nI��Fț�bB�)� 2� �#A��P��l)W�m�s"OT�P��+*n0��jT}p��e"O�LaA��<����aI�Hmc"O��{T���u��dhB��[J��Q�"OH9��-Ђ ����`hķn.��aq"O�1W/ߍQ}�)�2xqd"O��s&��$4%�q�� ٨Bu�՛"OP�����X�O3]=�!�b"O�ՊW�Hz������4L�"O^x �Gǘ��S�DA�\��	D"OHȢ��
XM�i��3h�$"Od`
�+̓O:并�R*nWvD��"O���4�
�G��Q'�ҐMA�@Qt"O�����;Q`�(E�&|�%"O^�*R��4|pb�ص-\�s�RQ+�"O�IY%Vg5@��"o�P����"O�T�B.� TÖ��pD��|I�T"O*�J�H]�
0�Y�CH��<��"O�`�fʴl��͹shBa��%@�"Oz���ʄ!U�z�z�&7���ɦ"OR����B��j��٭1�vm�a"O�p2�	�0�<- �E�~�^xW"O��3�#/A�iCJ�%Hȣ�"O�0[��j����h�u�p�Je"O΀��Kz_<t1E��Pv�is"O.�V����A$.V�=�l1!"O<����;Q }��k�d"O,!��D�'x<+E��`��8�"O����9T��5��N֒)x!�"O�5�c�X1�\�w-�"w Fa�4"O� 1 D�-.�� M��6��|��"O�Aa��R 8Z�
6�q��"O\��BGǥ9ʥ�U`�$"�I�A"O�X�1G�bn����h"��"O�m���W�x��k!��kfܩ��'Hda�׈ݷle�L�Q,�91�̱��'�9H�N�-*_�P�ƃ�(�:H��'�T�6�§ �j%2s�O>#��Y�	�'��A��³K�dX[����غ�'NX8��C7\�"���ͅ���mx�'>����#�<AѠ�$�QY�'����O�k�UALDz2x��'�p�#�H�d$�S�O��}2�'������h�>���R.(�a �'  � ��SN�s�Q�yHZ� 	�'��7c�#jenI�RN
�tۦ��'IvD�%�9JZ0�j�#.	�'x�]��%��f��G% �&y��'>r����A�qyh��U�9-�9��',ܻ��'QS�`�"��#��X��'XTQ��GS�5���D�M� tY�'����r6�R�JRL 'K����'�*�(�NB�6q[��E�xK^T�	�'�-�'@@=V�ç��<kϢ���'jB���F�~p�E���đd�F��'���H��|�̠C$�@�o`��h�'[T8�0��;$4|ы����1Z�'AT35��.���I�e����@�
�'P=��3C2șH��5
MV�
�'A|�`��̆i2�)xЬZ��2���'Ċ)iBBP�v�ч���\�}��'.0|q�A�"�6�	�A� zql�'�&M�v�ҥ{�����y�Pr�'��5z�r59F���v������� �Lbb��%X&���<�t��"O�K�n�p����9d.��
�"OT��®ެf�j��E��3fBYH"O�!rN*o�F�2�N�DSzA�"Ox+�,��r�Ґ���
 C4e�c"O�����W0a�
<!E#[�$&�4��"O\`��O�C	��g��JLp0"O�%Q ��Z��ibVa���|�a"O��0҃�VE@����ʶ�j�J�"O���⣀F��1�b��!H��H�"OZ#��Ȳb��b��#a4qj�"Of�b�72vQ1�HGȀq"OV� C�1Ț �w�X� @�Y��'L�|rQ!M���M�c���
�'9��J�k>2p�����ZƠ�'� -��<jG�]���QN���C�'�,��>e�"�	��ӌFp��	�'��	��L� '"����/��>��͠
�'�Z(v+V�N&�a�c�4m��
�'����g�,<F��$��;b0����'`��h��*@.���[�1��(	�'N���	��0����R�G��	�'��t���u�r!��$9.��0	�'�H}"��)�L�`��Ρ4bތ��'h��e�N�H٪T����-dQ��'T*��T ��
�!qG&�"�����',����[�`.�ٓ��E�8lZ
�'F60S�	
�A1�ԡ�ԈDZ.��	�'��]�5f�"�@B�חl��5��'���ba�?*����MN��@  �'��@�r��>nF,S��N7����'�����!@nּbsn��VX�	�'9R���ₗ3��ZS`�>�2���'sf�{5���i8��Is�TuPl�
�'�������\����`�T�	�'�` �!g�*;�
a�jY�R���	�'�
m�$A�l�l�j�ʌ/ք���'��4[t�ҹ`z�9����*0H��'��ұ��9%e^�+qJ���l��'��P�Q��܃�c��V ����'5���Q���=֊x����"S����'���I���B�nB�;�<��'!`�ģ�T�跥W4�܁��'����/Ղ��8H$�Z��(��'�(�v�
�ΉѦB�$|$��i�'�V�yBC���R�16,�y�H�s�'�p)y4F�6ew�3$Q&n��*	�'�0�@F�S+6e8T�S���pG*Lz�'�rU�enն>A����懐u����'�f9�l��
�4,#�-�^μ�	�'Jv��`c��(�`�:�d��3�'��န�4�!b㋫og�d`�'|�1@j��y[�8{q 
�����'^r�`�2wj72�V] !����y���1X�d%����A�L�I���/�y��8)!w��4p*�V�8�y�L-t,��,6�e:H��y"D�02A@��W� XV9b�k�?�y�T*��r��M<|��@�0G��ybL��l.���"y|��c`���y₀3@�m!�ʧl .5���S"�y���.~S`�ˤn	�_�4%R�A��y�[S�D)s)�*U-�$2�H��y�D�*�0M��S��ܡ��Z9�y
� D��kRi9v j�/�[���2c"O>D�v�S	=�:�ʐ��4��"O�����J� m�@���Q�m�d�"O�P��I2-��1%e�$UŪu�"OX���b:�����2-GT��"O�͢U"�=u���+!H0E�p�g"O��`�
Ԕ "�����"O�9"���E���:��(�V᠁"O[�U�F�v�B�h劓9`8��@"O�8	ڎ���	U�#4�M�f"O�pЯ�y7�]��(W�F�sB"Of��%Iٗ:�ش�SŃ�shI8�"Oѡ��-h(A�$��S%^93"O�kU�I/6�98�mXvD�
V"O ���m�=��H�C�&�t���"O�	vH��y� ��G �u�D�G"Onx ���7�t[-I�jp�ۇ"O��$�_Y���I�F[�( �"O8�d�������7�v�@ ��"Or0��B:~�PqU)��c�J�r'"O���4�O�����ˆ?l-S�"O�M��cԴ~}��
���# �ʸ�"O� 3AÖn�N��� �P�
 p�"O��Vk������Q'�9�t��"O�K��̿9z�)�k!NX�l�Q"O�b�� g=vJ���U�1�"O2��QB�J,cTD
..��	�q"O�|����-ur�l�P��X�ux2"O樂a�ޥb�h�ӣ�5dH���`"O�1a/C�$i�y �BE�C�P��4"O��S�"�
+��3��ДO�|X�"O���A�إa���is�
�G�j9��"Ob���1O=���.^�[t����"O�+�
�[9*�a��6��-�"O�&N�M�VM+�,J7F^�ś�"O ���
��U! ����P�=���"O�����;%��;�c��.��u6"OLԍ�>l=v���#���~�YT"OJr҃B�{Bn���O�[�\� "OJ��U(��?s�����ld�"O���@NKĂ<�u��	hM�#"O��p���e2�EV�_����"O��s���9�B����#@t�"OhU"�lA����7ꁡo�*��E"O�PP�ʕ�.�!E�Ew�9#f"O��PG���V���Dآ�r�Z%"O칐`��\;eˀdl�̫#"O(@�� �*A�mR�bǧSb��iD"O`�B�5��	��_8`O���"O�ॆ@	n�5K��f�N��"O��x�L!#Ǫ	&��"�6@"OZa��.ͽ �iC�gU�E�*��6"OL�:�B�0ay�s,������"OT%8%�	�u���Q�WD�z&"O~����<f��k�䌭P:�"O�A��D�<�Paz�O�e(���"OZx`$���l�@�K��H�T�3"O�i��8� )��b�*c�b8C�"O��Ѓ(O�2�X���[�x�r�)a"Ov��7&U!6@�3"�FV�~��a"O�|HjQ.����G8W�xܳ�"O�����X~"�q��٘w�X��"O��s a�J��tjc^k�N98a"O0���c�)x?`;1ኰ%��<��"O� T��T�C�7$�"�/RG�*ܫ�"OV��g��@��zP�3��i�"O���x��X�P�tu0��"O�Q�!ON.9Q�BG86ь�{�'[�H,s��L��@�4���'`ș��aK�Y��ʒ$A��j(*	�'4�`*��_o�l�Qw&���z�)	�'��X����j8�a�1+@8a>~���',ୀM58���k�nI�\�& �'"�����D5�����	�~���'���ѦL
}!�P��
L���	�'D��\w� ٘b���m~`A8�'��A	�Ǜ7p�F�1��{�l��'O:4�����8j��ޤx!^Xh�')�ۤ#]�SK���5ɾ�P�'Y�aa�	=n�×	kJX���)��`X�M�\l��.^�DS��y"������	��C�,��W��y����]:���SZ0����5K��yb��]P���FBˆ=��0ֈ%�y�.�6@�D�Y���9*(�425�Q��yF�;|ud��Pщ'a��B\��y�Q	\|�:� ���P�船�!�d��L���eK߬�8t�wb[>����%F�s��NH�4�uD���ya�G0(���&�5JG�y��?$h�H���4 ������й�y"/�9j�SE�	�K6���ՋR0�y��7J�@;6#G09݂i�Do��y��A#y�		�d\�4G|,�����y��-0��AS5₇5O.5����yR$�2����$E�A��!b�nT��y�va��i�͐�16�lkG�M�y�C�(���bM�0����FIѲ�yb���]�;p���&:Fi�V!���yb�޵��S�B���pp�4�y	�4�(-To���v���]	��D�<����'r�I<3�<�2!ޏR�<ig�?^��C��1@޼��1��/@��8���3b��C�	�1��8"F3$�N܃
G�Y��B�	�W_�D��E�xj24)�i��4�vB�	�@�<�ɶ�G�^�0�(&K%��C�	�wl�u����Of-�f�JF��C䉭V�����4Zj�* 		\�C�I�'��%{�j�oPA���ƲcthB�	�\%q��֑2�W�R�I
�B�	�V?���dԬF:X2v�N���B�	�H�,�
�	��x2E�>'D�B䉓$�&-�� �t�Jy��"
m��C�i%�2��-g�^ 2G R���
�'d �Q�	W�*ξ$#W�И<�#�'�@e�0�U�(Ҍ�����(����ȓMV qaǄSE����_\J8q�ȓ��9qծ�<���q��I:R��ȓ/C�ݚQ��lr�k��̇�R=�ȓ>��
�C����=;���>�� ����-ҥ�£_��e��D���e�l�r�:O�iw�׎V���&�\��	<z`l��J-}(@�4��_v6C�	/?�~��cýq9D��B�Z�"pB�I<�Y�Ǆ�#�<�8q#U�-�xB�I)Y}�\z�j�*���C��`B�Ɇ���(�0:C�l!�͊2.B�	 ��ʓ�g�r�	 Oς-�C�)� f}�ף�U�|L"(�f����"O�؋��"F�ŉ�$L:|�Q��"OD�sC��X���yC�5C��1��"O���w�E(k���6�� b�N@��"O��ЖΘ�}�Ƙ���d�aU"Ov��*F)��[��.+f� �"O,�3͆2RH�p���2ֈI�"O�=�� &"�I��-�p#��[��|�'x�Oq�F�Wǝ�%ox�Y��ܬ�"O����JK�z���P@�%*��z�"O,���$�^Ԙ�:�o�4֡�R"O*��A��.���{�N`I�"O����m�$,���
���:(��+c"O:���	ԗ2�z@��,ϻS���`"O��;����l~�D��nN�r�����p��B6�Q�y�ڍZ�֊��P%x�!�$%S����p �3V���kV�*�!���tC��#G(���hp�K7H�!�DA#"_̰&�R�i0���<3!�$L,V�z�k ���)Bi�����u{Qk�)���g��aw�ȓ"O2,��%���*�����M�I{���������
h2R�٢�H,G����-D� RU��^Ă�C�dE.27�����-D�$�e�R	󀍂e�>f�3� D�䣖�.
(L�� ��~�@|j�h?D���0�R�dGr���)Ih���<D�|�&kÑ'�h�r��$#�|���:D��&���QߘU��ҿBS`)�'�8D���u��:c��sOքY�8�2v+D�0��T2"��D�wDӆ"���Q�!)D�����؂$��,8�3r�����;D�L��(�z>�� �X$rF��X&@-D��zf��K�����Y'~(rMbR+)D��`���%uRp�!�<+�6���	&D��S�==�M+d�W�Q3��."D�"`�K�C�� #F3S������>D�`Agʈ�z�ƣ�*r��pS9D�(��>o�8Pb)&Q�	0%1D�DP��(^Ʈ�"ro�P�����C9D�`x�ń�J�Js ]�wbn�a�$7D�h{����1�a���^�6d�S��:D�H��� }Ͷ�q�gZ�'�,�y�o�O�C�ɾ]��ak6��9<ۼ�����9+�XC䉁4��yt�z�ٸ���)$`B�'rn�H$
݃G�:����WBB��-9� @�%��>uN����Ik'
B�ɬy}`��Ĉ^��Ri	�h�C�ɈR��0f
�$�T��"C�&cRC�ɥ+/�ڀ��Z���)A�^@rB�I?{l����U���- "n�B�	蒑��+.�&Y�#�4W�F̐"Ob��)�"7�&<RdA@�6��-	"OĨ3)
�vh<����#-o
(s"O�	T+'�9��K@ND[�"O (�dؽe�(�9�('el�&"O�;�`��:�ּ�'�'z��l�P"OL���L�~��y�&�$l�j�:�"OD[��Ag��Dң��+n
��W"O,���i�o�Q�d @�%����&"O��;ԣK����=e�F�8T"O: ��T�y���œ?p�`"O�(;�M(a��j� @��"��"��`�Oh�����"�#��Z�!�mc��� 8a8W ��_�����'�-"O�C�d��c�Y�#�в_&�q�""OPA��2bEP�,�;fp>��"O���E�K0.�Șa�ch�A �"O8�"���� �j��f�\��"O�)�˅ k" )�b@�^�HI��'�ў"~��-т�9P����|,��B��yR@G�I+��Vj�)j�.>פІȓ(T�qE���mJ����J3*����`�d,~=�h�MA�7Ū܇�g�j��t]{\\駬G�n�T��>�ȲЬ�"Tf�0��� ����ȓU���&���;���|!�d�Iy2�)ʧ'��axŦK(X8�JD�Ó=V����l�h1kC���x&��� �|8��ȓbH<�rN @'� i�J�L8栄ȓ/
~�+�cU�|)����Rqh�ȓn׺���eT�bc�Q�I5X���~g�1�.�ș��L�?I:t4�ȓ6�&m��2FN܊�*��N�콰���.�	d~�튡rQ~��/P��
ǥթ�yB₴r��#�P��a#���y2j�bd��D�3��9�$E:�y� �	\�� ��.B���+��>��O��w$�p
��ƪ�0Pͫ�"Ox�t$|��#Hx�����kr!�D=vbSk;��9�b�%:���zybT�4E{bg	�C��㴣Ύ}KD�����!��R�6�"E����%Aư��K�a!�'�Ub�Q�:͘���
Ac!�Fq��e�2e��`���|]!�d�3������
4\�q�pk͟5;!��'�tP@���R���"�LY<!��#@�0@Ӯ�@/����+�2R!�Ę7w������EIȬ���'�!�ۃ���ɲ��_Xd��$�39�!�dM�f�y,P;FK��HD�{c!�նD���:�HK
3��q�knL!��B] >���e��5�4��;p5!��G&tZ�8�W$/4�F$���3t!�D� 	�@Hw	�����g�[�J�!�� l�-�#��s�A��B��j�!���vDD�*��Y������q�!���Қy�'F��B�M0�H�=�!�D�3-�&#����W���_�!��b����w�L�^5�(�:!�	�#��xXA��!U����*�A�!�$^2|}Dؘ��H�ctp�5��^�!�Iq�$�%J�����K�ae"Ov�P�����4�G�ro`䪦"O���A�X�a^�js�Ƣ��qy0"ORQ��а����,/�� ��"OjhB# �( Bl,�CN��A�H�"O*p�ϡLU��80n"+�VŠ"O�<�P&B�#`��j�͖���y�	��

^��'JF�e!F�� N��y�%ܯ3 �8J�GF(d���*`NX4�yrj�6�������>Y��T!�@K��yr�&.�=���YU�0�gN�&�yr������P7�T�4�D�y��`<�� C��zB%�cfT��yңA`&δ��,P
s�XQ�0CQ�y�n�RϠ�"vo]$Ơ�X�d���y-D�C����e{a�]��dJ�y
� `�B�\�0�:!r�n�M�y#e"O*��6���d��(B?��R�"O���!�0;nL���g5x�ȓf�T)�"H�Yw���Q m �y��g|��C%)��)䜪a��xP�����ܟ���� ��i�ĥ֚4ޘ�!`��N�<!5c-/\�9#c�7�84	��H�<�g��F��8��.6O�A�%�|�<I��ϝ����c�+pf֘�
x�<�s
h�dnn�D�a!u�<j+�8@��.� j�d%� ��Z�<1���X�7�S�b��\�$�_�<�b`J�h8"��wK�� ��53�f�B�<�f�!G�U�k��1�� Á�{�<�"�tlT�%�׌-£�{�<A�n��D��1�Hu�4��1)�O�<i��-�X��R��)��fdM�<QuaM��j�l�R"�S1�BF�<i`�,~��VኗoĞYibb�'�ax!��`a�ĦD�"����aO��?��'�����%|��a�fɂc\<=c�'�
��� �ʁR�^ǂ��
�'֡y���R�&%+&O
�l�@�	�'4>p`��Ґ)y��V��2|��0�'����IJ�z�d �5ƨx�$*�'�`��>%��$���A�mW��(M>�	�'w
�����n�����Lهȓ6��L�M�&j� Hs$!��%�ȓk��,9�o��^Wh�ā\a�8���Q����C)�:X��		%+Z�$��@r�I�!�^�PQ��ӱ���rA$���~�"��'S>�J�#�!J$Tf���z���둚NeJe�S�O����IQ�'�L��7-�)�!!T튰#�F���'��� a�+�ҹY������L8�'C<)c��_2p02�B\�����
�'y`�Kv�p�B��b!�'D�4��MŪFrr 2�j�+��
�'Iz�R��N�K�l�k2�X�
�Bt;
�'��e(���9=ل8�$ҁ���ߓ�'�HȨf�1	�Xa���cM���'�aA�Õ?��0u�ғ.��`b�'>F�8��/ �l �D\(9͋
�'�J�	�3=�^d��e&�
��	�'��H#$�ݏ7޺��'�#���	�'k�9XV��9:��s$�W�F���b	�'�4(�fk�1uwf9pM�8����'�jQZ7��;(�B�(B9` |�j�'��`�Wk;�غqFǂQ��
�'������(�l� A�ǳv��8��'AT��0���l*0AB�}^e��'�����D�2��
��)<�!��'���w�	-g�|p�g������i�'Ypm1�$�= >�\�"@��:���'L�	��K��m�:���R�v>l`�'�dt�d�_��2kA�@;kfά[�'�6bF#+6� �E �=����~>�0�lS�o��b�ȃdb�ȓ6ȼ���h�l��4�����D�@���^E����`��Y�1�+޾bX�h�ȓq��C�R0`�~�c�͔�T��H�'�"�)�ӚY���ap�ުXb�ٛ�fQ5���0��z5`�%� 	���
�UH<D��a7�S1��,0ӥ-!�@�R!�'D�� �q��׶5s
��F�D�A~� �D"O�(B7��٘9{�%�]m���"O
u�E��+s ����=A����"OA���i�d���̌�U�0���'�� �a�O�mN�٣��BM�qc�,D��֭]5wrș�e�L���e$&D�0P!&��	
b5�WDہi�lB4M#D�����23{0��I�1��x�T�?��Ԉ���c��9F�*qK��_%N\����"O�dA4OA�_��� �i�FEnш�"O�A0V�3�Uz���,45��zWX�4��`�S�O(p��|�p	�:"����'ɂ�SdE�{�y���k{ �+�'��"U���Z��r�^�H�x�',ܩI#H
"4l��p�ͻ�+
ϓ�O��i��4d>�p�V+=(�� ��"O�S��<T���k�)L�:��tP�"O���������jVnԚ�bXY�"O��R���9���q��;(W�Lٴ"O8���O�Y�ZY�c��"C�F�J�"O�p��h��>!⫀Z����"Ol1���6[˶�����<C����q"O�mЫX��]ү�7P�Yd"O���
	��5N�D��u�!"O�`WE�ϒ���y���b�.�y��P$>
�+w�P7#�Ipb)!�yB���XX�`�����b���IE �yd��H���ɣA�3��53a�W��hO���dT"26(��`AB1̀C�^�!�ȖA+�L�-� _vMJP��%/�!�DO]��8�b
P;H�^P W	�+>�!�$'F���g�+G7z���ˢT�џ�D���m"�as�&�9�ެ�v�X��y,^��fΉ�H!bD��y�M�/;�ش��l�h������y"��$UG�(�7�ltF� ���2�yҡ��]lA�VgǨ`ZL����3�yR�ҙ5$��&FC8f]z��2ş�y�j�/nl0;ŦسbX ��½�hOD˓������jT��D�G2ٸ�"O Q	AEO�,�K@,�;�8��2"Oz�cB�*uv��	�Q��1Z�"O^�	��c��yS���Q��!q"O��@��!�x' �O�<��"Opu!ǒ��t`{r��([/>uKD"O�d��O�8_5ҝ��A�H��@ht�	�X�	V�O`(�4�N�%��W�9o����'��(�!/ XЁ��I��\�$���'L%��.Vx����B�� Sz*$s��hO�6�
�4���޳a	�]hT��?#❇�8(BU��Cȕ>���h3j>3�(�ȓV���Qe��~�vL+��	�x$�ȇȓ<��M�>ƒP3c��W�($�ȓ,e^���1 =q�@Z�8�1��@H~XɌ�c��0�&�^�jtR4��7b����X�<P�HU�D�p�G��S�{K����A�m���`��C䉪!�t�D��-i��n�7��C䉓3����� ��k�@�:=��C�	QG����-�jn���OY�ҦC�sp�@��-5�]��X?�C�		+����"@��I�0��O "C�I�hj�B�-�,�����5&a��=iÓ���fЉD��<!uL�  ���S�? b���&^����b�N�p{��v"O �Qf��jG�A#�↣`lN���"O�)�&ާ�<������Y���"O�|" AE;a������;U���@"O���d�.V�Mj&-�K>�px�"O&�����]d� ��1|;�)z�"Or5�ՊVl�P�FJ��
L��"O�E�T��^��0�+_v�ź�"O��$*!��h�A�=0��{�"O��C
�]n�)�Em^	m!�� �"O@H���<Kw-�J��Ey��c"O�,ᐦU�[�4ti$��3B��H��"O|�G�V�GļDB�!��3�"�c�"O$�	B-�"C��
!��2t��$"OZ8S��)s~�<r�!�s�f2�"Ou@W%� f�^�B���*2}�e"OL���I�CFլ8x
�W(��B䉡��ە�I�t0��80B<��B�	�;���1��Dt�����X�T��ds��YK��t���MșO����M3D�̑��ҟp��K�ǀ	c<%H�=D� !d���I'^�;Tņ2>q�Cc/D� ��`W:)^��:&��i���)��:D�칇�lk�ǫ̻`�����:D���v��Izڭa]�N��;�8D�<
��Y<{��Q�����P#�f4D��³�ӗ_�,�"�M؅euTHG %�?�Sܧ�D%��P��C���	o�d͇�.��]����,D2�2#c�U�ȓFt�3�K��ڟL1��ȓ��[���6�,:T�D�� ���I{�'�윫�X��0�
U�p�~Ի
�'S���М&�P%�D�^8c����	�'	HH���k@�@�d��j�~M#�'l�8�d�Q�0|���+j��R�"O\(��aF-��I�蔵.��pz�"O��Qˆ"h�4��3�\�`��y"O8ՠvdϓ,݀��1N�/}c
��g�'k�OR�?]�OG�Zamͺ"��*����}Dz1x�"O45��(c�z��@�4��aZ�"O��f��/����t*\d��dE�'�ў"~2Ï�G�"����.S���&-�:�y�h�a�����Ըi4H)��L�yr�H
��{�9 �Q�J��y��_0GG���bI5t�NY�p `���Pov|Q��<\��R�δ��ȓR�$�c�-{��qг̀4{�\���ff�<�֢��pB&$�T�.Fj���Il~Bm�1K`�B�	�zbXt���y2
ʍ(tpR���l��@��EX%�y���B����G�,g���S��Ҡ�y҅R/���r&�^ڑ�
�yOO�AǪ��p��� ��a ��O��y2��
�b��N�e{�����y��QE�m�61J=�p����>y�O�y��C`Q�po�8d�.T�6"Od���LYVJ%p7� �^6�0 "OȤ%H�FmZ��ݙw#&�t"O&q�D�)t�y3.̔T���"O�����A���B_����g"O��'aބin4 ��Y�D�8�"OL$a ��X�r��$gu>ts��A�������� ��zy��#�O^˓��S��{b·,ԅ[�r��t�3�R�:-�i���� ��9�˚j��%K�J�6^L�!�"Ol�� ]7T�L�yU%�J6E�B"O�u���ؐa(9�#"i���"O( �Ù�K"$��ļs���y�j�U�1R*U��%�aa���y тbج$��U�\ő��?y	�'��� �I9=񸨰T�O�}xx
�'nА�,�V-���cA�*� eC�'�Pm���\K�mX�
͛$��L�J>���IL�~kh�ZG&�/^��89uJ �B�!��(&�MASm�q��mi�C)��r8O���F*R�@�ζ)�Ԡ�"Ob��]�"��b�G��
P�5"OJ����U�t�����cC4o�P	�q"O�h�mXl_��Ka�UW�0�"O��r�$΍nS�pɴ���W<ֈq4"O�(���_����j]/ۨeS"Ov�2Ǆďf��q�cȇ!r I�$"Oɲq��t>:M1G��#U�d ��|��)�ӟ���r%���vQ@Pǖ�s����(x-Z�r�e�_����&�?/��Ą�t�ۡ�Zk���K�9{e�0������rGڜqQ�]��� �ȓyR�)��@��)Y���D�˔���Nd��I�
/	J��4��{�6L����<�'�&jP2	2�"�[D���n�<��c��;h�Trrn��xhZx�A�r�<yp�Vu�x�Pa�Bh3
�i�O�v�<I��,<Ǭ�h��	D��	L_s�<q�,ԧy�(�BFh�c���Q�q�<��TX'J�k�Cކn��[��D�<�6%�`�&�Y��Q
M]�4�R��D�<Y��ˠ:�TŊbP�����g�<A �3�P��ed�+b���8T������9�0ف�e@-1�(��a.D�d�'$\(c�Y �gK�A�b�2�o.D�8�cȓ=!�ReK09�g� D��QQH����K&��5W-����O=D� �̔�>l��N��*2q��5��0|b�JX�8�{ca�?Q�6��Ah��hO`�G3��4B�r���FgED1 �B�'5���C
�R�4�񵪓�1薰��'j�k��^.��e%�0��1�'���q�
I�1,hcԂ�.U� 	�'6��ՅO>W
t��nՃ.�Uh�'�8@0��@���A���g�&�	���hO?� ÕO��߉jRLP'�Gh<�AmεG��Q�=�Na�ק�	�y��CCl��4-de�&�I�y҅V3b^��V�������bEU��yb@[�����	)�K'���hO���I�mI�,pt���(a%�\Y�!��E72�<�����n�s��ƎWHўt�'c�����K"a�(���%�A\̠���O>B���c�c���,~H !���]~ B�ɾN����o�3��j��@���C�I�/�>�8a$L�@�ĸz����(��C䉢z����!X�&l��X`.Y	4�C�I�C� ���C�@��x���C�,a�D���O�)����t�mrX��d;�	:8V���M1on��B��0e�C�I�?<.̓��|�l��OV�}B�I(T܌y��V�\Xh�D�C�ɞU��1R&B�-L���+�͘B�)� ���i��,fHI�d�z;N�J�"O�܀��<u�@���$:�l@f"O�����	O��˷�щC&9����F�Os��8q%)MI0@���(���'\�CMP�H���ʃ-(>�lܱ)O�=E�tcT&8�X۶�X�5����^��yҥP�y�&��p���+��p�#'���y"㊐`T���kK�!K�!�r��yb��F&�ݚ�bĩ}�!�r-ޯ�yb$_FPР�`#]�H��eyg����y�@*N�R�匮?Y�)7$ɔ�y�Eݔ�S� ��0����
��y��0Sl(6H#<4�i��ɉ�yrDB�J�D]�(ލmXʴ�uE�ybDF0X�~HEќL��I���y�	X. ֘Y��	}D��DM�.�ybK��p*��G#0�� D��*�y�藵U��(saCVjK
`0c��;�y�DN�İ�2�EA�_$0ezwM���y"�ݏH>4Y�%�.]�T`	�&��y.��:����A�R�Iys�@8�yb�߁Uf��i�!��6��3�Ө�y�h^.&̀�q��z�T(D���y�DͷxLZ�r^�L�,�Ƀ�Y��ybM��Y~� e޷o2|18�/˩�y"�ް]�d%8�o�[p�0c�[��yr��	}h���AkGԿkH���v�I�AnВ"}�`i0�9KCp��ȓFI �)�KNfH��a۵A��t�ȓ
���g��N�z����A�]��j���3 !V�$Ȅ��C�u.��ȓ�d1ҕD�Z��0�"��H�Ԇȓ0�@����^�$��F�Vӈ�ȓx�@A�dϟ�\L��`f E<K.��m4$t*��>Ϯ0!��F����C�t�����e�����gϦ�ȓH�ȩH��%n6j4�p�YN�Ȇ�� +�=]�*�2@�w9r�ȓ>
�x.U��B�ܢU��X*R�;D�8��	���lx�N��Y.hY[ �8D�$z�/.^��L�įF�;-,!QD9D��b��UY*"���X��E�Ё7D���h[�^��IAȄ�8=~U)�*6D����9��x�.E�(Sh݋Q�3D��ӵ��$p��X"v.�3{X�07D�,b&'T0N��Zs�	�g�H���5D��G
����v�[2\��)3D���2o�����^�.���"Uj6D��K��X�co�P2&�;J5z��!�.D�(��F�4��	���|�z1㑎8D�X�a��O �б%�	e���ۆ�+D�\9���:<S���@ ^����)D�P�) ^���'��6t�Eғ�"D��b׉
��`m���=kF���d�2D�9RDQ�A� ���W?]�d���.D� S��5r稡���%�Ri�-D�䛁g	Ju�5`��s6N���H+D��w��>2�Q�b�Q�xa�F�&D�l!󨛴V2@����R�b1��)D���&ԩi�Bl�[$C6u���#D�tض��#S��ѻqɛ�I�X�xSb-D�@�b�z�\@�_7G%Z�-D���D�\�SR�<"��
Z��@5!D�lqaF"̠aȷ� �L��7j=D�� �!��D�D��Nr���"O�qaF.�:9�u�U��#q��"O}�a$&e��h9s ,��'"O����!D�&ٚɚe�W8o��""O`����}wN��P���#�|� "Op��s�Y��2PB N�G�hh�"ON=;�@�N�� k�A�8�`���"O.aQ���2��w�b�	c"O�Rŀ�>N�N��u�Z
O�V�"O � ���,����0n2��%�"OFyqr�V�j"Ǆ�"5��J "O6\�v(Ͷlbj� �_v����"O¥c������u��`b�1�d"O�3&�#�f�R�+A.{u^��0"O�h˔eܿY���0���e��x�3"O@���G���
�7g�:E�ȴc"OR��4�֕w�h4z���lup��"OT}��'�s$4�X�AR�`f��c�"OF(pB�=9��\:�!��(l0��"O,y`b�+S��U3�+�%{\�)�"O��:�,��
?i񏍪XAn��"O6}��n�j��d�%D��^�<�b"O��GiΧ`����i��f��	�A"O�+��r��(�3s԰�"O*Q	�"ٽ%J`y0g�)�Qqg"O@�(@'�uU�@� � �h9�"O���#�ȥc/ �
3Ɋ�7�q��"O��1���M��r�ؚ����"OX� �f�\�
P�AݍP�d�8�"O�i"W��7)��a3A�~'4}��"O�{'`�U@F4� Òe:p���"O�i˳�@,v~Ա�pΎl:R��$"On�8��[����T�='�0�t"Oܴ@��K<\͎���{��t�G"O�	0�I�y��p�J	g�>l�e"O�l��h�F��ѧh�1[���B�"OD�0&�MbZ��k凃'M��!I@"O�ಠL�"I\���"7��I�"O<����	4VĖh�$�	��F�Y�"O"dy��̞0�L0�f'Q����"OJ�:ED�>l���2W��g��8aG"O�] 3�
BS����)X*UB��U"Oz(����ތP	L	\F"��v"OR�*�V$
���	{�|y؃"O>aq��J�E�	 g��h���K"O�uZd�_�Q���5��C��ݲ�"O�� �OA�X#ʰ�R�"���p"O��a7-�7!�dB�"Q�`!!"O0����&V� �ʐ��F1�"OZ P��O�T��J�T�;�"O��2���o6�s .&��p"O0��C�?�B����ό&���"OZ���l�. ����C�H�Du#�"O��B���%vd�@��6u�&Yh�"O�)�w��<������/y����"O��)l�(hD4�����.���R"O�3��/J��R �
��Т"O��Д��� q�dQ4a۠(�La�"O4p����m����3uJq��"O|mi���?R�a��ߏM�q�v"O
�@ɐ+c�̄�V㙺e-
5�u"O�]�/O5j����#U��xB"O�4�v+L�#g���G�H�%�S"O.�u&&�c�mQ�c<�y�""O� :��c�a,�-�6���"Oļ�$���CBl9�0���F� D R"Of!ZA��L�R����3~^���"O�Q�?e����IO&G�|�#q"O�����ֹ"|@`{6B ^V�� "O"Q�pN݇6d%�U�fr��`"O�L�t,�d^�U�6͏	xq5`"O��Af�	�e���5-���zq:�"OT��VA�NI���j�H��@"OV����&�(�B�kE�[��q�"O
h��)H���(��5]r<1E*Ov���;XC����"($��'J��B�R�n׺�����0��ؒ�'Լh�`�S�gg�$!�΁_BQ��'�Rջ��
P���A��@�&�\P �'?��J��Ͷ�ԙ���:�<��')��J�����2�Z�	ڼ��'�6)8�'�HD|�`*Y�����'m�hiei�ĭ�IΞSO�	#�'�X,��*U/ �6 �G�(X���'[��!��]�+!�1�G��{��d!
�'���Jr��|����r(H���' dy��Z�dA(�C͟W�J$h	�'���5��."r�Xa� �y�� ��'}x|r.�88=�%� ��-yn��'�h)�oԌT�j� �/�
n��a��'��t��ȃ�ՙ��(U^�
�')�sJ� c ��2F��8�
�'���CU0g���Yrǋ�Wnn���'�:  a��<���	��W����'堸S`��c�J�p�M�e�P���'}ޡ;W�א'	( �B]�_k�i(	�'�A�r�ǩ0�='�ٝQ5�H��'5��n�H)�@+F�D>ȤY�'
�`��.p�y�5B�;�Z�!�'?���j;��$⍧�%�T�<������Iޒb�z��6CXv�<�1�[�.WBxJ�!@�yH:|�FXp�<	f��(���C(]b~8hУ
j�<iA�W����3T�F���\��g�<ᤥ\!EFh��Μ���h�傚e�<q`,�
A�(���ė�&��|'mA_�<a��ԣ3�^�@�.�n�0��@\�<���ӪC!�9p�% �LZ$�[�<�%�G=y��|��
9厸1��!�ƣI��Q�!� dz��8�`,hX!�̔�b�s�gT2���j�ʂ�QX!�DI��MX�L�G�*�Jv�]j!�d�\������ P�⩢ՍI�s.!���BE���E(���F��6mΕ^!!�F|�h4ж�D*}�l�:�I�!�$�7�<C-Ɔ9����ǐ�=�!�D-@KZ�F� ��C�J� ��j�'8���e##s.���F퇔�x��'��j�AF���HA*� }&����'�.%)B������.6hӄX��'�Li��
�U$�!�h]_rTċ�'-�%� )���q���Q���J
�'�8�Y�C��V^m�Ԏ�1�d<�
�'bt�+�@�P�)7d�$�v�+
�'7, ���m#�mJ��S�:М�
�'��a�#�@ @��;(� Z�[
�'�i�"E��&��c��g<��	�'����c+J�[l�(�f�M��
��� ��[ԋ����˖��2��Kf"OR��S*  �n���Cͩi�Di`"OV��L�3+�4l�'�8*��퉃"O��S��_�L p5�Q��-̲�k�"O|<4��8�maUX$̀MX�"O<]WIոe�0 *�f��A��Y8�Щ�OI�	�����@]+j�4`.D��i����2>xX#*%�V(�Ch�O� ��0&B,�=�<��o� wԄ�xa�d�OF����f���)U*��dx�@"O����:'#�TZ���	 `a[T"O��0e.ˏty�-�ĉ��?�T1�"O���u]�n�L�:%
�9�܅3�S����:�S�OZ�5��#��%��	�� �j�.�P	�'����D��$�J  /��2vX���'Z���Q ћH��!㦍�{du��Rn7�>3������ -Ī��Ո��r;!���)8l!��咉�����&�5j�Q��D����35����< n��e?�y�"�!}��GL79������yrhT�=���PukK��|�y�#��y�ï�i���y��p�g�X��y�O׆IQ��4g��}���!��O�#z�$��F|���q�8򑍈z�<�E%q�%9C]qUlْ�mE1�Q�E{*���V�	�14���J�:\wԘQ#"OZ�i��.4� ����2���@����"d�,{��u���Y� �thrB���>��O �0���3 ��P�Q,����Ǵi���$�1}��xAԦ�\��Y �Y�\O!�$[.���!�Н�l�a�<!򄑴>�ya6bˣ��ڀ��)2�)�'F���8�6xj7��e�L|;	�'F�X��#Kny�����XjF�`�'��$�N1]�J�y��a��ɱ�'��p���;�:3�b�p����'ў"~dfB<w��d��M�\
\{�d�[�<��+L�f����O�'.�F\�Ȱ=9E�
�ڔ�+K�q~H!A`��8�<��4G�~�����$�M*�dڦt�"]��]s�ѷ�".���۟L�6a�ȓ\��8��@*s�0� �Ť\�lH�ȓ�l%P����b\��Ś���<l�q����0l����k���LmH�N�F�C�ɵ/���ϓk4a�)�-U��C�ɵi��q!W��PP��?]�nC�	��Np�`+Ù%㞈�+6�:C��>ag��c&�U7F+>8A ��Qz�ʓ�0?�2Ε!Y�ҝys	_�<��Tjx��3*O@X	�حBHR Q�^�����"O�Lr�/L�h���A�>�Zex��ɒ2Q��)��^<a���7W��HG8Y�Vфȓ=f�lq�A`��}� �W��F���HO(�}Bp���
�kg�[# ��yc��K�<1c�W83d	Cc�6]~�	1�N�<B�-xӚE�0o�D8 �J0@N�<q ��o��A_4L% !2���A��F{��t`@�ȐMϬn�R��FHN*�y��-g�N�� ��B�FgP��yIÜ
J��@c� #Ԙ![�H���'Mў��(��k� �8��R�k���۶��6lO��)���,En�éB*���W�Ib8�+���x�\< n1/�e�&h���S���	��H	U�S:2�09�-z�z��DC1򘧀 F�; ���Yеe(�ye&��d"Op �d���Moz=��1wI�9���'8ў`���p�$p��F��B���it*.D�ti�ϝH����3�H I��R�.1D�t�B� c0��bG�\N@���.D�x�2 L�Y�X �����WX��rO"�O�扁 �j�Ђ�:(ȑ�]�d1B�IjN�y�i
���9��@�� �"?q��ɑ�#x���ƛ3hK�a�Rkݑ �!�䒇K���:R�W�lI�5�����������]y��I� <�q�,E���*c�ޱUJ!��ҧ?U6:�� �ڄ�N�@D�'�|�t�m�C���Dъ\IC�˫�yR�P5`Bg��5^E�U��O>��Z1,��0ceFI"O���sO�ߑ���?�O�
��EF�nz�k���:w��\a1O�|	F=Q���IŘ�����<G�Ԍ�~�d���
:P8Y��F5�yB�[/N�;�O0\$����yR�ֿ6�F�d��^�QE�٠�y�
�%;��!�4A^��@��J��OV���
9�p��kѳ&JL]���Û3!�d_�e��HS�@�7��ꕎQ2&$C�ɴe�d3�J-k�.5Hd�ϞB��B�I"@մl��I���m���4O�b� ��	5?�����U�(��P��Jh�O��=�~�'�ӻ�vL
槞&xR���o؞��=ir/�u�A�a��2�L��Vj���=�f��$q���+"O|�fg�<��
�#�t��i��|	�r	�c�<��K߂M*� �r#_^:PB�-Z�~���~ښ'e�p|Ƭ��m��P�j�0L�Q�\���۰?�����|����$bך ��m�O|��w�$�	�?O��D�&/ƴ#��Ҁ�H)�:O0���K�h���Q�(K����`�L�I�!���p���Y�]�z&C+�!��ƽmʂE�!N�c!��kR ِ|֝	��d,�S��/�1z���Cō2g�֑q!a���O"�Ɛg�)yq�3L6.Xȓ����G{���'��`0C�,��xAF��O�n�m�������)��M��О^�
��4�	$C ��`Q(�O��0�^��mD�Y7ZY �%X+h���6f^(�,�8X��I`7��Af�d��#t ��`�[-�;���$�����v9�v��0�P�C#ڜ� �ȓE���Ūz��c�͛I��D��'p�a[�H�Tz@1��Ѡ=p4��,,0�
�`�\��w ��66�H{�'�T�0�U7�< ѳe08@<I
�'W�P�בd9^I�'�B.0�%�	�'	���f�T ]I��j��3/�x�9�'m,�,��4�b�K� ͻ+İ��
�'�$92�[V�~�q���)"�$ �'�rsvbkW��Z𨊦�$��'��@�w��_��ᇌǋ�>]��'[�%��^UE& ���I]H��'�B����=)ن�1�7J��l��'Ʈ�u!�B<��WJ�V��Y�
�'��`�3���)�M����'~��C�6�2����\0=ε��'��@4��i^��J�FߡJ_8q�'O�Xk��)z��sf�2>�����'��X ��:T�kФ:0ļ��	�'���H�Lٍ�∢'�>�0*��� \�Y�D�]�z��� �_{��X�"Od`:G��/ZX4Q���:|�A�*O�(:�ˋ�~x�G�	l�q�'=�3�i�G�
�2a�;ňA��'�&��#j�x?
�8��M=}���'~
���)�:��A�WE�y���)�'V�j���S}�����O�kB�
�'GHqt�ٺJ�va`���[���	�'�*=Cs�ߣt���ǈ�2\>���'�R]D镩C�>-�&�	5�͒�'LN��D 3,j�GP�,�V�"�'%�;��ɺd�F}�eM��5(��'@� RO�M�>��E-!+hzl�
�'骡�ՍųW�����͑)8VhP�'[��2���QRh\�t�&9#=c�'0��
���>#���)���g�� �'J.���c� "Q���v�/S�����'���N��<8F%Z��f��'�j�#RÛu��٦�ıcK�I��'^`̩"��*?�*�A��݆YWr0�
�'��O�P}�z��ˁSv��x�'dp5��͏#mtJ�Y�N�!P�^�B�'l��2��J��)��RS-
�	�'�ȔP��W55�n]J4��'D��p��$���֪��Jc@�z�'v��;��"R~|!��A�.i"�'̚<�"e�Ui��B��I�'����_�gy~�bÅ��^Q�',�����Ƞ��"��"�8Y�	�'ȊHj�D�v�1`��]�
���
�'8]����8TFJ% vc�<$�	�'���*�!�Ey�Q� �lU�	�'���I"Vz+��B��5��#�'��	h�ϣ'/XZu�]'�D��'�"0L��/Z�"T c���'VHAJ�F��"�4�{���.0�
!��'E�������J��X�m�+/W�H
�'�d-AA##&�\���N�"1
�'��1!�%[8I�(�(��^;E�ȉ�	�'���ip≚��*�`ܸy��'��9x"H˚��}�c�	�Y]�ur�'��M�@�%����Ȼ\�%��'��!�"X�7<&A��ӜW�-1�'������~K ���VE�.e��'���s�Y¤<�!�D8S����':h�t!��">b�Ҁ �3=%>���'��K5ŝaN(1�,a��i0�'�ּ���V�n�n5
m�,
0N<
�'������Z�4X:F�ґHO���'��(��nX�DNb�yA��L����'�\�0sA��P���e !Bo�pX�'��|�g���]0d���A��o�ʁ8�'��pQ�K���>�d�*Ƨ�)�y�`\������0�J���!N��y��z �Q��A�"��\Q�A��y��>	���	ǌ�+J�"�Q���y���)�VQ�Á�>Y�LUR3�y�dۋSa
`�W1�x�����yR*7qJ (�0�4v��$�%�y�oR0b<%z��3�J�Z& ��y�/؁(E`��&-�(4G���J��yB�Z�t��á��4���2N��y��B�8��q�@�8�60[r�7�y"�J8�ؐȳ.D-0�|�{�߃�y
� ��{7a�h)v�?8}��r"OL�i��_$T����eY�zo�p"�"O�ej↛�_<|e�����Wo����"O��玱j������0zk>|�C"O�j1*	<u���fJRG}�1"Od`�EE�^�t�5�'6����"O��2w��]�T�ڦ�� T����&"O�ī`�3-�I ��o�H���"O�\���J
^�X�樜#Q�t�a"O��C K�vӨH*%��G"Ox3��.����� �a�����"O�,�� � J����³!�8��"O �`��)w��yaCq�z`�"O�1tK�<|�ex�"��z!�$L ���roJ���*AJ�S!�O�;�qPd�	�%3���Ys�!�D�����O&�e��`éI!��*~`�� "��G��`�'��Q�!��	�J��A(�3���WcL�^�!�d�) )��Ӱ��p�0��� �)+!�U]2�}�FdQ>��x����H!�$�ir���,�;`0�pk�'_�N�!�/w��l���+E"�83Q�×C�!�ǻEd�9� ��������$!�d+0��o�.D �Id�9>'!��	�eB�!A�U�q�64�'ʵw6!�d�:mpb��_�<�>�+u@�P'!��T!z����M�8������)m)!�Wq&*�`c-	o�	
� P#3�!�G-?����폅E>��Ů�	
�!�Nw���b�_'�J��S��Q�����v�?��(��B�f���c�MZ�&D���'J"~"jQ�6��*?�yQ.|V�0�g�Vu�)��<QA��s�^Գ�'�9u�&����](<)!�B7[����a�"`�mQ�O�-E��\`�Zy80:6aY��=	 ��.6'4��4�6R5��C�(�G��)�I�&C����ф� @�0�޴x7 ���̆z!��Z�D�4��)�ȓ�~�ac�R�b�#�-��v��8�'EN9�%o�k�!r" ��Zl�F��&I`ܙ��oVt�	SĊ�<���pA�]؟P�!Q,�Z�B�n	?�N���Z}
	�"ME)e������#]���l/H5SǄ���c�R
#k��$dN�IV*�/���S*��*���/)�����7G�`�B
�1|���򂀎O�"\sA�'(��K�@��B�_��8o2��d�;Z�fQZCB��D��?٤�ȑO�p���)��Jp�{�iZ'-�Iw��@��Ԛy��Fh��v�F�'� 8���Qb�g�I-)��bJ1m���ڤ�]�X˓(��Y����{ul���JD�~�?A1���	@�u�u/�(\a�-�5�V�n�����[�a~��ƤW�4��%��4i��RSF��@�vp��ÚZC���MV`���a؟0����X�3g���O(j`�F)��d��h]L<���',	Z?��ӆ�7t�<�cѱER$�#��:kt^dC�Π84s��>���"�SMń<�BҚF�88[�!9�J������ ¦�X�C2ёu:O���p��-O����Z�E,,��r	��
U�9�Tx8#�3�3��BN�D�� I�5����ǥ5V�ɶj2Zac5F�Hl�@��	64T(��D�H8 ��	aWL�}�,�ʁ@�5��;��w�a~H��cx������%<����ӱ���g��X�( >s�2k�0a}��Ҡm�$>���ӼKQ�ťE��]����Lk7��N���s�CE����gMN�l3XH�l�T}�p*�����@�v#Ձg��9Y�GLg?�v���  �Ӵ@��}��j�"�J����,6J@D}b��;�*4�K�I��	�rS?]��l���}#W�G�TZ�Pe�<��M\��vpY�",O�)P���8v�BT�d��J�ƴ*`1O�{W��J>8 ���* �!X��TΌ�� ���8L�5 "/�3rbt�����Z|�ē����ǀ�v?T���,S��^r�x�Åc*Ԛ��@-��ѩчA	u>��yG�ʔ$�z݂DJ� �r��nP���>����hR�A����Vk^�lo������q�X��뜽d������?}2�8~�`�ۃ��4a�� ՚������~�J�`� ;sў�Ab�ȴ"�6��&&^�0� 脮��|� �!�惒�e?F�������J�\��8�/�;��F�'�l:�D�:{����V-�#t'�ɀ�N���G�Xmؾ"�b��[�d2I~JW��[�b �4o�0��)^4��-[V�ӪZ�B�I68�*8�rG�

���גjH�O.t4������d�A 69� ,�2'J�i��;$�A���p$�������*�O���U��Fi�L�/��6TM� �J�
�AÔ��W�j$0��	�O�pyd%��')B;싻Bێ	1��@�d,��ú�;��8}2EE	a!�Y!���2'� 8��l�$bS�Δ�4x� ʿ*&R�G���7�!� �
H9sp#[��0٣j�&	���T33d���K�8��M�@.����A�if��D/���G��.���Ѐ�uSR�\����ܵJ�Dl�-��*@(Oʸfn ��N�G��\˖O�0���k�f��N檁2$IM7���	�v�0��Ā'�B��3��ׂ�<q1��s�$����/?���Z�~�AR�L�A�Y�bLZ�zqz(�q�dl([(����K�d܊��p�@�)��I�.]�#C��c����Xb��>�[�V����E�9mީ����-sH*2f��8�̍|�p�1$$D���	��۸��S͗�N��죟���T�n�|�7,�aJ��Io�D��&�&{��S�*6h�S�	�3*.dm؆�ٽJ����$[d�2AJsJ��|(�u�	�X�:y��	�
ـ����X��䓶H����H���3�	�Bی V�DQB1�$�@�Z@Ң<�E��Gј9G=�'��)�傳:�t=
��Z���D$$^$4��m7�ON�qC��.+ ��'��8�!"�T6�����@�}�1kF�ᄂ� �槿ta�J��h[B�
����F�<�r.G~�Y�e�9��([�}?�#GM�+�f�i�9}��N�w[����H+��j4-�����=�
��d����>�4$�r�46MZ�C�(�0�S�EL<��5�
0J���X�3+�c6���Ջ�ޜa��T+O ���GKfG�~BÙ�U(,T�F^�q�R�R�����b��6d�Q
�iU.d�a}2n�n_\`�gU�q��i���O\x۲��=1���{��*bBZ��&H���ʑ��!��u���W�]H�C䉕y��*B�%�E	��|���x�X�P��-HE�4��t�?=�c�9xG�!85�K,V�8��"%D��c���bs^H��(H8�VP��?3@�v��4N��l�3�Ŕc�����'Bց���T�h
� 1ynP����4)	��Ξ2w(�##��]�f�;���*���y�gB<4.0A�(6�ONI��2D��E�,�5~�d�+����u���p�b�R}�t�٤m��p�q>�0$Ș���E�Tx�� �#D���E�մd���3�`�	\�be1D�	YaRYcFlX:%��U�֔N8���5���yWo'����+A=m.)��j�9�yR!��%�tm�<���E���S���2Iиi�cڌ*\L�bQ�9 �9�����Nf�$+���*"q��A&jݧ�z�
�"o��
W)nq,���X�ƽhլD"mm|����I�А�����U�N ��I�]}���)K��8��E8R�P�La�b�Z��ܺ���w@E�6G-ʙ��Oin��EV��Fi�#h��,[�'%����UsP�p#�nϓadJ����^�Dm	W�L�0��,	f���H'��?��39�$[b
ϥ"�
��l�P�n੷"OT���ME1�1�
�&J��Z�GE?s��$1�#�t�
e����tyax�H�mE��@��5I�&�cW�ݩ�p=�0���̽*�j	#�M� $��n^�S�ʤTn DK3,@@�<i��Ă'f��{�`9���Xܓo��A�p���V 49�􉊖:�,`iT�؇xoR(ڱ+ŖHP!�$\�䮽��A�^��ͲqL�J�ʁqN�:[|�'��#}�'BH�'O�f
&���]"Re�
�'���`èȧR٤P)⊉�W��Y��6��t:���0>y5aC�'^�[�JX�}.l� �`
@�<1�F>\�>�yB�I	2�Z��gK
x�<�K}i:�k@"�p>�� �x�<q�3�f�G˛<-9F`bMy�<a4��!v��.ټ�y����z�<фb��]�.|҉?�&�h��Y�<�B�Dk�AB
�fd0��%DQ�<9�h��-[3�Rq
Dc��L�<�e�ا
� ��b[�H(Cm�O�<���$6��Sf>$�0�J	G�<!�+\$ܰ�Y�&�'(�^�CgM}�<� �	 �C�$<��<r���R���!�"O�pA䠛�g�}���ڜD��بv"O�dbI��8�V�@7���v���y�"O �X7 ]�~��F�B�M��t�"O����6zr:�J%'�l��`�"O����B3_P8iCF�.tH�"O��e6Uҩ�Dd_�o$n��W"O�):�.B�o�-@�B0�4{�"OD�'dT�+@�I�&���"O�p@4$ӗ"�z��e�^5g�>�"O����fH V�q��@�^�6\�"O�i�!�ԓ=>)��'�I��8"O2�����bp�l3�i�3�J�"O�TC��A/z� ����
���"O���WbV6�&Ȓ@��O��!s�"O����-�'_��97 ++�i �"OFU i	
�^ɸ�j�rg�|0"O`ͫծ��K��銓��T�#"O�hp��G�^��J�.J����"O
	����xԄ|;%�E{i��{�"Oz��԰F��h���4^|�s�"Oڱ	�,I�t�c��=D�x��"O���-?�J��O�0~d��rw"O��;t�U�Oɰ��H.Ch�"O��ҥÏ1eH��"--J$��K"O�̫���h4иv�H�N)<e�"O�PDʕd@5LƢ0+25pr"OTp#�B��b24�b�NR'��G"O&I�f��
;����
;+Aj�"O� [cB��{���%��P!<��"O
��MǸ'�^�*�`��s�"O��A$hL%�<h��>%2��9"OFMxv�O+��u�c]&�Hy�"O&ɺ�m�4zǨ�sp��u�:i��"O�Ո�K�%�t`ۆa�4R@��:r"O��ȳF��֮�) AVAh"O�DP���	!��I����K�V�("O�:�f�)I���� �
5 $P"O,�����ū�צ3
D�hB"O,��T���;W� �瓤}�0L�R"O��b�EI)�p����j�>���"O�HA���D�� ĨU#X µ"O�1A��B �*�Ͻ7-��4"O|�0U���8�M+Q�K6>��9B�"O�4*�A ,%���A�1�h���"OJ�B�cN!?�I8�L�{�<kw"O���nȪ4#�q�G%Ѻzer0�F"Oh���B+6�ƌ�҄��,k~t"O�mq�&5O�T(2�B�'vID@"�"OX��a��?Hkʐ�wH>&Ya"O*5��l�I�TA��9^�D"O&��s�ǾKV�ҧ��'6�\��T"O2Q��^&h-� �*(׼u�"O̜�qDR)c��X��Vm��qD"O"��U%�8aDblzGj��0�rP��"O������'_/\(�1�����q"O hä��w���GaՓ{�|	:"OR��WIE(E��a��E�&ƈ��"O��b�`%\ڌ�1�X�-貅�A"O4�D��\)��q!�7μ��F*O�+$�KR_$�P c+]:�T�	�'��Pj�Az�L��Q:����'�⍢�'�e�J�&oT�x�h��'����bM�:b� ��[�z������� <ܨ��R�7�y`堞0�h�5"O�It�=qJ@ԎڇF��,h`"O�� ���z���- ���A"O��!�ـ�,h��O�8t�'"O��+)w�T���Z�^4<�@�"Oj���C�z�=��I�(.�r"O\  Ҍ�7��`����/��"O�-�s���~�{"�@�r�4�P�"O~�z����N�2�W�q�$�;�"O��lq汈�/���� �3"O���H�lڤ3���f��!*A"OL)�t �(h�)�A�X�Н��"O���#�ˆ/�Z� ��5$9y2"O�i���i�%��C����y��"O�!r%�k2�u��cL�{@��"O.)�@���p)+gE,D��"O�hsr��o�xkq�_2@ rQ"Opx�J�H�VyJ�-��bpPl#�"O�e�7	�0�!E��]HH#�"O0��c@��8�J�#v^�3"O�]���8	�Y���M�jK���a"O��"��$�:snۇ)R޸j�"Ov��n��|��g�F�H*24��"O2�Y�c�%V��1HR�(1�4� v"ON�*�b^8#\h�Θ�I��t"O,�ѲKC]�Yz �L6<�lc "O(i�f��	t�����.�']6���D"O���@��>(�#lX�+p�	3"O����QWȜs�+йQڸ�"OL�ڒ(ڪ;�c�L�#_����&"OKV�DF�E�g!�+LQ�S�I+�y�ˇevID�Fl$��^��y���'� ���n�
?I�����F6�y����~Wtc���5�ޙҁ�C�y2�دw�T�Ab���*��a��^�(O���X/���*@�c� 8S�U1�ĝ�B�ܬC�"OP8��㘜 ��9ҒޤZ����,i9��)�J=��s�x0e��qф��2"
i L� :�8���CC~\���^�Cnr)���Џb�\9*$���l����f�B؞���1l ,�VOK�h�R 
D7O��@S���xX�]�4B�"���oZ�2���;D/W�8�.A�#�/XhC�	*p�r$�Q��<����@+R�FKT��d#�H�`QD�]�9��|��"�v�|`���9+(� ���?(fd�A�*�O`�1G�9"����D��[۸e[3��8OnT�S��K� ��ڴ1e��I��p"G�o�Ā4N� ���=�E�M�z]��e@5K�œH�s� �ؒ�N�~�h��Q?l��`ag��)+���GL�:�Q\��O|BEy��H8wE�&W�@#	�J�'�i����t��B&x-��;�:1K� $4�s��,��ݓ0(�s��ZV=��L>�f͙Y���B�N4Vv�����vy��ʰ>�@�i��-TװEC6�x�'j�"��Gꙿ�$�t��lDcdA�e��Fφ4�0?�$�%��q���8y����=M,�q �
��MgϒFH� ��O'��!sEC;~��8�'{0	1��ٶ]I� p��&I�E���ky:	V�#t���P dR%2e� ��%֬X�p z���J,U
��_WlٚM�P�d�ܑ
�@ ҒF�fV�]HwA
�D�axB�6�. �B�øZ�4�'Z�Ay�%��'�8T��̿|�X�%����	�}'�l����|%;J��DxG�Z3
�H��	����I�g,H�KӯZ��0sW�)�yS���4'��PĒ�	�
*�Ӣ�u��ѫŬ�0?�d)�7w�����9N��ȥ���J�xiS��9�� =H�zi[�Y�/������9%�q�!˧)�v����9D�܈6
�T�1L����VF���=�R�1*�U���t"V�- �>�K���r	
�P���'�҈abX�<	��V�'NHQs3M�1�H5�)cybMM56Ҍc���dX�x��k�>F�%�������"�O���B��4{�����WQ�l;�H�9a�<�&\���x
� h�3���l>ɚ��M�WC�Zr�I��X��g��M����@Z���%��$1��C�ɉw"O`|u�	Wr`h�ѷ3�vP��'�� �' �S&u�O?]��o�B
q�cK��IT����y�<����*B!�!E�̼��ȕwy���8<tDp�"�cX��YE�E�;-�h�� ;�: c�-$�O8K���V2P��F�aB�G�,eA�"f�ސxR̖oBpE�ӡI�M�;4�\��Oh����H�
p8�?Y���gc����$��Pm���*D���ǡ �[Z�y�I�Z=Hf+��@���M36MqO�>=�qi�x��a�FѲD�9���OIx����������x��[�Pe���6(H�,�pa)D��%e�4G�2T�F�e���4��>��!�7g�%��ep���G��TQ�m9��D��Ą��.X^�b�Y�l1��tK�=���C
R�^JN��F"Or�/�b��j�) ) f+��ɱ �b,R/��`�O�v��ŏQ�d0Õ��;Qs8bF��Z���z�l�򃞄D���g#�2L6���'�.3�ytkY@�DO�,StĻ�H�s����ICN�g�N�@���3&�Pe�"O�1I*@�����H��]�'�Opz�H�5:<�XL�� ��Q�hstܡ��\0�ͩsVD,�����P����n&�OFuk�Z��P�l�%u�Z�9��s�	Y�G��I�%��%B�Ԏ�axbL�>ӊhI%��-C�JL��.�(O$���E͊;ۆxYM<�u��qL}a�P�
5K��.tF�����T�!�$Ǯmڵ����
?&5`d�۝}Or�ʖ`��:������>��m��p}���'}��8���S��|޼\PG��,d pM�ȓUOvD�T�U�)W�9@���3f!��{��u��<��'�\ͻ"��&.�O��LHq�R?㈜j��;@��	�D�ˁ*n����ƣ����`��T�U�>	���%Sˬ��v�6O(��S4P���QR.��D�Kg�'�֍� ���݀���DŶf�ڱ�F�ٳJ5|(��MțiKPd{��'��y�#S�iP�a��!S5�:��$N#���h�*��O;���/�?A3%/��j��;6�C��<��;D�@���E�<���_�y[�؉a��>�ǡ�M�������h�,lHb���H<B��ݿA��*/K���$�W����(	xǤ�Qd^��)���M���'�JB��q�~�?���O�E�����@��P`x�a��4��;Ӗ�:l�=Y^�	0�Kԭ|\A3�nK�ϗ�o����ɢo�D� %��~��s��	~��⟸)�P�D�ȕ����t��ۘ�ͧ(�̈ ��P=��a�������ȓ9�;�J1ݴt��oA#�J@��`�<d��@�J��a���<	��~"!1�&�ÒB�R�b���aѻUY�i��"O.L�dBCh-q� ްu��e��&M�<p)�a�=;��_5t�.H�4΂�@�(S��
ox3��_<3Y�����0\O`ۗ�͔4tf
$T/�4�@��աoa��kT�Ӛ#�zԓ�
G+P�vf<�0>�G��1LPt4��Q�7��h@��\ܓQpH@�Ə>��y��CI����!�Dse�)�4�ĸ�%��"T=d��&���`!��<ʖ59 �B��yH�� >8@�c�X�U" Q�A݆�z 갃BG�'Ar�݇�T�	B2U����ڪJ��C�	?)�����#n��:��4t��r��5��6N˭R:Z�Pc�9OP9������v,	e$4*�ʒ�'IJ�!������bŸi�P��^�)���!J5&.�U��'��!��=9:|-+V%��  n!��{���a'�N�͑>e��M��T�����}�X�0P&D�L(�jJ�K�4�K�GS��:"��p��0��Sz���M������[,d>2�jP�Ln�!�U�5;�l�s��>n�����CH�;����'���sUB�<� �68՞��'�2�ę+h�����>�f���'�b��C/\^|��, *1�jk�'k�8XÍ_<)Lȅ�Rg�*+���
�'ð��!�S�b����bn !m����'���c���:%�n�A5Ou��'1Ԩ���@�Ȍ@%I�|t΁���� �e��.�[h�R�#҄V�usE"O"H�n��7��K��2{Č��"O4��;;�ZUb��N) ]�D"Oܤ�r�O�t�p�Z��P#""O��1�LV�J�������q��)��"O4��`
{$���6r�I��"O�4چ��gu�غ�У7`tE�Q"O�%�� �
f�8l^�{^I1C"O����^SҤ`r!kW'w�y�"O����n�;R��3F������"O�<+6�hT�0)ǰ<����"Or�k�J�8 �����ٝ0  	�"O�,@c`أ":� ����q�H��"O^�C�闇cȑXW��1m(@�"O>�ٳ� 06y�q���K6\!�"O�Ejզ��|�h�#��	 3����"O�1���<S���j����qz)C�"O,@�pC��S�"Y���JJ�AH�"O�� �((���93��%S����"O�0�s� r*>}�7��S3q�t"O�x`N�<W���eDtE����"O���0>nA[�N�ob� D"O����D8#ߐ�a��Г^X^"O��rP�'��ڂnԜ8S`�R"O� c$��j�5�0� �9D���"OB��� �$1�u�î�f/��#�"O �Q�íw�b��5`͋�"O��i�f�P��$�FئRА�"O(���j��+/�PV�,6��"O�t���Ĕ,vT(�n�9?JM8"O��oM8��R��-g��#!"O�QK�	�Aa`��AZ��a"O.��$�4I1:I%�n I�"O��J�-�(i�|Q�&��0�0��u"O
,���&�� B�E�3k�A�"O2p���T�0X�K6�ڮg�^r��'�uꀱi�f(ʓ�˚Q4 ��-�>Z��K�{R[/��O1�<Qrr,��FAS�K��1��	�L����@�Q�S�'M��h`斥&a�����ZH�r�مMe��̒��Lv�6I�A�S/4��� ���(�RIɟNS%�Aʖ�`��-�%%�����t�Q�d�+���s?%>��}:�@�<܄���I/M��C�l�aLؓ�@M���ٳc a�t��,1a𜩂��bE"���2�2SV��rP�R��xb>��W�{j�Q&��X=�f��y�'�g6@@@��2e��������v����Ӂ؛O�U�w�\��X�H7	��>��٤NQ�z���9a5�'A2x�&fր<�t��2D��}��� Q���hfn��?�M��R3���<��^��FMпt ��B1�Ɔs:%rVf�k��{2>�������)�/��O�T r�'	0*���#:B\d��'}���B�,m�p!�cD�>E�����_1ȡ��W�iI��B"E�-T��U;�re�քYp?��ӊ1<�$�� ~�ȡA�f�/޾�8��AJ���7;O��آm+�h�9����wӠ��݋MVfQ�r�a�0�[�4@�j�[�I�-(_���i����!j�@��JпA� q#���y�	5n��;�
5f��Q����(�l�V@+V�(@�.�����Nơj,�B-O?7��
.mĐ�Pg�%*|`�
L�J �����q�L�J>�Ϙ�j�O���faD-�$S���C�<��鉄Bc����!F��ږ�@�<���\3 @  ��   �	  �  �  �  �'  �0  �;  �F  R  I]  �h  �s    J�  w�  �  e�  �  ��  ��  ��  ��  e�  ��  ��  /�  p�  ��   E � � _ �$ e+ �1 [8 �> =E �K �Q X N^ �d �j Zq px �~ ǅ P� �� �� ĩ �� h� �� �� �� ��  x�y�C˸��%�RhO5d��p��'l(�ɱBy��@0�'�F���A��|�^{���OM4�@hC�N�\��C����V����Oʁ-^�A�fJ/j�I�&�Id��	h�<|�S,Հ���?/�����	k`|��4��V���	�I��6xE
SA���O�,�d��_w!8����O��6-��0��(��N�t}��e����I�Ji�@���`wԸ#�	D`d�p�ܴv�J	���?���?q�7_<���d�A��9��KB;N������?i���?�)O���?����?��h�\��H�GlK�~��Ժ/�:�?���hO0� ��ia�$�O�]���O�:c���^�C;@���M,�O��ɇGR�\�U�
[1�k�a�'q
���*&��\K⬀�ȅ�P��~:�*��P���gߣ�~�'À � ��+"y�혠*L9�?���?���?����?)����Oj8H��g�
b|L9�(ȢuPL��}��i��d�>���i����p�:ʧV�Bm�$���W+�`�ǇOz�LX��D�h�O��X��B� �.ѻfd�"v_6Dh	ϓ�O�4�NF
J>����=b��Š"�'�ў"~���'{s�Q�H!(VrIzG����d$�O��s	�yda��䊄D��u���Iay2��'F�E�D�)k4Rh⠭�G(��)�|����S�KHH�HVA�2P�5��8�I�W ��S |��h#o('V��Q�� R_��$=���O�?�'$��7�C$	 G��{i^���'�p(9V"E�wF��Z&��>k�x;�'��(6J	Fq�u*��
6V,8�	�'V�ء���<U�aIQ�K
�*	�m��@�N�$T`��ӛJ�������hO"�����{�(�f%D�R�t�YT�\�}�@����d��	k����l��H��t;%�}#�B�I<:�c^�7�T�B�����B�I9+�<d�db��2p�) ���	ذB�I�Y{(E�Q��
s�i��*֘Ҫ�?Y��S�hz>	�'��g�d��%��*<��L ����H��m~2
̧	�
aY�H�Đл���yj�m�6��`̅�d\�i�i�y��ױ)��Л��  U����y�B-{-��FI
[Xa�jΝ�yBG̾^d��uL%�8�����B��(��|P��;w}��@%��1�`A�Z�b4�������o�)��610�/+D��5!�&o�NC��3E�Ƞiԇ�U�̵�%K�9K|6C�ɖjFb|�!i	��� W��v�fC�IQ\~Q�!���ICt	��X�BC䉯6pF�Җ��5�$���L�p��O�p�>t'*6ݛV�'�g� ��;$�ip�$jE�Z�x�rQ���IҟX�����h� ����������#+������d��,A�k�PP�㚱rOF�b��
I���(�4n{��ڊ}���c��x�V̅�	�D���$�O��oZܟ��Q 6M�NT���RSc�q�|˓�?)+O���I��.OL�Ҳ�[�3t��3��N��!�n�ƠA��J ±���M�=d�l�&�Tڦ9�'n����'�Ҟ��'��O27p�� A"lf>P[���w�r�'"����`N�츧�RXz6U#<]��q�.A��䙟���A�nvqO>�h��ϴ��|�4���lQ��=?�TişT�I|�Q�'8	"t)�Fޙ*v,����s*�&�l�	��hh�/̬�{ ��)Ce����6��%��>Y�0!/�R$�U��|<B4�O�]
�c%�	�?��I��'�|����	 ?�E �燁�P�'��Ӡ���1i�L���t��'�9�'FV?Y�v1*ՇS)T����'�"����W�p:D�P�F����'A��y"��-@GV�+Q%�7(�$:+O��Fz��i��ʲ�e�6�<p�Ï�%Iʱ��<A���?Y���S�)�bL�+�� ,校�b$L	W�M��O���f�VD$DiGD�
d�Z�C��d1!�DH�V�K��#ML�x�쌺��T���'4��'�2X��g��|� ��U�|Fzq��A>��Q�'b4�XS�̪Mx�e��ɓ0p�O>aV�i�_��#��O.�A�i� e�d[�=��*S�  �r�	��,�')=��Ex
� � iVg��'ly㇮r�=���'ʍ���$�����M/0.D��.�=�ax� ��?��y�P�V(i��B!��8��HŰ�y�+�9I��K��i{8��6瞋��?�p�'��i��ɠL&�Jw�Ήa����N>�D!�a���'N�t�'lL��"	)�T�ZM΂�>x��'��-�1R������[� �	D1.��,[7�Ù(���%Oʜ�C��#dA&��7Ϙ�"��n�\����eY��#�⍉L�P�*L�F��O*�x�vl
4x��ԋA�UĀ��O�0�'E26��O���-�	�O�}�׃
2l��`��T��bU�5�O8�d�OT�5LO�DY3��%l(\�rf�̍������	�h�B��$#&B�v�C�-�H`Q�*�>���?���V8���'`r�' �Ɍ�}K�n�*/ì�*!�c���bCo]+g�>,��Jǲ3�-0��W`�g̓O{��A4��?،8@�H�/"���6�րwF,�qK�u�*U#3gCC�g��Z51Ca�-�x���${ˊ=�ٴRe�	'I���������)�I�jO65q�!+r
9� �2�D��5�Lj��(���щ�*k3<ɕ'�\#=�T�З'.9�ˆ�T�z���/]T^D�i�h�n6M�0��D�O ��?����l�/l2 �2E�
��%��1n�,�PT;:Fe��G���0=9�!Ї�
����/�b��"�z&�)�h\?@�iÓ�m���P4��.�8���?ge4������Φ��ߴ��'���?!:����->�!�1j�c�h�'D��#ґCT��9�D҆R4��,2���}}��|�� �Uӟ�H��� �jp��:���5�'	�'�2��>7�J�1�����t�P�j��\�<i�FT4�Z���юW� ��bG�N�<�ű�>	�A4�>�Y��BL�<���]� l�Ps��
򰸹T)�P���:��`�T��W�;�R�"�К�F{���ꈟ����&A�B��*R#S;n5bG �OB�$&�O��ᴁ��u������|��Z�"O�]҂�����Å���U�"Ov=�E���r���t�F�,V�tr5"O�A��dʿɔUi��q<
5���,�h�B=� -$�QZ����p2����'-�����4�
��OD�^L�'aKZ����@eч%�i�ȓ~J�ȵ/�5G�x���J�&n-��8{��XG% �"�[�ņ�2�]�ȓr<�I�H�5�$S1l�Uw�̇ȓa�a�So�FX�E��`�m�'��"=E�$��I]������U��a���D<D�V�$�O��Oq�Xl� Мr6Lᒕ
h�9��"O`��V`�e<���3U+M�Fy""O������@����<�t!�"O����hӫ
źU95�ͱ�>!��"O4�s�Y�ӊ��D���;��|" (�>2�짅N!��C�^9`�CkҠ�?�J>������	.i��|����tF��
��Էi�RB�I�tn�A,ԯ6�Q�G@Q�|!�C�"}��|p���*r�  "nS�o��C�� kP�#rS	��N1�H��d�����L��X��3OO�}S<���"1�;]^�D�4(��xxP��s��Qp���/�[Z��'�a~R�	2vPt�+pD
3(��t����.�yJ[�dvP,)N$$9����S��yBb3����&[�y����15�!���Y��;%dM�fHTH��B4?џ����	Z�1�z��"�M�4Ep�x�cT���  �Fx�O�R�'-�ɉ	�V�s��ĨR@��#�ڊB��B�I4CR=�'��O�&a8��? #2C�IS��3.�d`؈{���.4C�I)$rڥb��Q�h*�hSe�υ8�.C�� �*������@z�ԡ��`���m呞�|���[��V��raZ܈(��JHy�	:rE"�'1ɧ�O��P
�J�B ^��2m�%�81���� ����L:O
����U� 3"O��9�f@�Müи�� �x�0�2�"O.��&�M�o�F��Ł�@�\X�"Oz��!Q=d.�����p��H�T�|b#�	�ڌ��Vض�@v� v��[��ό%�vu�	H�̟���O@)!�r�hya�B�"OL��f�.5��Pr�K�)�"O���#V/M��:B�Q!�bIIC*O�%��BZ^�A6j�1t����/N���;/*��Y��c��ի�����hO ��ӗF�,|�c��.s�dit�$���������	�B�� nͤ�4x�ql�B��B��2(�6�U1��sǠK+v��%��o}�8��}4$9�)k�Х�ȓq���e%Lzy��r
�$Lt�G��(ڧL�<�֊*EAV��l�����	R�#<ͧ�?Q���$�9��Ȑ�ѥm��D5i�!���	|t�3�l�T���BLA�~�!�H� �!�Ѯ�F�:�CS��+�!�D$@�6��2Gߎp�b��G�7�!�$�(*�"���n��.Řl�S)�{��I�HOQ>U)  U���D��
Դ%��,ps�<��͕�?q���S�'uT�m+�@Z�H!n,"uj[x�ņ�,Wȵ�TJT��u+�j�@�D�ȓ5���c�J~�8�aDS?g��	��e�䙺�KA�.-IqGܾU�:P�ȓ7��$kG��� ;� �b\��&�����d��Q;�č�� ��B�,R���R��6A�R�|B�'���ov�p6C��8��RIM���e�ȓ\g�����,>�p!���3���������̅�(��KĒ@� ��ȓm�%�fYw�ųv$]W�Ȅ�I3�?�#��
�6�G�Q->70MH���F�'�����i�8	�������頽��K� 9�B���O����9/��%�Fc���#` [*r�!򄔼cQ�P!6-�q�l	r��.L�!�$��x�B���R�b�b��^0>b!�
DJ�dS��X�'�~|�5 P�hNџ�B��)�	P$��I]�~�^ W�j��ͥ�O��O���<?�0��?1�D��DI��a��Z�<����c�B��.�f�Z�5́`�<�!A�$�[b�N�\��)#�b�<y#�C�2��#��H3a�H1��`�F�<9P�V� h0���C��<���FLyb�-�S�O9��J���h��L�1r��(O��X2l�O�� ����)c?|�(��8^�1ش��:u!� sXy��ԮP��,X�-��, !�D��|#`a# E,\� ���X�!��?-����ʃZm�,h2F�3�!�.fn��JwH�7|�Ic�܎m��'d�"?�I?���h�|	lP(DHQb�I
�?H>Y������%E!�ޘ���Q!�L B"OD4��@�3���6�Ë��zB"Oj4S���$�$Y�Ո�"��e"Ox��.ԮB#�����1x����'����L%C��q׏W!
FTx�q��hLў�Ҥ�6�'!�8���Q�r1��!M�^{������?��Ha���b�߿����ԁ�3�D��ȓ��ضbşx`x�Q���?X�D�ȓi��HaoҜm��H�b��F���z�
$P��I�d
0�1��X&+��#?�W��d|s��S�s��LB�-Сw�����F���P�Id~��;HLޤ8�J��������yb�)c��1��:=�0G���y
� (<R�]�Ro
�	�T$B=Sq"O��Iq`��cØ �ڟW�]�"O䯦�u"ř]|8�L�Ay"�7�S�OD&����U2�њ+���R.O���N�On�D;���O<`����DA� n�h%:DJ�P�!�dIJ��r��v�d�Ir�G�O�!�D��[�Ф��0��L2��L�c�!�D�J8�u�I�; �8����Jw!�䘼9�Dq� ��t���Q��4s�'i"?��%�e?��E*' Z��ɑ>ߪв%gA���&���IX�g���; E��zA�'+T �!o!�̂"�����T;��B��m�!�D�z��aZc@͹ D�������!�dəc�x0KقQ֊��@��#�����O�-�da��6=���Y�����ɉ4�"~�@��e(	�РXJvp�4�D��?Q��0?���XҺ1�F�3w��d��E�Z�<1&�V����V�ݗ&O� 1DIOX�<AT��"�4�cm����4ĖW�<�!��K���ە
M��t(��O�'�Т}Ce�77X�8z��% $�����ɟ��tj2��|z��?�On����T�+�N
|آD�"O&�@G���Kr�\2���3��퓵"O*X�U�8|�E�V�:45h"OJ!h�k��P�0�@9�p�
�'pe�dO�M@ɃA	T�ꈰ)O��Gz��IB�n�F��p	�5���$gV�A&�	�k(����ğ�$��>��3b��TjJy&�����!D�ȒSEզl�x�h���!��[%�,D�`�u-��d:����M�>X2:Is�*D�@�u��:�t�����,2��C�j(D�B4Ǔ� c^IF��~ٌAYr�$�$h�'9^�B�'�r���=pv�@C�![�nyC����?A��L��P K�(e��
���Ffm�&�!D���e�	�<vt��c�߭PP>�g�?D� ��,]6�ptA\�<s�8�k!D�ȁ��Z�W�,`j�Ć�c�9a7�2�O�4��1�y+�gI�jvx�q���(u�=����s�O�T� �ͶUd���+4	�@�چ�'�B�'Wn��i�:d��4K�E� �h*
�'�lu�2Kv-��A�!lv8
�'f`Q�ץڒ ���"�7ּ�	�'���Ԇ���"�B��fPX��čd�O�d�5a�s�1�	�+LĞH��.�MDx�O�b�'��ɇ/*b)UdX<Iۘ��#'[�e�B�I�g���0�+7:��5hY5:�(C�ɓ}�	xp�ӔZ;>�{�DԹ@�B�	>9`� Ӷ���0!��35X�B䉣q������_�0y�7k��m
�ʓ8둞�|B� X�=. ��q�R�[t�A�C�PyR��5,�'Rɧ�Ok��qdIgde����$pz��	�'\��ǃ�~�JEo�sD�)
�'���33��PF�h�����2	�'�ȼ�U(^P ���jH��i��'{ڠ��ʛ_��<�R������H>A��	:"��	=ن�猑J�f��5@\��:�d*�d�O��?�'�h�R�j�YQj��P�ٿo] ���'�����A[������g0���'�Ѐ���Z`GcɾX�4���'Jp��S��,a<�Va_�R:��A������l� UH��d4�CD�*�hO�I��6\�J����ݓ~�nq��7�D\���|��I:u��̘�E�W���hqfܐܺC�I�9<i�b`�  +�պ�酲~�HC�)� �<Yf��7~m�&X;9�X�"O�U�A����p ��
��"�Jx����2�h��u�'�	Vhj����9�c�'�,`���4�����O��\��Y���H>?G��-O4^]�\�ȓ&1d5a��K6ʄhǣ2f���ȓS��(�6E7C+(<��#]�01��Ob�i��)O-E�[��E�)�\1��^ *((Gc��l1���	S�Ȁ�'%L"=E���+P
	0����S�t�(`���$ӉQ!L���O"�Oq����0敉j�&i��Ȍ�ME(i�S"O��Rq!Zd�J��̈́,���"O�����8=\8<��.L�M� K0"O8�/�$A��*�����q�"O�}g��E��ɉ&�́_�v��қ|�+3�D:���N�ڰ�"�
y��r�iE-R���	_�	̟H��O�aJ�G�6z�Fm�0�ʅ=��-�c"O���c�xϬH#�-FCyZ��"O��9�FE=9�(	Q,P9���G"OT�b��GӀ�c�YX'��� �'/��$ێ��eʗ��"v�j�J6��$�ў`0A?�{�V8:A�[��Xc_� �����?)	�>fl%�a��()(�Hǂ�f�j��n5���#�)R(8��nF�c؄�|��auf�� �(v&D]�ȓ^��Qz� I7�h��F�B\5��G�*�'C����3y��19C��I��$��/D�"<�'�?a����X?�V``#�[/BVy�R�X��!�䑖A鬩A��Ǡ.D�5o[��!�D���%	Ҭ����N.Rc!�DDrB,)gbڑ~\0��풺�!��]�X��Z�e\>Gm��B�L�4(��(�HO>�ЊI3)�&��@ǈ�~��eh ��< �`�`�O��`����]<���I���ibt2�F3w�@B'fS�Y5J>I���?��K�޴��6F���%�����!dF܈@q��r5 ,Z�M�7ˈO���* G"���
q�x˧u���������J���a���D|�N��?��͘OU(GߤT��d
�"B����)OT��d��V�>@c�Μ-��P��F�z�}2��<���!�# R^�i�5m�Dy"�
�yB�"
��i�OșFc���Tͱ��@�N|� f��O���i|k��E@(Vo��)����H\B�m�w��) [��Γv�l%���M�s#R7�蟜1:�ᕔ}µ�U���z�<�A�9OPEy��''����tP^��5�K#PȖ�iSk�w7j���1�NH[�OƎ ���`q��]��iF{R�3�i.���I1�Ԛ�ۡA��-�6�?�����t�i�t�'b�Q�x���!�ljD#ŜA
1T�_�I3�䇼u9����M>�0�O$��቙h*�� ���;���!*M�,������M;ES8GSؖG\i���d��/Kh�ɷ�˜=Œ�ʂ(��:���8{����O,��)���|B�o֚ex
�:4NL,S�ƹ��R[�<Y�U&G1u�vk�'M ����̝՟����4����9��hM �qǔFP!6�P�@�~��nr�d�O.�OQ>���+e�yh�Fȫ$���j��!D��"L݀S�����o��	���<D��`B��K$PPő�YTh3��?D�d1FaP�?a����"O�d)zi#D�j�cL3��������z�L�<�I����'�Tp��c��l�� 탺?DV-)H>	���?�Ó1��@��ŉ`���&�.i^��ȓ"&�,:w!R�I��L��D��0ه�m)���eOW.5y5�E�0+���ȓ�@A"�����ZF["�\�����򄕲3��9�Gܗ	��� D�ՑP��O�L���i>����]��y����Nf8J-פCyR���C<��OXi���s�Y����A N�j�<��Aڝ"Rh��,O�&�
�	2�_b�<� \ݹ�� �y�:��7�H<|�J�)�"O �q �jX|i�fMS�� [%�I�������$ I\|���ۡ6>*�"�� �O\�	�OR��)�$�"n֐�V�ҀE�μ���0<B�N�"�hT��pʰ �9q�B�	5-R��G�ȃ��䨅c��p��C䉛9�bx{�䙣SUZĘ�N��~��۩E�u	K��J���1�L.�ү#�S�O~ �G���A�ba)��ǚxt"t�B�'��4���'�B�|��i�
^/�[g.����v��>7�!򤉂C_�DK@A�#d���[�B�!�d$�|܁��ìR^�W�>�!�ݲ=��9�ӢYN��.ȯ+p!�� ?��ɡS��*P�:Mk2m�b�2��'���'2İ�M?I�-�3M�2%�&$��͐Ci?��O.�d�� ���ҵ�7��|
Q#�T�\��Č��z�p RtLU{�'r�XR�_a�|a�}��5PX(�f���ȡ)tǐ\�'R����?q��?��O_�U�F��X��YÄ�Z�2�u���?A���i�93+�;���P�,��#��Z�\��I�>ג��EĊE�h�A�� ����?���?������O\ʓd⭚0�2YJ�r�-���
��?Y���P=ԍ�EPl��c�BP0�OR6m<��6��O�"!9U*�?�$�f�N��a�O6I��O�-�O�s� ���)l�$U�6Z�"�B�r��D0�R�'G�'ȶ]jK�4�I|B��?���dm�*:gl��#�^F?&�'pl��W��y�'�11\�iW̐�w����@�ək*h=�L��3M��@QG"}��~�1�,e��c��;�0�j�'�ß�jf*.}�"���f��"F^0@�xb�h@�%�`�Ol���>	D�>)!�IN�D��U*����fE^Ī$i%*�-�Q%�<)��R[��Sg�Of�) �DU�����&lî���&�����n!}*��$�	\��I1-��$�3�4%�@r���1cX�"��Ry"i�����I�H�U��*�@ �'��jRy��'����<�\��9O.���O��A5���=��lݽx����'ԅ�	w�v8�Fk��� ��(i�B�	�ϐ�`�I
�*-�t�\���7m�O*�Ob��~�+��օJ8/�d)����=l�\ł��0���1��8�S�M#;�Fu[�@2X	��� �y���`-���� F����ͨ�y�������e�4kf��b
��y"�]E�AJ4��/=�ر,��y��q��"�3��=�b�:�y2���A���
,� ث��V�yB�݂1�.�bV'�� E6� PO��y��;�>�#L]%g�^��'��:�y��]�jZ~�H!4L�.xF��y��jT P�`� z��c��Ĵ�y�d��?��ԫ��ɗu5�5U�E1��O����O��$�O���؟h��+�g��B���	����g�����O�d�O��O��$�O��D�O�����\͊�o��t~XE̞ v��m����	Ο�������Iҟ�	���	=~ȔMJ��֎`�rCsE�����M���?����?����?����?���?��9j���� č�}V����ǣa����'��'���'��'c��'�R��!� �A�˙b��XC�jǹj�7��O����OV�D�O����Ov��O~�� |;l)J�c͘hG���A E ���mZ������	���Iԟ��ş,��!E����K���aQ(�:�p��4�?����?q��?i���?���?��ua2�#�朧'����"H(3��µio"�'�2�'�"�'���'�R�'��X���w���i��^M�(BiiӴ�D�O��O���O��$�O0���Ol�AL� ���#�"|*� b��̦��I��	ğx�	����I՟����L���:;`�q��1g,� ���Mk���?��?��?���?���?�B��p�SM��ִt���Bћ��'r��'}��'`��'gb�'�r&��.tz�hQZ�r8~�aqm� E��6m6?����7�CȔ�[��%`ֈ��IAS�܅H�O*˓�?	����t���	�a�p`q̏ d�q��~���O���f}��r3���O. �SOZV��E�V�O�C3ܘ��'��$���:$�i>�͓>j�	��`�/"18Q+�!��T2T��$����D4�� �"�e�?}6=�ba�OlV����Sj}��'=20O�S� t6���J��U�ᲄ��J(��?@�^�o�l���$����ܠW1O�SԺcߔ)ّ/,e���P�x�'���Xʡ�_�e��@ЗK�*>�=��m�O|-�'���*�M����O�Mc��RH=R�o�!�bP���'f��'��+ʛ+��Ɲ���'U�$��.�CT��&?���K�-�/� x�t��Е'�1��)��I�7�����kǢjK��P W�[�O���?)���g)Mx޹:G���*�d}�t�Ԇ;���?���y��)�Q���[U&��F���U*�7*�.�b��X>U��IɟL���'���%�\�'a>Q�c��R�&�ye@��)zY�@�'G���y�䗣tmV���b�mqc��1�?��i�Oʵ�'}(6��ͦ)[��Y�`ؐ���H�Ep#��w�L�G�¦I�'ot���?�c��<ﾘ�ŗ�m���Vꏑ[\"b�'Y!��ҵ,���掀�n�{���`r����ʯO�����DԽam~�c�J�.%z�ôS8l@O
�lچ�Ms�'c��x�ڴ��D��6��YgA]�^��`"�+D�-"Z� �?�%�.�$�<���ބR��h)'Q�W|��d��U��O���'��Ɵ�OUb!xƵm��*H��< /OVH�'��7զ�N<�����׋R6Yk���p�ɯ5~d9�j�;D�����S���?m�c�'�N�'�h����ŪQ3i	 V~l`�0�ٿ`���,�O X��dN  Y ��Cj�԰��'O��'-.7�-�I�����O��QJ;�U2p�U$k��2�c�O`��ݔ$wr7�,?����L��S~�T��.���� L�Fԉ�w��?�*O��DV�Xc�c�+%�M���G7�H����O��?1�ٴ�yB���2h�="ׂ�;vJ[F��D��V m�̽$��'?��tlZצ��M�\5Hgv�|���ӖQ����I�����'�<A%���'Q"�'L��٣̈��kP�يix���'���'�S�XB�O4���O��DZ�?`� ���E�d�Q��]-���xx*O��$f�`�%�<%O7X�(x��JO7OA.@�J�O`�$�76�^�#  �2�˓��!o�O�@؞'c�U�%Fx�Ԁ�A�Z4L2�T���?q���?1��h���	��0 ���xN ���l�����P}RR���ܴ��'����P,F*ճ���
w�A(o3��2�5����g�rnڀm(�n��<y�{�,�#�h1��=#���w/�?kzp��(�����O����O����O&���z)���� @&\E��nȤ:� ˓��IП����l%?版�4!d��Z�*-K���1:�AʩO��n�"�M�x��T)\ $T֍F�٣-}^p�q
K���d�qe�?���(,�B�+��'c��&���'�j`3�n�]���V���a���'���'h"�'�Z���O:���^�(�R
Э$l`�RHƳ%u&����?��\���ܟl̓u�^�Z�o 8ޡ�F�����jW����'j�B@@��?��}J�w�4M�EF��~��*Cø������?����?����?�����V��� 2n-� 7J5�E)`�'�'����?���ng�&�dB30A��P�'��S'aI y��'v"�'�2�����t����r���RƟ�cL<c�ϳS*]#��'o�'�T�����'���'�^�a�*�
t���\5.��l[F�'�B\��˨O����OH�$7��i3�|���PL)�jyK�>��?!N>��رؐa�D;R��T,��$��`�����A�u"�	��D�^}��"��OZ�9�L�>��Ig.�3bpd�F��O��$�O�D�O֒�\�'C� fPl��U�Ap��%� 9�?y.O��mj��Gp�	ş�:f���}~����?Wp�E͚۟��	�ywV�m��<���{����基��'���b%M�3�����HU$'�ޡQ�'T��㟀�	ޟ���h�	g���G��,z��R�:���A!o�	���	� %?�	�M[�'[|�H�_�y*DOPur����?yH>��?y�0Z4�ݴ�y���ܦ�؂�ܻf�blK6IO���m
�-uʭ�I�d��'w�i>!�	0VN� �U��+	�؜seb�&c\�����	�h�'����?����?	�!Q0IU$L{ ��B�LԾ��'���?I������f��4ds�&H?s��I����?Is�E�l��}ˇK~��O����>��D?n�(��Wkb�g�9A�R�'�r�'����<)��A� �ZxIe�Õ�@����{�O��1Ǜ�D��Y�N z[X�Q���X �`�/�O����O��d�U�R7�)?�F� ~#��I~�mHb��DC�T�� sy�%��0�d�<9���?���?a���?9��M�W&x0x1�����;����M_}2�'�B�')�O��%�b�<��T�R�%�Q	���,O��j��V��O�O���(�)Q�a�P=(�f�m�уF U�;\�ct�΃���U	n�5��O
\O>!-O��(Jk�hk�-��JXq qI�O<��Od�d�O���<��S���IJ�? B��U�ٱnՆ�{0��~l��:T�'Κ7�;������O���O4�R��H![���͞S�h�q)?]>�Ɵ��J ��L���A�T��鼓�bQ�Paj��t�ͭ;eP�ؕB�`��џ���ğ@�I̟�E�T�H�+���1%^�V*��P+*�?����?�Q���	ԟX��4��'	�s��_���0-��h�h<Ã�x�Cz��a���|��s�p�=	�#����F�2�0��ķP~=Z���cX�dR�������O:�d�O������pBC!ܭT�`p�%�?<?��D�O��X���ɟ��	ߟ��O2
�� A@�H��eK�'+#4l%�.O��'52�'ɧ�����96σ)_�}Z�BI�t3�� MP�<�awU���ӷv���W�6p>� B�C$T���9�.��2a������ҟ�IH��Wy��O�uj���:LD�\����n��q��'.�I,�M���>	�g��(����ഈy�#u8j�Ù'�& X3
������`瀍qP�4��x�Dݡr��D�1z���
�?1/OT���O^���O���O$�0�h1�b����� E��z�O����O.��=���O�!nZ�<Qwl�.H��P	hafU���U7�M�"�'U�'=�O��6�i�$T�P�J[�6'�y��#�$9R��u��P�I$+3�'��̟x�I1U���v[�t�
��3�A�"���។������'�(듁?a��?a�OͅN��R�ѭyT�w&B#��'��~�����O�O:��Dm�c����� �R��!�<I@�7f�r0C�� e����y�E( ���P#g��r����w� 8�?	��?!��?����o��$��Eg�)��nOh7�q���O��'�ɓ�Ms���On�A0�Hȥk�dX�#���D�t��'��6m�̟�oڳy��nv~��D�\��3�~$R�.��J���D�2Y��0&�|�T���I��l�	ן��I�x��H�f�@P�8� ÆA
iyR��>Y���?A����<��aY:��z��AYE+#�������I[�)�S�Z�pt'ʁ-/�D%�����=܎����p�`�i{�A�OD��M>+OlE�q�O�We����J�?F9��8E�O����O����O"�D�<� [�H�ɛT!$����Jgyr�Og0�E�I��M�R��>1���?ɜ'�������)F ^���n@��IX����M��Ox&��'�z��49V@(��8r�M�e$��7�'t�'�R�'�R�'U>Qٰ�At+h�%N.68�%�O����O�a�'���M��y"#H�&8@�鑁0-����6���?����?�TA���MÝ'�rMF�h>V͘V`�P5��`Ԇu���rCB�͟���|RR��֟���ݟ��딺C�U�VM��6hr��Yʟ��I{y��>���?�����i^--K�l�-ފl�eb0�R�f��	���d�Oz�$)��~�dV�C����A�g�zA�H fՓŇWۦ��/O��	�,�~B�|�ш*W�2�d��6�,� q-I�o��'U��'����d^�`	�Z�e���N��EcG��5�z��	��h�I�M��ҍ�>�N$�Y����+Vَ��j�7_=��x���?�"h��M�O� i�
���d�?�Ȓ�T/d*�Qb-_
q���7D�ON��?Y��?y���?�����	ݬ��$��V�:�<5{w"���L듟?����?	N~Γk�f<O��2����Q�(�GF$��qs�'���|r��tm�"��O����+;�Rb�ϑ>�a2�'��l���4��|2[��՟��+�_�8�ŉ 6|(�4�ٟ���ݟ���My"#�>���?A��8�r��@ ڙ^��9�f�^�<(���>����?yJ>�0��=�@X�4'�0]ؙ�!��?�nszA��.����'����]埄�1OI�)] ;�V�gB�V1� ��'���'B�'��>��Zc���skݡE ��@�uZ0�ɉ��d�O�����?�'��)eOQ+|8���Hͺ��L���?����?�r�ˣ�MK�O4<R���8����
�M&:�[��!�r8ё��9C/�'��˟���ܟ��Iԟ����e0��kq�6���WM
?V��'GDꓸ?��?H~2��Yh&ʵ!�azv�H�B�ปqQ�,��ӟ&��S��$�m�,��DZ�+�^ 閲<a"%xV�Ϧ�)-O��	����~|�Q��J����?iZ�hs,R�~X�A0�IIן�Iǟ���ɟ$�	MyBj�>a�Ĥ{ՂS%!�D�&�Ź����)/���dTK}��'[�9O�"��ɤ s�%2���B��U�V�_7p>�����V[�o��i/��s�8�"J&N���8�A%',-�� �O����O����ON�d�O�#|R4e<:�� �	!��!`
�����؟h�Oz���O<lZD̓ �P��9Mp����y#��&���	ߟ����^M"QoZ|~2+�B#�4ij��R��W�u��
�
O�V�&���|���uG֟8���O��d�wa�ar<�xͻQ��lKV���O��{>�I韐�	���O�4�A�f_�?�f�1Ed�Q�������?����ģ|��B�~KP��%fX�1PQ.8Q2�Y�Gl�0z��Çŝl~2�O��5�	9Y+�'�n���IK�5�ެs�$�=~�����'���'+��'�O�ɔ�?� �=ؤ�1+i����g�*b���'���'��7�"�	����OD*��ۯ(F�S��W�_�$�J��g��nR	�(n�]~��ך���S-d�Ӓ\t��˷4H��Q�+�,5�4��<���?I���?y���?Qϟ�q[nׯ��y;���0�&x�v��>	��?�����<��i�R<I��|k�AG��{�+S>,B2OO��� ����q�H��^�"�D
.��5�UKҝ#���-/I����Y�6�O���?��OV����S�.�BD�գ�Ft�\���?���?�,OD��'��	럔	�VŤ �c���
� NX)2�:�O@�n��MkĞx�ߎT���%��	u8XUзo�*2��9��}�V��I��)&?�&�'��Γ} �@�ā�g���	3�)Z-�	ş$��џ�Il�O��$�&/Ö���N�a����]1,���>!���?�6�i��O@�I��5��+�LW��8�I�k�0�d�O$�d�O$�;�d��Iɟl�q���i�'e;��Y�l(�~hȵaN�Q���O|��?����?����?��2⮽�sDڼ̩TL���`�/O�P�'<�'~��4�'�x��1�K�����K�,&�3�η>��?�H>�|�� �U� ��uCN�G�b��欛\:��ߴi��5g���1�On�OX�[���@uH�.H�`��M'_OJc��?Y���?A��?	/O��' �[�~�����	�/b�0X6爗E�&x�r�|�OD�mڌ�?�� � X����3e9�!��/O�0W&t`�b�M�'e�|�Ъ��?�kq��t;�����}�|e�U��5@J��Ц�'mb�'"2�'mB�'�>)Gm@ D^�r�N4z!Z`b�'�O���Of|�'uR�'_h7-&�hH�Ņ�&c° ѕ
�C��$�`ڴ=���O<��*�i|��O�p�ƃ;7Z4���1'�ڕ��!�����\ڜ�O�ʓ�?A��?���	�1*��!N��,�{x�����?Y)On��'���'w�?mh��9
�}�1oO2M$UB�	�<��]�P��Ɵ�'��2�\٠I.!���w��<(��՗mJ��\y�OV���	fy�'U>сG�Z5-��Z �A�EHq# �'���'H��'E�Oa�	��?��"3�*��ln>�p���̟��'��7-%�I��DJ�!@T�Ԛ{�Ȅ`��B���2�d	�?�ߴ%����4���M=dp$y��W�h�'��ݹ�D#dX8�HUJ��\�	]y��'�r�'"��'mR�?��@�� oV�;V��^.�,A���[}��'��'��OB+i���I�|��4@	�<�R�C�d�x�l��?�K<�O~�T��Mk�'xV@J�ATp�@`^�$��6� ���O��8I>(OL�D�O���ej)_�4M�t�.lU�q��
�O���OL�D�<Y�^���	����	v^��p2�P2R�4|�R�K�?��(�?��W�|�I�t$��0`�ηuHf�H(^?���f�؟P�	�$��R�[�UP+O��֊�~26O�,�Å���zv�ϫ �ɹ1�'��'���'��>��.���F��J��$C��-(��������O��$�צ�?	�'"��qY	�Xaw�8�2 ���O����O�����5L 7�;?�6NM�I����`s��H���*���aA)~�H�&���'�b�'.��'���'� ��f�'C0&a���(���Z���O�˓�?�I~z��O;~�x$B��&��щs�ِ_�^Њ�S�4�I̟�&��՟���"��8+!Đ"ۢ����	��z��ݦ�,OH��蕋�~��|�Z�(�ED��N	NIc7_.v�e)v��۟�������	۟���byrή>��D�2�����P���]�dr��T��V�$c}2�oӰ��I�H�
]��la�ͤ\X[U��]�T7-*?QamD�h����;���y'�Z-o]��(�G�0r"�{��ݐ�?����?����?����?��IA�G29��'$.�Z`��W"�'|�%�>!��?�iV1O 0:����[CBaCW�R+i !�V�|R�'	r�'����iV��9 ������;| �ڃ�a%�ػ��R�P���7��<����?i���?�!��p��i���X({�
d�qO��?������On}�',��'8��*��7���(vRx��_-	���'J�ꓢ?������|R�E�h�zԎݪdל��`Ϯm}X�
C���jW�-kܴ
�	�?���O�O�o�x��F��^�2��Q��O��$�O��d�O�����	�NJ=9���ӳ�a3�( �'^ �?���?��i��O���'r�G"_��`*�Nץ�L	��o03�'Pl�
пi�	�9�
��5ٟ��']��(�.
>��$�f�s�4I�	My��'�r�'iR�'��?1U	Gn��u��/�&^V%���XB}r^���	`�ğlY޴�y���
c�1J��� `��q�I:i���'�ɧ�';(��۴�~��G�^�j0�r,d�K�iD��?���%"b���<�䓤�$�O0��Qoy��b �U����4IL�K�����O����O�ʓO��IX�I�`��ע�M�Ν�N2���Mj������M�5�'��'���� `ƅU��mY�L�Su�$S�܂6�i?-�����':�䘏�y���X��4�$ �&��(A�7�?���?!��?���i~�� h):�'Hg%���=�<����'6��?1�����D��|����]�n�ٶ�W�L1�IA�j�OZ���Ox��6�&7�"?�![hSX�S��L%�lN�,�
���� :�&���'���'Ir�'���'����ۆAtĘTi�.�,� [��`�O��$�O���/�9Or�sq�U�*�e�D����rCx}R�'�d5�4�����dt9���+��D�2�ˡ%Qn�8d%(^����<�ѣ�O�l�D�����N�z�08��U(W��!��Q�1w$���Op���O4���O��{%�	�� � ��:�JD�"F�: �8���ܟܹ�4��'��ꓼ?q�'b��V�:l�E��P=�� �'lz��8ߴ��D�K������p������ӲĆ	L�.���8�x�d�O>�$�O��D�O��"§cl*���-]�4��|aE��3�­�Iʟ8������OP���ڦy�<)d����`2����A�T�A������� q�\��%.��7my�,�	�B�H![�,J�r�"��C���X�LJ�� $�R.�o��Ay��'+B�'.",5�tl鴪X�[�%pֈ�;d��'��	3���O�D�O�'R�8QN�1l�|��E�
`ܗ'6��5�v��O�O�	���0򧏎zD�łX�.���@EZ>�1��I4\�������OdI*N>1����C��L0�8E؊ȱ����?����?����?	O~r-O@��	7m�hɺ������A�G+��Ķ<���i8�O��'��7�F)#ubp�RD�4nc*ب6FB(st��n��M;d��	�M��Onx`V����6#ʧ�� F:1�sk̥)�ސ�`�H� �'���'���'{��'S��2a���U��^Z\�b"�!Y[V�'��'U��)ᦩ�*|�M�Bk�RZ�l��,.�D�O�On���a#��j�b�I3S�v�*F&��q����B`�m1 �Dרxd(�8��*$�O,��|r��FM��0W�	U+��h�
f%��!��?����?�/Or��'���'h���%/��k��?Kͤ�s�a�)OD�O���'O��'��'/N=CaQ�!Քd���H2�����S�PSҦ�,'��L�#�9?�'\O���3�y"/C�	^�;�H0�� J��<	���?���?���e��0� �i�D���O��v�D]CE�Ob��'��'�|6'�I�?�(d��$!�4��a ��+����G��<ڴg?��j�~I�S�g�����t�H�y����&Fu��B�	�b"�+5H*Kh�$���'��'w2�'���'��dhp
�>��1��he�`�BwQ�l��OJ���OX�$3�9O�\�Ȇ?\T���ܾn�I �lBu}�,���	D�)�ӽBn��	�e�7(NĘ0K�(��-�Ώ�@T̔'�l�`w����li��|"Y����� IF�e�PN�6T^�(��MS���	ӟ4����X��Ty�̼>���+ۺ�����n4��j�N4&�E���Ex�v�d�^y��''��'�V}"�w,)I�&ZV4�C��p�����P��V����_���C�H�6���:��ea=���⟐�	����I֟t��̟�F�D��=p�p6��*�b����Z��?!���?92^�<�I���ٴ��'�\ G�`&&<J#�@�����x�bt����X�+�fr�b�
�(�����4Y��I�ek�$$.��(���䛴����D�O�d�O<��R#Q��� ��Bq��aCgǞO��d�O6�=5��yR�'1�ӷ"����ꙶ<_޽;Gb�~tʓ��I�x�	q�)�BR�NX<|��d�=K�t5���٦:$�Zb��"
A���'��
	ӟ,ir�|"j]c��:��T�Ve*�䛳*�R�'�B�'���D^�h*��t���3�ۯ8-Ĩ����$l>�\�	���I��M���>���i����墚�Z8\xp'á�]r��S���M����Mh�OT\S+D�B4'"w�y�4�����'<�\XSAПd�'�"�'z��'�"�'-��Q���'�V�5�
�Bs��!.:���'��'����'�
7g�`s1��3 ��r�;$ĥQ����*���ē��'&�8���4�~�쉚k	����ʧ\v��+!i���?����4����<�����O����??.�(�̒Bಽ
k	)~�$�O����O��s�I�����PDG�^�����\�yo�`�K��	��M{�i�vO�l��錳���fD2�����)�O��DC! F�C�Q�;"���r'��O�@�'��x�W�Հ@��@��Y>E������?����?���h���	(Dv�p����-n�Y!d��f���$�D}R]���4��'�����;y��T ��-W��˜'�R�i�
7�F.W��7-0?�U���-���i͏w^�ć���z]1-xd�ө2�d�<����?��ӻ���Ov�D�"��غG�*(F���jE'|�C��IJy��'��L�Q�LA�|��Gŀb�l0�]y"�'��$#��šmS�pI��:G".����Tn�ԭ���O�{��ɞS��)J��'\�&�,�'�8*r"��p��#+)�41;V�'���'m��'P"Z����O��I�X�ty��KG�a8�,����i����צ��?��U��	����KVH̲��Ӻ%s±a$��v�`q��J����'ص
��TO~�w��9f/�s	�=	f��7t,���?���?����?������ �\�����2z��!΁��'��'�<꓄��Ʀ��<��D6�챒��3Y�)!�@I�	�(��ɟ�`�%�����''2� Q��xd��0�h̡6͔�Y2�4!�xa������D�O>�d�O���H��8��Q��+�R���Z>'H���O��K��ҟ�I�X�O�>�. ]�1fI��,�,O���'A�'aɧ�/O6�0S�S�V�lc AC1	p(��fC��(�7�oyR�Oe������3!�H�g�Kp��	;��q������?��?y�����$�۟�%�
쨻����`A��O��d�O4�!���O>�M����:h ɸ�O��?(9Pc��?�4�i�DD�׽i��i��Q��A��~�d��@�C}Zc˜�ɄD��zB0%��[2t�q������O��$�O�D�O���:�am�7"�����B�Q��TOܯ��D�O����O������A��ϓdޱ��gR�Yt+�Nʼ��B�4�"�xr����D-��&�O�D8�k!2����׌�2�����'���"�i�ߟ� ��|�Y�������f_�3�ؘ�7��f��X�w��,�	֟D��{y�,�>���?1��@DR@ᦂ��m��-�1,����*�>ᵲi��7-HG�	79$�{Ŋ��a�iqT�Ub�I�'^��9�')m�V����TF�蟈21O�遗��c,��Ӆ�hg�����'��'uR�'��>�Γo@"� P���gy:`Y��W!!2������D�<�ҽij�OF�I� #*(hӤ��iE!O� �
���¦��ܴ4G��M��D�֙��9r��;�c�a�5��l_�EH���b⋄*�M%�З'R��'b�';�'$�x���sM��&�-\ 6�1wZ�0p�O���O���)�9O>�3��%a/��0#�/ ��Bˇa}�JmӢ�n����S�')z�u;5�ť�I8�m��q�����l�&CV��)O�I�C��3�?q��'�d�<���'*�xk�Q9~����?1���?��?I����D�]}��'�����3e���8�k��D["�'%�78�I���G����4p�b�V �15.J�:����,J�Z�y�4��$[�e%�U8��JvX����ݍo'ܸ+�GUຐ����+%�X���O��d�Od�D�Ov��1�'ȍ� �.-�<ŚP��q�T���?���+{�I�L��*�M��y��T�a�U`O��֠#գĎ�䓥?!���?�$���Ms�O�:�� g>>p�cK�2
�\�*��"��R�'��'����������	�Vyd0�%���-Mt�y��@�b=���	Ɵؖ'�듎?����?�Ο��YW��Pj������QCP�<��O��$�O�O�)�O���捅�??�D�K� t��x� <Kނ�F�a��'���Hu?YL>�vf�P�&��D��# }��[#�װ�?����?���?QO~j+OV��� 5�d��S?#>��0�������<Ųi��O���'"��I���4)�P�~0�D� f���}Ӏ=0�x�z�J�"�1��t`̟xQ"e�N��&��)�9��-
g�'R�I���	����������b��cQ�_��X�cF��TOJ9��I�yw��ܟ�����&?牙�M��'LP�W+��dq�`M:zmJӴi�h7m�\�	@�(+�In�O?�6B�-h�����? :�y�S(C����"O�n���_u��NyB�'�҃�W|Pr��[�EP�}�fp����?����?�+Or��'}�'�g�!��аq/V 1���zb�"�O���'��6��5�N<15(.�ҩT-N8O,UIsb)���P�u�������	D�������R�,P��MׁRJ $�pn�Qt����O:�D�OX�d;ڧ�yB�Ս0�<`G�i���G�A5�?!�^���'��7$���?��C�5@�h�g�%Fܥa0��Cڦ�z��M�s�F�Mc�O��o�$��!|W�H�ˢkH��喞(5��OB��?A���?i��?q��R5^�A�KԷ]Q�@��n�NX]�.O�}�'���'#���'��CgM��^�a�Я=�,*c-�>1�i��D!�4������rekt�>AO��AU�32�LA�b��m8��Co�<!	�9Mm��DP<����d�L;N!YC�K�$4k�g�?���D�O����O6��O�?��	��(bR,<,<\�r���
w���wN�ٟ,��4��'����?1�'Mra�- ��`ԁ�CV�¢E34	dUS۴�y��'�@a��B�?q�AX�@�ռ�����,ٺ�Hl&|0�PПt��柔�	ȟ��IܟXF�D��d�z|���V1�l ����?Q���?Y�W���	��4��'R�x;#n�����Z&NY�o\�X#1�x�n|��u���00�r��R�xk�-J�]�����-��Z(��
94l���c�n�O6��?	���?���CђlsdV_�(H�l��L(*���?9,O�,�'��'E�?�)`�G H��S���tR����<��_����ߟ�$���Ɵ�Y�	��o��9#�i��w	v���O�5؀Uh����U�)O �I ��~2�| DF �Ї.Ҫ,�11a$6��'��'T��dT��������#��7_�8��uɖ?�:��I��t�ɲ�Mk��c�>1�i6���R/qP�H6B"w�a$)�O,7m���7*?�f���$�P��;���U)���s@�R7yNq3��3URr_�8�	ޟd�	�|�I՟��π ��",�*3D*�8UiD&l@�qCEG�>���?Y����'�?���i5�䘔X�DE��2_\`qӄ��k،7-���&��&?Y�ӉG�����
cX�!Fꝫ;:���a�ۡ#����b�ޅ��'̼9&���'�r�'4�=[�o�=db����	8
h�ذ�'���'�RR��+�O��D�O �������
Ϡ���ОDj���ɫO��m�	�?QI<q4JP� Mf��1/��wUh�Gɀ&��DǼ��+�
%$�����{�$���"  �����Hi��Q�d�O��D�O�D�O��}�'�:(Q�*E>(�x0V����!���7���������M[���Ok�\����T$D�B��5pzX}���'�J6��ȟ0o��xlZW~b�Y;pp^U�S�q�2HAW�-Q�&XAjܬ8?~$���|Z����ٟ����D��֟��Em�L��f��*�,�P�NUy"��>�)O6��>�ӹ3<�9I�	��j�(����m$J�)+O��dp�`d'���r�H�쇻 ����O G3��2�$l�\�#��<�w����$Ȇ�䓋�Dͺ
,�qr ��?������Qv���OT�D�OL�D�Ov˓U���ş�'K��`���C�7l9������4��'����?)��y�m��S���ٲ	�,��{CM�:*H�޴�y"�'$�	[GI�a�*OJ�)p��"�BB�>����N�g#��pT��O&���O
�$�O`�$�O0#|�G��Z$�X;rkБX/
�cS��4����<��O����OLm�A̓]+��+�Fǁ1�*�ؔ�)�J�&�h�����I)m^�m�J~�kך3�*�0��6�r�ѐ�^�Ѓ���z?iN>Q.O��D�O��$�O�x�c��?os�P	�L�}אT� ��ON��<I�Q����ӟ$��R��W��:�qr�G�d����;���Wi}��o� ��a�)�4�@6��8��/�	gE$���2D�exq�@�'��e2.O���4�?ɖ�9�Ć�Ze�0�G"�+DU�=�aE΋}s��$�O�$�ON��/�i�<��'�t�hć)���6�
Q�����?��A�����P}Ot�R��'���JHބP�Y5J~�ts�ߟ�oZ~V�np~��]$vH��&?}��)	f�Q�]���B��/���d�<A���?���?����?�ʟ�	k�#ɠe� �a ��@��Ʒ>����?����O
�6�e���E�U2���vDGF�(��+H��=#���ē��'i��]��4�~�G�I�F(c����|-y)_�?�t(�7�����䓷���OJ���<����e��Ŧ���dˬu���O��D�O�ʓh����������l�Q39>�23� pU`��g�v�	��I� ��@�I3}<$�w'�#Q�(!`Ҭ�!&��T�'�De�$����F�;���~B=O�J��'� �2�C.L|����'l��'��'s�>��i뎰*�%<�D|pdJ��e�	�����<)�i��O*���oDN0�N���q���LRi0���O���O�ݒl���p���@���ם}�\p5BF�lCTۦJL�."�O\��?����?����?��5������]�s>Ap�@�0(|�{)OL	�'c��'����'dV3Q`_�]����3�ܼX(� "�>��i��7M�E�)�%G^b�)э�9��`R�Źt��CBՇ��8�'��J$#�ȟtS�|rS����|�l˱��<�F�I��@��	�@��ȟ���`y�>��A�0�0w�g�B�*�㚶��Z��-�v�|��'���=�V��OH�DN#[o�@q�E�:�z�ҽK���W�i���On@jv�S����ƪ<��'�y��[�E����$
�J�"��<������I֟���ݟ��Ir�Ov�����ɴU�(yi�i�G�t!.O@��@u}\�ly�4��'�z�A�%D�mR���Y'T*v=�@�xb�qӲ�l�?��&'�	��?�P��q���A�14~p�����H0��O�hYK>A(O����OH�D�OH�dl�\�foI�%�Τ` ��'_�I�����O����Of�';H��Y0aN�3����j̆&�)�'����?Q�����|"��y2��>l���	�@�R��k�F��4#(���?�v�OB�O���U/�]ǖmra���Tzf�$��O��$�Oz�$�O��B˓ccҨŀ]$(5
���KZ�p$ɂ�?����?Y��i��O6i�'k��W6N�p�����5��9QM�((�"�'zJ�ҽi���O
�xWo[����]�j�Nn�Xه�ͤ!�Rm8@�AɟL�'��'��'v��';���,n��N^� ����S3J���'���'�����U�<D�І솱J<�9�#��ch����8'�<�	��D��ly8�o��<yaS��L��E%2ྈ��N�?���$I_���������4�2�dɯcע�S��\�\����1�8���O��d�O�ʓF���t��ş<#����T���ګb($`SNx�(��2�M���'ǉ'��E��Ȁ4R!F�
��؇Y(�R�'�bg�p%���`��,Z���?����'�hAϓz�(�c
Q�T	���q���r�@��П@��ߟ��	a�O����'��r����W�����>9.ODmZj��Jeb��t��Q���R�95�]�?�W�i��7͞��ؠ�Φ��?	eΈ�]v�����|��p� �)j4H���6�v@#J>�,O����O:�$�OJ�$�OT� �i[�M4N�xi�9�T�uQ��I�O���OV��'�9O�(S�A�5�U��Q��� "�
B}��y�*��	O�i>��S�?�y��P#a�bUa%,�-s�Б#c�6k� ��AWy��#~¦I���T�'��IWl��cC�*5lTH$�?A:�	ҟ���ȟ�����x�'b���?�Pƃ�5�RI1C�ɭoT�0����?���ib�O�l�'�6͐�ɩ����l�:(h��G5d$��j(j����̟����Q�4�py��O5��i|� ��xt��7���8!��' ��'��'(���,O0�� ��&(����5lx�D�O��$BR}�V>��4��'c�m�e�;a��`�(h���x"`v� |�韂��1)h�L�*c�l�B
?�n}�EȴN
�;w�2�ח�䓟��O��D�O��dL0���@4���w�$�cŢǂ&����O��>E�I�`�I���O^�۠��5YJ�� �֧+),O� �'�R6-ן�&��O�4)  �~�
l� $+	Q� [���ɳJA�����N����<�OH���`��\֖l�G�Οf
$�M�O~�D�OP�$�OV��j�uv҈_�G뤤y���6[]�m�G,��?Y���?i�i��Ozu�'�7mU;M�b�AA��-4%8В���x"(��	ߦ��!�K榍�'���"Ri��?u��~�h�s�8U{��1���2.�OB��?)��?����?���i�9�4+7LӴ,V�L��s��?����?�I~���@j�&3O�A��l�0nE�)�s" �T�٨ �'OҔ|��d��5қ��O�$B�%ې`v�:�#�>P�+��'X��	�������|�W��S��9���t��i �?�@�V͟T��៴�IVyB�>q���?���H?ļI@+H�-O�ɀ�mQ�PM{�"E�>I���?�H>I�I�= 9;�MO�J�C��O���Ą6'~���I7:��i>�  �'~ֱ�RS�D��<v<t�g��H�2H��ßT�������N�O �$�(���pb�׭ ����D��"?��>A/O��le�������l5̪0�1>`�����?����?���+��!�4����<�C�'�uw�/\��%��M:>Ab)�mB�����D�O���O��d�Oz�S�"���"c	-|A�S5��9\\���������ӟ%?��,r12�T��<�$���K5�~�1�O����O��O1��=�7G�Q�N�+ ����bk��?7�0J��� ��Ɩ�{2�i�	kyr
�*����.	Y���{ƤH�\��'���'l�'��I���Df�`��")s����Uc]�([|�`Gg�O��nZ]�����ҟx���<ICE�/t����5P��M���O!o�(�lZP~"�N�?�@�Sxܧ�y�B�;$R�B�L�i8B݁��<�?����?����?����?I���F_��T�)� �v�B�'�r.�>�(O*oy�M�x8"��$6q� a�-��`ZB!$����ğ �ɞ��ml�w~@�1�:��D�J$��!H0�G*��q򦄓��@�|�T��S�����ߟ�S�
�<���Bqf��}pҴJ�֟x�Iey��>�.O��$5��Q/����*H��Р#]Qy�D�>����?aJ>��Tu�G��cN��)�_P��z�BU:|�������d� 4H�#c8�O$��S(	;ܘt�+���.81��O��d�O
���ON��B�3�ү���pÀ� Ȝbဇ�?���?���i+�O `�'���� �< C�͒�N� ��A�73��'_�1d�i��I'�PU�d�OB�O�ұ@�� _ʦ\2lG.4��!x���$�O��D�O&�d�O���)�ѭǨy�X��.	�"c8퓲d������O���O���dԦ-̓C>p�Ə5%!bA�S �~��	ǟp'��'?�`Pʇ���=)���
Q?c�t�*h�r2�-����;��'�v(%�ȗ��t�'Z�mf���a�t�a�d0cJ�?Q���?a����d�d}��'A�'��V��-�b�E��#�ޥQ��@{}ZT��l�O@O��2�MѬp���רEi��&�<)��oӰ����4��O7���I7��Jb��"/ t,�ga�w��4�	ҟ$��ןX��y�O��Ħ?�v�Ӳ��&[8M�&�����>���?�"�i��ON�霒�0��Y+��t�o�"]�X��Ц�y���M{�B�2�M3�O�|��O���r��'���rq̒s*b���a�.��Odʓ�?����?���?�9,�d���%-��0����a�5�/O~}��'���'R��y2.T=*�)i�A�D�&ř�cyUF˓�?�����S��xrhJVɝ6-������6�2���\�d��H�'����b�ɟT���|2R�h뀅
)�^�*$� F�xp������<����,�IGy��>y���P��F�6A Z0����0O� ��Sn���
[}�C}�5���l!4�
m̑�K�^"�@�W�W7m:?	O0^��D��'�y'f�XX䀵����,:!����?���?y���?9��?����d�pQ�g�+y�]	�Gr�B�'qrk�>���?Q��i�1O�Ńg.�i�`a�S+ҷ-����9�d�O���O?����i���/ey���S ��d}{�˙� 4d0���J�<
K�u�Uyr�'�R�'"� �0#��S�c����GnQ�;��T�!�'D�[�ԓ�O����O���6�aƝ6ިaū�4
F��My2˵>!2�i�~��-�~Z���'PZ�l���i�b1R��
�5�,a����3lć�' �T �՟�1��|�ü5����WG��/|����R(���'W��'�����U����5�"}K��m��2�썠!S���I������M[L>9�S���ڟ0r�a@-J`�g$R�d1�ht�G㦗��A!���=�'> ��c�?1��?Q�C�g���Ud]�t�^t�!��O���?a��?i���?I������="϶�q�ۣ����bB8R��ꓒ��OГ��$YĦ��\���L�<��	�NT*o��؋�4x9�C/��.�i��b�~6����R�*a����0�����O詂\��?9Qa2�$�<����?���+B恨��!i�๨#�e���O"���O`ʓpK������	���"���<q#ޥYd��f�<�C��Tt����dP�O&�$�O�O�=҄-�2Z�"���(B�u�yf�<��+ʢe����4o��O����y�x$��e� �jD��g��"�?���?���?����v�����F����j�,b� H*�,�O|��'���'��6�6�$�O���ֲ*��� $2l��Z�-�:��ɦ��ش�VhƋm����|Ȱ*�2u\��W��9��0�@]���ǲz��&�X�'���'"�'�"�'�4���(Z�f���+�a�-UL2cW��:�O����O��?���O�p[���+A昢ÄۡJ��J��w}2�'���|����(��3�֜d]V��2�J�n���!ոi�V�qV"t3�篟�$���'#��˖��8AR��,�j� ����'lr�'���'�R����O6�E�jc��a�H~5Yr�W���DT���$���ɐ����O��$d� j2�hդT�`�~)���6*vD6�7?��"9�����ؼ�(˺�"P(Pn�"��U�!l֟��	̟0�Iܟx���HE�t�.<�36EҊ*��*��0��D�O���'""�''�6+�$O7NSZ\�r��8X�x+\H��UF�w�I��Mk!�i��4D�~��f����f`���4@q��Z�Ը��P-���ʑ�'b:'�Ж'�R�'���'N�����~ ƀ��	�r<R`��'rV��9�O>�d�O`��&BqӎR+B���4F�<@��iy2�>y��i�T��4�~z��+�x��7M/1���v	��GC�)0#ξ~�Xі'��� ϟLc՛|�g�QJ���⯖�]Z*u2PF/z���'�R�'�ҙ�P�pk�9n���D֌V���a3$���I����I�M#��H�>A �i% !��o?D��WH�:[\�:�@�Ot7�X�=�067?ɢ��7'�������i	�A�����ÂRuz�#EO*u��[���������4�	˟X�O���A���0���¯�=�
h��\����ן���t�s�c�4�y�Ş�,�:M� �x���I��D�{Y��!�OOn�����Q�b���	�vx4hR�O�G��eٴ�M�&�ă&qp� �J�
�O���?Q�-u�!xk���9
kuAMߟt������Iay�	�>���?���kBJ���q�5����p���2��>鷵iB��D>�K!vԥI����)�Ƭ�#�̋��˓pN�jeF}/tL O~�5��OjLh�'}4U"'f�!P�t�% �h�I���?����?9���h���I1It �DAդM�(LYvgZ����s}�'���x��⟴�ӞY��Xb�ŏi�( ��R�ODf��ɩ�M���'�Fe$E����80 �7MK���+k��D�?l� �B�"��e�`�&���'���'���'�r�'a����Fo^t�(����E\���O`���O��d-�9O�4���^��5 �=���Lyy�'�B�|J~��Zhh��Eh�������0����f���DFB�{ WY�VH���"0e����4H�q5�ǰK���R�^�	m�D1Bd�'8-¼��hZ-9�y�L)P^���¦g�^%SS�=���c�9U�Vn�Y���tDؽ,(��U���O�����-�9JS��+B�ګj춼��Gr�<xz�"� ]p�
���<t�Ft�GK�8:�H��%�Ual�zqo� �V��F�Q^v��UGԶ!�.�s���"�����i�=��h�:9���@X|���J�=�@5�aM@�L�@U)=�t;Î9����`eNT�r�CȲ9�H=�A��
 J�!0��#H(��	ٗ{�e)PɀD	z��6�5w��-���[�4��X��'IVo���4ԉ>d���Ώpa����#[ߦ�i�F_��eKg�(0���	�tĉ`�O�u�v����/{+��ɰG���1��T3���M�WH5�Q�Юr�N]@�E�6)��ӡWI&��'l�b0�����P%#������߰N����FB�,$A$�"
\8t!�S�
0��	Ĳ�RY�$�ԇ^b��E)M(/���ڂ�ۨqD��9R�Yf��aj�V��OHx�w�Z;�I#d�)H;D�j�B�O��d<�d�O����aG�c��'iߎ �l(�/�\Iwb�ON���O|�f3O��dN���'���'�J�D�������O�X������|��'���ɪ@|��|�8�4�	�$?ע%�V��^7�<2��'�	�'���n���$�O����O��',m�#	��Ppv<�C��)l��=���'��'�������|"��T�I�D�iҤ9i����u��2��y����?�0�i���'���'� 듄򄏨i�lpÃQ
��Q����$�
9���O�:Uq�'��CȂy�����<#\d%�Â#�6M�OZ���O��d�P}�R���	�<14	صx�R��k�]Z����i�D�>���X��?����?�� B�i��Bd|l(���Ǚu��P�T�'���'�z����O��O�����
6;�`��X
Q��]���<Y0��?����<����?�����)�",M��S�W�=r`k�<T����>,O��$�<���?��xKl`�5 ����B��/Ro.���F��?!E��<���?����8�t)�u��	����?I(Or�d&�$�Op��Q8��I�IR	�&-]�\0��Ď&�H	bf;O�D�O��D+�)E���'�z `%�c�Fy���ե#e ���'�r�|�'���� %�1Oԑ�"Z8y�RU�eE�..J"����'��'���'ORL�~b���?y����d�oS�c(t,���ѥOKB��I>���?�v	Z_�'5��m��0"F$:�����m�pR&Ҿ�y��'o@7�O��d�O���h}B�EtN�:��f�P8"�G"^��'
"�2u�O$ʧt�d]x�&�"�@�b�nm��^��?!�Qw�f�':b�'����>�)O
��s�<��I�%.Uv8q���O"��A�<�Ii��a�<�y��'��09�A�2`�\�9�ME�!B���kӐ�d�O����O�t�'��	ǟ�͓V��)���7��(���L�9f��?)��ɴ�?��	\�<���?i��%x<�b*�8Z�����ĳk���H���?��t��	cyR�'��'L��@#��4r 
��!�&�|$�']�`�è�Ɵ�f�a�@�I� �	p�D� �N<aY�d�rp�,�T*�?��x��'�b�|�Y�����C�)��!�7.2nY�@������!�L�	���Iʟ�%?��� r�q��
> �KĦM^2͖'Q��'��'P�i>u�Im���JR	GI�@}z�d�)YN�)q`d� �I����g������OR��Ņӑ]i���W%���O��/���<ͧ�?)͟�!A� L�VZ`eX��݅��A� �'G2�'�$���'�Rn�~���?��wv�����V�D1��:"�M�<[���J>1*O����OD���KcL��5��y���R�P
K�:�$�%��˓�?����?)��?�.O�\jtÂ>P�� �$��02��!%��O.��<yiKK�����d�}z��ݟc��4���@�$��P�P���I�p�'��[��o���"�R�d^��2�M&UP�XC+Ol�"q�i>e�q�,?AF��*ھȹ���aΔXW�M��?I���?���?�-O��z~"�*0�����];΍�UB4޼�Gxr�O����O��du�9�fR@�*	SQ��#�f��$,�O8���O�˓��2��$9"�4�
^!=���+��_p$�h�b��  ���?!��|:�'ޔ]{�!�)A���p��K�������O �$?�I��ϓ6�ṱ@�-E�U �+��~���!d�z%�Kg�x�I���m����׀m��Y��ŏ�1AM���SQyr�'"�|b]��Sڟ��΀�$(ܕ��Mz_��5L����?9����*O
ʧ�?y" �Q���J�9��,���Q��?��'��I7+���'&�KPKC!|���+�z� �����?���tEl4��?	g[?��I��hϻu��`ʆ�
"
�n</<�����a�syR�'�2���'��T���ѱ(G<@ka�S0\��*A�'���p�'��aӘ�$�O����O�=�'�^Ĉ�o�K�h`�O69.�������O��'��|R���X��=�B�>J�Ir�̆1@llP/OJ���O����O@���<�Oᲄ��O�\*)�d��6`&,1a^��SS,��|��,��<!�+y����㕅	��=���$�"��i�"�'T��'��O���<��#,CP���H�)M�R�����ʟt�Ij�	��<���z���	ޟ<�I�&x1ɲ����B��4�K
6�X	�Iӟ�I"��S���|�ĕA���rF�>Hb���J^�'��D��yb�'@"�'��S�$b��͟9mI<��!���,Rx�$}bY�t��vyr�'���'�&S-�;<`���O��I�ǂA��y2��>6���'��'=��Z>{�'%Q`ߤ{ !YQj�:@��z���D�O&˓�?Q���?�GB�<� EU�*H*0S҈��'���pd���h����?1��?������c�4�'VJ`$d���Q�S⃧y}&���'#b[���I����ɚ�p�	]yrbĽ#�H��Z��1 C��''"O#�y��'ON�'�?i��?�e�ݞ-�X2f�0sBT�)D�����O��d�O|�+@0O�ʧ�?A�O�������lh�Sw�͢Y�bX��qΥ͓�?���i&��' 2�'���ql�b�h�wtА�����D�~Ɂ���?y�k:H$�'���n��n�-Ͳz��*ո����/����'��kӎ���O�d�O�q�'�� /��c㉅>3����3��&zRĭ���E�"<�/�� b�0O������(z��ټt%a�+Q\�LTlZߟ����7��Ĺ<A���yb�V/n�K%O�2Y%�IZ	��?!���?���t$�̓)АḨ�?i��?i��X�%��(��8�R��&�?Q���?1�P�h�'�R_�lϻcdn�  ''wо]sS�,]����'�����'O�t���'r�'���y�#�Bݘ���z<��P���R�>�)OF�Ħ<���?��p?h�Q�B�	�>�Ҡ�@�zk����/X�<Q�ܒ�?a��?����(����3� z�m��ihh��\^S����'�� �'�2�'�NC2�yr-�Y��)�J�b�|X�Ă]�Dtma��'�B�'��O�Ӆ��I�O6��V��w8< �D�?$&�)B��O����<���?��*(����?�'�&0���]?zUxM� �ͭ��e���?��s�&!��?��V?��	Ɵ�ɱTc5{f���:)$���N�+����'"�'he7�y"P>�	�|R��O
�4)�M��V|K�o�ş\;�|���	�M��?!���?��T�\���1\�L�8I�����Lٟ��I��+��-?�)O��'M즠�!a��#b�����ܒt��T3�䓇�?���g��F�'���'rC�>1-O�,�#�8A~Y#��נ6����-�O�!1����'��> ���ڟ`��c0�Y!ID�II�1���ޞ�M����?a��?�]��'�9O�mz�&.�ؔ�C��W���oY�P�'�lp*�'�I�O ��'A�F��<�`c�`A>	�8�I3�>1>��'or�>�)O���<��w���vh�ˠ1�EEUΐ��,OD 6O�ĸ���O��D�OX�����DX�L�4�& �^.e�f`��C2�D�S}�Y���Ijy��'���'|��piJ�,��t���<�^� �Ʈ�yB��8�yr�'02�'��O�j�i	�D6�0vŚ�z�ڴ��醹C�T�X�	by��'Vr�'E���'~��Vʘ u^"�.�;=܊ H��?���?!����.����O���
>�$Kr^4i�)3a	-���'4�iyo���x�������*R.B��=�ţ�07E�x��O\���O��;O��$�n���'���'��ӳL6s�Dd�6q�{'[���Iџ��MÎ���$v>��VBŮx|�) � ��:��w��O�q�>O|�DI���	�����ן�r�O���-@n��;E셲���+T��O ���O� B=Ox��<a)��!� �8�F�D'O�`G$kC����$�O�ynZğ��	����������<��i�[h (��a�&�qbӱ�?���P~S�ԖO$�9�O5b�(}B�SĤ� �6P�!���6��O����OD�d�C}�T��	�<I���zN�3�+�E`@)0'��}yr^�`�T	r��P k>�	��I�z�(���PO��)[f	Ӷ���	蟔������<!����q���7*�?Ґ'�B�-��i�Dů<�tC�<qP���<A���?i���I�9~��*1�X�Dt
S��'r�>�(O����<���?��,n`032@��t��P
]�,֬�v%�<�0F�<���?A���T����A^�Qcƶd-P6&ݛ�?Y,O��$�<Q���?��Ј�Dm�U���D�3�$<.�9 )���?���?�����)�\9�O��-:�Ĉa�@�Q+*ܫ�+J2�r�'���<��ퟜ��Dy���O��4��+W9SLx�z��a��c��'��'!֐�'$BE�~J���?!�V�:�j0��%}Ū���H,_n��K(O����O~��q��|���T�n�$ LF�nl; H��?���<1��zC���'*"�'F� �>���(	T��.].�{����?����?�#dB�<�-��$�|"bK�	
�Th�V-~�5K� 
*_�<���?q��i���'�B�'�2���,��{f�W0)�i$j	!pm(�d�)8�$�O����O��'��tͧ�?�G�[i܊�@&ǡ)�j:�)�4���' "�'G��>A(OL�dp��h1��G�Ƭ�u�G�yL�S��O�$�<Y� ��<�W��|���?)���F�rb흇q�~����ì��� ���?�g�O���;��I�pɾ!A2�8G�-k�J��N��ʓm��M�s�����?y���?�ȟ�Ę*?NQ@S���H���'��O4���OP�O6���O���d��o�RY�F�U���e�v+(��J*�$�O@��OV�������4���dw���P� by���?]E	O>Y��?�,�<Q�� �A�B���JJvZ�]*c��w��͓�?���?yO~"�U?����4tV,�T��k�Je��ʈ�<^����ʟ$����ʟ$�aD���'�h+E���ܽ�d���x��[��?���6itD��?irP?��I����I-~v�	�E�K*`

E�E9O~x�&�@�	��dȂ�����&��Χ@~N�+cG�E�t6c: ���	-ψ�	����۴�?���?���(t�	�1�2(�5)�QDK���=Y"��O��S�+-L��2�d�|r����P��
ϖ�:��
(����?�żi�R�'���'N�O"��M5w�h�#$�J�
�ƽ�i��~j\��˴]p�ԔO��:�'([-ynv��BB�7ܾD���S�/�7M�OJ��O���w�I������<A�ղV�Ր�M���P�����$'� k6+��А�Jc�,���� ���+!X�'C
8��`���/2���	�$�I���'(B�|��Z�ĥ�v�K�&��E�W�qt�ɞ-�j��I�9�4�	�����L�OiZYk��D�v�̓$b�>�jp���ʉ'b�'$�'r�'-<�葃��ᒧ�0d��\����$8B�A��y��' "�'�O���N�-Nv@9�(ُP'� ��o�x��'F��|��'Gbm��x����	ܴ!!̐�.���a�����`�'���'��䤿~���n���8WKn&B�(� /\C�l��?i.Or�d�O�dX	41H�g?��I�q:�BqA]�n�b�T	��X�	�!�y���I��I�O��$�O� ��
�&L-S��%l���$1��|2�'�R(�7�yR�|�:�N�5���y�0�FaP+%�Ι��'��c�'!"�|�x���O�$�O���'��!���DӠ���{����(O~ʓ�?Y��O�~4�'�U�V��Eke V'6IX��`/�_\r�'�f7��O����O���	l�i>٪#Oש7��Y#HQ�x��a�{y��'Z�O�I�4|����O$�����".�`1�l̲K ��Æc�O*�D�<����?�����O��I*
&��  o9ح�'�$a�Z�[U��?�����H���<��$>�RCLO&�+a_��'�'�R�'��O�˧�?�(O�I��̍<���(�@�^�&��<�@�<a����<1��?���2�O��1��^����ՆQ�Q@c��?I���?	���?!I>��yR���@%�A2�ۑ@�P�kr�I#�?���l�N�Γ�?���?9I~Rf�OWF8�%��-��9�ӤA��0(O����O&�O����O�H�g�OVQK-*��l���ؓl~v3Āʺ�yR�'<�'��O���?��.�
Z�J�����
z��ĺt�D��?������?���$�=�A&Z!� �3��
$=��k�C������X�%p�,�I�����O��d�O*����K��%� ,^f�
7��O�������yT�iH�B�\�|i���`����B9���O>m��T��ܟ��ɹ��dG���X)1�L�Ph��C(C:���'���[�O�ʧ�\�ۤ�!zW��H!_4�ν:���?������'f"�'��"�I�CZ�(�F�!x�N�! ��~	�	�Lm�#<I,��q��1O�$V<K�^Y��Ȏ#\�B��M�Y�F�oZ���	ȟH�ɶ��'3�<O��V/�K|Z0��k�5��Ojh��'z�'<2�'�BHK�`��ă�GҎE���Yq��c���'�>��ߟ|%�$��S��$5��"ȏs�|%�0�jyb���ybo��y�'~��'���c�|����Ɋ�k���UK���q�	埔��u�I埐�	\��Be�+HǪ!�A��-̺� ~�Ly�Ce���	��d�I�?%�O��i�6,��zQP�pڽ2 ���^�D��P�	��@�'[��8Ŏ�*2;��;�Țb.,�TcC/
dvQٜ'�R�'���d��~��5 �f����pq%�>��L`���?����<��kDK��'�!s`l�:<x�@�ȉi� ���?���vbE����?a(�Lʓ�?�FT�7��`)D�oe���K����?�/O Ƀ��ɛ}�^|�n��0i��Ĥ�9%T���	�_�}�����I蟬�'�B�'��i�3}ڔ�2@�(��t�0ZM���'�	���"<ͧ*��a���?(��c�Z�� �u+��?��#r���'��'=�+.�d�O�!�Q&`]��;�ML�u�����3|O:���7OF��U&}6�Ͳ�H�g��IƏ�5��hnZ�l�	ٟ0�I��ē�?i��y2j�9W��ɠ�`B6�����f��'r�A�'Q؀h�'�'7�*�|���� �%)>XP�p"�'n�#���O�D8�Ē�ws2q ���*L�Lr%�k�x˓t!��W�Rt��?����?������/U�,��<bt.��� ��"&��?Y*Oj���O�d+���O�	:@��E`�O>l�pc��w��^�#�->O���Oh�D/�)��?��Ҧ��
HЈb�GfH�kB�<	��?�����<���Y�7�	�,�����G�,\ƹЇ�O� |d�Iџ�I۟��SX��]>���R\�PC'@;þ�b�!͆N���Iퟠ%���	myrd�9��IP|�(㕢�)�e��ȟ�/J>�d�Ob����Dp���O.%�O<��'���O�%�����Ś7���L�q��'��'���ӈ�z>)름;Jd"��t�^kj�9s�I�O�MX�9On��J������@�����r.O@�U�Z�l�܁�C�C#X|�����'��'�ޔp���|��Ki�����:
R�&��3�j����?1��i�r�'���'>O��$�\4>MsRui�0�c׷v����C&Sr��S�r��?���"`�L+Ю%�����ʺ��&�'��'72�?��՟�ϓ=�����y����"��8��?����<�ϑ�<����?A��\��3��*=I���GA3j�������?���W��uy��'����seh�2�n�*�kG6k($�a1kyR��yZ��;�'b��'��?a�fӒy|�7��NܨH-�O� �'��	���'���'��cD0/��*d.CM���\g�jQ�� j�x0g�l�P����	x��zhS"Vl��3/Q;Q>������'�RU���ϟ4��&%���I	ZtU2���(�l"ӭ$܀h[���O����O������'C��S��đR��S%E�xY�}���џ��	{y��'Fr�'1����O��I8A��	pC ���<Z�
O�1����O���ZR��O\�Oh��']b��bK�=�EB��*9�8BW�F�	��Iɟ��	埰�&}��$�ϧ��a�Q��C��Q��(�C. u��	cʦ�I˟*�4�?q���?i�?���	!��(��i�^���K��
�����ҟ�	��IY�I�ĩW YK@�>wlD���+�&L�#*�'v�<��1&��5��1QB��17�����N���ϺqV��Ґ-��� 0�)��71؀]�����q5�'?b�i��7�@��4�I͟\��v�R�0"A��nMe;�H�2r���V���Q4�"��Ƥ@�X�!�bW(�P�*4��@ǋ:� %R��9L��3��7~#r�� �P9C�Ab��"M���Bt��48��œT�#xlxrt	�!R{#��[3@S*$h6kݡ�p+׎ެ�ģtDS��#�/O�&i�g�.���e�:(��@���;4D�&A
���{��H)�hr��S*OX�����-�v��S��;=��G�4#�8I:2�E6A2��X<c ұ���
h��F)f�B�[�h\-h���NB�6u�ҀJ&�F�4e���1Nr�����O
��n�"��Q��HwX;��(j����'� �����{W��J�U��j�O�1��	�sc�����m��8��k}40s�`�kV�ص�>iQ�>w�[�i�\�Yw��6 ��z��Zp0��'�	4��SL�T�
���C
����J�"	���n���f���=ҥ2�"�	!�HO��Y�Tl֪qP�c�N��0t�%Y�����?ٶ�57h��'["�'��	؟,���1��l� r�~U����#p] ���i�N}Y�h�'=��mq�'LO8QT���r��ACI�T8��i���"�^&a\(@��&LO�\�LB:>a�y0OۖtV�{@�i�Ip���?y��$-�����R��>�L���>k�!�� �(��Ւ�����`�h�Q�lq�O&��&A���O�!��o81)� �b�� {B̀џ��	Wy�'V�=���!LU3?�R�s2��
N���0���;7O�<:�b���3<OrU���Z'*��5�Q�_�~���9`$6O.U���60��d��#<O Y���'�"�i� |+`MW��(��
d,�$���D*,O`���ס�L��G+��!;3"O�a�w����4(vd؄-ĔA���މ����<�S㋿���͟�$>��3�;����UBǙR�L���a�+�?1���?��(��rJ8"P�B��R�S�����8
Rb4a�V)��j�<�9���=5�\��D+�XUG�dmP .bH��N���v��cm� ��'r�X����?�����ear�iD�G4&@(��#���ēw���+F��\t, s��>x/fU���"��'t�Lj'h[���y�K��n�l2�{��'.����	C,�H8�"��m�
l��'�!�C�>({*���B�>^�v;�`�<�~��BGC�X#JЛ���3$џ���:�����٦7�l�A#$D�,2��ȯҭ���*��`g0D�`Q�kЧk�XG<'��X��n.D���V�ۀU�ZI��/:����&3D��Co�;n�`�A��|��L��C5D�|Ij�2E���Sp L�Y�vP���4D�@�BP5�nLQ C�;�R����!D� :�a�	?(։� Z~�Z�b�:D��!��C�HvE`k[�\0�J�+"D���3�-	�eX�i7{i��) D�2Q�M�7pJ�:���+�uS�2D�0��E�9~�#�bO�YX��+2D��DNC��}!O�=B*�(�	"D��Ԍ�7cc.8�Q��'���e�"D����/H(H�(#$�� z����� D��p���S۬�jGB�u�ddڅ#D�d�c�)��VLh��K>D�<*B��63����K$%�.��ի?D��)s+�0�Ĝ����$<��U�<D���ێ}��ɴj�,h�P�p�=D���38�<X�V��<�f=p�'D�\�e�t�6
cOB�vf��"0D��0�X�{������ 9vha�L0D�	��I7VL���Bއ@Z!�M D�P�	�7|��DS��\�bv<U�e D�8K�-u�4���]7	}�t�%D�l��	c��@� S�Hys'5D����dD�:)�8�ժ�(s�РS�*&D��I�l�G�0}�㈺1��1��%D��^$"x"i"���Z�v�{rL?D��a�kڤh��A���=�<  f�9D��7�/O�L��b�Q!}d4H��7D� 8��kȥ@�Â�U�<�q�.D�� ���0*";�~��@��JY��*@"O~Yk�ʒ�*�~%��ŏi5"�(�"O�	G��e.��VM�+=X0"O$��CW�r��b��!Q�pR"O*�Z2,5s�T�9��}��"O�l�6��W|�����&�b"OT�k ��Y�4	cb'X�Cɀ�9�"O䙊E���)p�� ��!�f�'��a�r@�X�S�O��PS�+Ү%��Y�E�R����1"O��۶�Q aÄl�6��@�l�U�f�[53,� ��I�D�N��`n\ l����#\�]h��hAA�F�L�ˠ�u�<Y�KO
<Xlx��,4D��8P�j��)C%M�#.�AD2ʓ@(�h��i��#|�1I!}����̖/f*�҇�Cb�<�ѩ�7%k\�Y����F�4���$�
�parFԞ���O?�$�2�Y��!�0��J"�Ďr !�D	�+��Ɉ�ă8$��m�Ԯ(�'�e���0=a ���v���T�U)��X�Λy8���C#H8i���Gm<��d��,���\a2��7s�!�dۤ,]���d}:�І�K� �Q�l �-�'+Q��0��Fj�  +U���a���{tC�ɾ��@�#��{�(������5�쫁J�68>Fi�7�"}���'1�H!���Z&��`��2?����T|.���SH��C�c�?S�����4����&������ �z��׭�8��@L.�|2�^2rf�P�`�sX��d*�Y.�U��E�;6FnL�=���"5$���A�+:\���aF=�n�
��N���x8� ��*���}jpnʏ$��鳄�i��l�gd�964�c����?��L4=��p��4u�d��%���@�Ï��?�O�٢�A�j���'�ʱSǥ@�������٥g7�"On����+m���bH�m.2q![��ه���$W���t�>E�4�ךq�va:P�̓j$p*PȌ��y���Bl�7�@(d*��
Y4��'*Z�z�`���ϸ'\T���*Q�H��S��r������YZ����S�Z���_2/L3�F�5	��%�O�D1�-F�v�d���f��Y���{���6NΡ���Ok�O�2!c�mF���a��591L��'���P�DL�:Rީ0����ؘ8+O�\AB�� 8�sK��|b��*º��klU�0V�<�wO
�gF�q��g X��И}��8�P&���Mk�쀉�*("K~�=
��u��P�`�@�{��V��`1w
�5m���A�R�L!Af�?#t	sƈf~��ie�a{��[�<���!�->mi����y�ˎ#���<��+��!��*q���%��e���<��9;&��*:�8��͆:n%* ��'ϐ��B@ĥL����K�g�r�k(O0�3f�i\�0��#^�b�J@`�&t�d�!�e�s�4/	�2���I�2,3��Q�-�/�>���+\������ܨ!;�Bű)F�0��,#*�`a� Z��4���E�E�g�I%1Ί�p��.$<�c�`H+z�Z"=��b�bO�%��+7��l�DBC�`I �6{Tt�)D�~���G�nDt�g�')�-D�S�1H�,"�P-X�%24�R�-`Ԝ>%>5���6RH&���h��Z��xs��w+u衬Ϸi�B�Iy��r�!�<!�Uxp�?����!�V(C(������	FV��H�ؕO�"�ypl��fd����-,�:��]V]Z���&>

fW?4XY����Kl꤅A!bgx9�##���IC��yBKϖ&��q�fʋ*{Q���Q�P0�HO�i�%'ʑY�4U#����\��<�A�UN� x A�9�~���(��`R�'���b�Ia��T�I&ʰ޴5�R�yFɌ~�ӧ�O<�8�&�ğ�&�)J5���gNІn�����2D�(kj��v�(h��`��x9�y2��<��i�o����p���JҋȄ!�I��nG�y�������Q�~��W�V�i����6�  x$���5"C�Ɍa&]y���C��4s�ӹ�\B�I��1�0�Z�.��'��xC�I�<v2$"�`P�.�6�6��C�Vc�����B�剂@���@��� ~4I0��6j��(2�Q>�4z�"O���$Dn�l��U�^�πN��\�p]&��
X���OZ�'(�M�d�8.��'�	*?d��
ۓ5��, aŧ�H�4◝Sih��թ�]����n��m#v��F�_��(]J�D�f"W\�' 1��L�=i8��#g�>pqΰʍ{�9:bR��8O��yC��<c�������a �қc���6f�X<`��+�4��q�?�O08���A	RV�:T��*�aNò�p�@p��O
�Y��M<�0 ��� Fqq�kћua���A�C�KT��="�-�dEV�:o��ϔj�<1p�Уe��0@�D��IP;Y	��[/�
�+������#0eС�?1pO�� �q����1��5�q�&�ڟ9.���c�(LO<h+�m�vZѡ��t�`���!��}k�Lp���/f�����:�Q����O�����L�;Gn���D�2,�zp��N������� q61O���B�� w<8���8���ʛ;)
��	�3/�V��EōH��bqi�����#ԛ_<\̘������ o���p<A"�%34*]ْ�X��#��W	"��y
��O�ء���� �x�H��36 E���Z��3�m׊&��E��#�T_nA�߃.Zd �#�[�J<�������@�0O�a�N�,\���C(�R�� DD��䒅(�>�((�P*E�yZ���cb݅Z��i߈(2m�V�6�]G�h��ؑ�O "��*.T�D�;�$9��1���b���+'DP� fd��I^=@�A!na!�у
rD�w��_?B�$�8������ўj��|{�)�A[W�S3��Fn�z���I�ta05e���?yk�'_�	�E�'�y�l�	Mġ�F�2wD��۳�剘k��AЅ̈́j��g�'�b�R��]�x
F-����i,5�Q�U`̤@c�͂1�?�BA�'�X:Dݑ;��$_�N��bgŕ�� #2$!- @ � �R)q\T��ɜ@]� �A�$6P���1��|�IQ<.�i���ЅL���1	��;�7��7�1�IҖ0m:U���S }\�H^̜1Ԇ�7-d��#�J����ǌd��r����(�l=^6m�nj$p3���SM�N�]�$ʕ�PAN����Ж�|A�A䙕M�NIH����	�
˓fR:�j�aP̧} {!?,���$蝹 �P�GӲ.���R�i��s7C��	�H:��D0zT�-���:q=F�Y�o�A� ��'�2�� DD�L�D�Fty�Cz8TՆP0���I16�٣
��8�&��A�S{$�`�<�t���.8.�q�g�4 �	�3J�=�*вYwT�Qش��\�c}F��H�s�#01�2ϓ�K�Ó�3�7�[�6�8i0 %�:��pջjR�h��҄^�K���BiD�����5�$]@��N{�5ꦜ�"/��P:މ�b�
6sHh�P�I-"`X����;ǅ_j�����2X�-�����Q���C���24-3�$�
!j�_k4��!I+LO���C����)a�ý&4��BRO�;�8\) 8O:�[��)!���[wW�CF�����G�ɼ>����/G�<.Xr��I"ah���!�^z�<q'�� *�.��F�55|X6��tU��Ȓ�8oL�!c�`�re#��!)�(�+��œ%=�N��m�+���r֋�p��R�"O�X���Ѿ���C J�'�K�)NU6}���V��1%���h�½���ҴN��� .~��&�l�E
&bX�1�	\UH �r�0lOd5��늉�?��[K�"�@S�]�t4�|�)_<_�J��n�2X��(��ϕ3�����0"�=����j���0�Թ1�����/5@���m݅V�ҽ�e�͙�����#����T+�x���UM_h<!�N;NI�@�GE�/?��pE�r~]y��I�@chv�)��	�)��q� ׄ6���K�+�=	*��A"O4�;D#�;,�èӿ\�M� .��E8D�01:�:��u ݖ�1�8�O�9���':rԐ�W�9m��r�O�!�mݖm!"��5c<��9²N���q��bӯ[8�t���ܢ-���_L`
q�B9qzLY�P�Yc�xrHĸ�VY��k��V�~N8���]�����Қ���c�ÆT�<�TFL�j����fTobI#D��M()�ܪ�F2�Đ!�<����a� �c�����k���a�"O�T��' v�!V#��亥�CϏ$8~�i) �2�?�p.[�:򱟉'Ř�`���4a�
�� �]Q� ͉	�'0�E��j�$!���j�!BM�N%D��L�X:��-$(��'�u�A�^��5�oė+z}{0&<O�m��Ė)rmc H��MSr�U�2��A�F�?#��Ybng�<Q%�1[��t 9<��&��h��|��	T*(R�#~j�O08��bVŤ�� *�b�<���jmd�"ׇS/fw�#�`�	������-�g?q��
"K.v�!�		2u�ms�OZR�<�e��1�@� �L�!��,����{�<����)'��3��R%8)�c�X�<1t��/&)f�A*,�v	[ �D~�<��^�Se$�[�L�/E�W��s�!�D�&�R�9q�w0<�HW���!�� �-3Ԡ�d��}C�mW8&�D��"O�9��2pƽ�S�T���9�"OέxN ���;q(мN�:��d"O8=RUmց$�<����`��G"O��(R�P�
��Q&Ls�Mj�"O�#4γ\�`5	s`�2Rk�%I�"OX ��b�"q}"��.�U@��F"O̔!��IZn sB��=ŠA"O���%ǆ��b"؜\�4�"O�U��*�4kD4p���>N�Z�"O6� �F�l�0i�a]<`8S&"OҴJ�"W�c3xͲ�i�$C�"O2�3����tP�-C��%�:�"Ob�I5FM;Kz �'nԶ�J�"OlI���[��B�Sq�T3�"O�2R��J6HH�$�
0>�vi��"O�� D�dM2J�'��;�^�#"O�y�'�,f�&]�"KX�N�8�"O�d�to��z� �����b�"p��"O���EX�C�V���숁7�H��"O&a���ް٪��C�bl�P�"OlH4h]���h��K��4�}�#"Or�U��4E1(�9c
"C&���$"O�m��MW� _��ɱϕ�}� ���"Oxe�ׇӆpC�ҔX��<@"O�����¦gb�`�cA\6T�V"O��[��<
�0�d�TX܀"O��r搈w���� U��b�"O�5{�(Q�4�V������)��"O�x�v+X�$Z���;y���sD"O0�����^���	d�5͸@�F"O�6f(kMN�۴����M��"Ol�!�&UE\� ��A���D)q"O��b��.6��P�����ڭ��"O�[dL�#;�r8˥EI;vxP�hgO9B�z���F0[U��w��q��?�#Cy�͘��"�&���f�{�<	b�ݼd2�<q��	�D�ty�<��+�<_v����
�9�����Ls�<	��Rz;� ��)]�@y�W�Wu�<	�KC��*��C�E��-��m�h�<D�U����R���P~��Ӡ�f�<�VK�/[րB��3- a�.�{�<�σ�nH*��4��-p0����@x�<��,�U��1�GS�]�H��J=D�<�Ƀ�	��,���RU]Pr�.D��do:e�ډ#ю�$�&hإ�,D��R7].�; &� (B���֣)D��0CV�����sM�2YZ�#1�2D�(:q�1<�.E#w���PL"t+0D���c�9X�l<�S��h�j��Ƣ)D��)�憲+R	�t��XJ�&D� b*��m`D��H�"�B\.�TB��?st����gF���AqŢN��C��9��ua D�dڹHƉ�! 5�B�/�0�S���}���v�B�I���Ց�o1]A
y`�'��B�ɘ�"my�fʪZP�$��G�"��B�I�< J�pt)�yv���Q�h��B�	�-���v�^:j:�a��(ϞE�B��M���+
�b/��*V
� �`B�I�D�Ơ3_	|�`���j�8�B䉲>ܶ��b㔦B�8U��@�n�C�� +=���o�F���i܏fi�C䉯	��c4興39�v*ͻbB�)� �1� �"��(�u@�qL��`"O��rUE��9j�ioO� �N]3"O�d�r�B�(r8��ĸ .�3A"OX�x��E�8���WLB5i��,�"O Ӂ^�ZI̛�F���"O�lӴ�X�@Id�j�*�2k&�Eؖ"O���ʨ�GIp|��`�"OnX�n�RG�=�`�]qe@ċf"O2U���R�}�D8*ii]0��"O�H�f��r�0�0bX�x��'�Zp(v��6���rm��9�$���'�ta�䎦O~�p���5'�����'���#��P^��:0���(�D�
�'���QS�
���BA00�TT�
�'ߢ��t��:f�@�,���S
�'�肱�i�h�W}��'�Ya��=d�½�FF��,tA�'�t� ͷ_�*�bv)-�8T	�'z�x�.I���KC�I���ҫO�h҇f�r�S�OjƼ��C�Z"ʥc��#='�%Y�'��〆I`�l2q�'*��%�I<q��J\az��6|e��Ӵ��?7l(T���ҁ��?y� h�8���C�'-����ǳ3p�;$"O0��R��sĩj�Օ^�y���ɔf�V�؋�G��JT��LR�H<��ѳ���N!�SLʬX�(�"F��@⯍65�ɀA�
�}���4x ����	4g���ɱ`��@!�d-C*)��ٮE2j`"�@���'�t��d LO�Uن���-� �B�M��'�2��2�F�)���3����� =SLB�=je��
�i |^�鉔��$C#?is�VI�>�Ґ�P�$I����O4ҭ;A�0D�\�dLQB�@���'Y>s���)g�>��;��O�>��HۃPpdA�I$B�6Ɉ�?D��w(Q!c�`hc� (�2� �=��,X�E���'Z�e���a�ԙ�������ֵF�S�
�x�6�q�
��!zGl	w�'��Ón^�5�Ӊ%��!gBCf�f�F~�.�u�^���c�>e["�сsά�%�)}Ȭpp��R��Պ�cF�qz�  N�&�'�9�F�(�	y�'�x�2����=�A�4N�y����'Y��H�OD!2^>�Z��8p,<E��y2�:t$�O1�hh��	ik�%�vq!�"O���!�C,izL�9����t���0U ;��=�"|�'I����F��$Z|Z���'�.���Ļ^Q.�҃�ɫ]�����ӳMG��p �9�%���ll�IQ���?�p=af+Y�I$<(� ���0��5�d�R�zB�	�/�@��B�A�r����=��B�I�e9�a�?�8�c��:w�B�I��:�Ӈ�1��M�ݩ9�PB�	i�D���"N�O&�c6)�- &"<����蟔I:�dR0r�<pM�)Q��"O�ՠc�P�?)ZA"���&�nZ��\>��"~�~�� R���तۄ�W�~}�ȓ��� Y5���ƭ�&DZ���i���%{��I#1A��}��C���.܅�	��L��' �	C�D#s`�\��n���'UXTJ��H�E�v�$�-��-z��T�AǺ���,�TC4�X�cU�iBf�� (�y�<9�dV"t�beH8���c�`~�<ч�@s�iyBY?=�[�&�}�<ag�� $o�tS�n'e�i[ZH\��3~��+kG�-�����1�6d��S�? �9ӥ]�L,9VkR>_[���"Oz� )x�B���#Z�p�Z"O&q8���;c�L:��X$D�Ti*�"O �!!���fe�����&6V�v"O�U�KO E�ӏl����"Oj���MU�D&�cS�5*+�4�E"Oܐ��^�d��XFK�2����D"O��Iq�	�l�
��!#�5���b"O���Щ�e������w�Rx�t"O�p�G� ��C ��wzΩ�%"OrHԬӜ,�T]�eMF�Vy���c"O���t��< �j��R�uj�<�"OX��W��>,6a�iK>e�x�"O���Y Z�V�`VK�_
8�"O �A�b2���\`[L,�U"O���@��)��3 � �E�&"O��ҷ�O7␠�o\G��Z6"OR=��B��F,�DO\5�"Ov	����%ONf�����Z�4z�"Oeᄆ)0��Z�o��^��Ix�"O����$ͯ�H��.W<]7ެ�u"Or�Yv)&VX�ȁ�G�?<~��"O~����7Tj�(���\Wp	 "O
� 6�X7b2P� ����`� "OZY��<�R����m�TV��@f���l���fh2�N����̏�e귯U7��{��Xa�܄�ɲw���R�wOv�h�����<��6�H�vGf"?���6H]�N>9ƣE����Cb)�U���rPǉm�'F|=�Q"A y����DÀ	�l#� � ۸`�kU4H��� Pj�L��m�)§|P�	���s��Yz�.��p⼭m&預��n8O'���|b����?��#�z}¨�j���BPԸ���0��'XĘ������Ϙ'ήxKƑ�fZ�9˃�*m0̠�O��R�H<pF�(�a'_�I1cq@@�	ĺ3��Z )��i�RC-C<ز��C`mѢ��$�p=�đ\S�N>4*��%`��$�����h#T��ǯ<��J�ia`���45(�;X
v9	b�˭���l�,�o�70�3�Ω!�R��d�E��5,J��x�ȗ>D����¥ׁQ�޵��ꑻG�� ��I��<[��L�[/�v�8�96&����:w���32�=Tc����#���џx���� 4Ќr`oR�<�)!��i���H	>4�c��
(������.
�M�-�B��8(Y!��Y�b�,d�'@�i�b���
��M�%*���&
���$X���s� ��@q�^� �6y�-�>c���D?k+�Yr�9'i�-��#���.R�E�ڑp��ў�"�9�0��4�;c�컅!�<Q2C[`�)���`�B��z؟�Z�h�(jˊԓ�"(A�=�0�ǁ`4s��P9�Ҁ���hK�=Vg�	�gن�;N�8��ɋ�Z�p�����V�٫�f7�ޔ�9��5e�fq���FU{��o,p���%$��O0�Ȑ���>�d� ���M���A���jb��$)*	Iy�±>�CE)��HK4�ӀvNX�Qr�\oqTD�
%�i� z�2H�H�����fٖ5v!�$_!l�5aK�r8jWd� OrT��:1�6�#C��V&�B��TK�2'-
M�'���@SȎ�\:���$F�;� ��L20�Cen�L�Ӊ�50�x-�]�|01S`�����+|��Q��g�����	�h�495!��or����1�f�"����dӔ|蔧E<5O��Aǈ,6������L�x��(r�1���`G�/�Ovl�D��
c�"M�A�@�Ի7��D��Ec�Ӻo:��8Ey�M�3&�&m(�gB)o\PC���\Pr��5a��r��M�zo:c��pĬ=LON�r��MN�m�g�:��DuO\$�G�i�Ub6B������w�<�T�X3Y���`Q�ҙ(:�yB��nX��Gy�hN71�����'�,f��'���y�ش "t��@zb��!�U��yₔ
:�"1��i�Pr���y� �-<(.�cu��(+��qc�'��yb��d8��!2N[!*YFD����yBM�$:�BviȂ!����$L��y
� H�BO���<�j�cTf�ބ	�"O�T�� b[6 �"`��%��9+�"Ob���M���A�ϙ�m��53G"O�Qp�	V3��x� ^B l�W"Or�����;֔�X�Ă��"OB�:��/GV������4����"O��z���O��%	�@<�I�"O�ݑwG�g��\��C+1�pK�"O��y'�˭1'�u`"#�#���"O��i�o�++���W�)撼"O�1��(1���a�&R�}a�"O8`�uƢ5І`;r�t(�B"O��K��9H�٥��Q/��"O�y�� K,^,IBoI�\��2"O�r֭ H��3qny�c�"OIp�Ԙ+@���m�(Pl��P"O��8�5j�%R��%i��z$"ON�33%�5@�|��`�vW<�"�"O�����Y�/&1j�/ C�5b�"OQ�4��x�����ݑ8��"O�0�[/��bUcËd3�,�"O ic˕�e�<h��ና?="Y�t"OX9Jt*�*����g`�� 1>�X"Or�xC��#L�-�$�7}Cm��"O:4��$HIB�ʒ�6�PH�"O�Dq��\�<ͦ�T��<ž=�"O}�F%�l���u�B
T�ݙ�"O�����Cx�,�j��_I 1�"O��6�I�6���1!����X�"Ov�H�F�$C��!٢ G�Q�8�bF"O<$�`�ړ��cgΫ���P5"O�l5�գ!E�(�d�ɓt*0تW"O��Q�[�~>��*�r%���`"O�(w�U+�t���I >�P�"Oj� ��p��z	I!K�d�d"Oh Z�K2j�Ab)�_�(�"O� �u��9@�0!�é��R�Y� "O�� �-J�7�ج� ��v�� e"O����݋'�����Z�Z5@���"Ory�b*�F}T�����%#t�Q"O�p��θ>\ԑ1��"�Ur$"OX�I(�6!Lzj$n�L�}�""O�D�v@�.t8J�H�L�)^��I�"O��
�A��.
D��!�9)���6"O b�š6�T�;��C7���"O(�����'^����_4�zr"O9(��K_.|q�$A4=��yR�'�@Q� Yp2�
�C ����'��X��S1=D ҪR�Es���'�f�"AkZ��Q)ao��&q����'Eb%�B��8D��[��/���#
�'���K�O�NH8gI�;R�rX��'x�,xŇ�v	@9[qG�L� �Y�'��
�c=>A��w�ܧ^�*�'r�q{@�Q�'�ԅR�SN����'�#��B�=�j��&��]�ze��'���@�F'7Ր\@����PWN,��'�������~���+6FvvL"�'����%`�x8V�bp�S�8n�Aa
�'Tp�)�-x�h�m�=��К�'�:l1V{UĔ薅Ҍ9K�@��'|fE�V(�lz�I��LϚ63T�a�'�̕Q�N�H ��u�I;z~��	�'�|�PRI�17�Z��ơ�"JЄ���� ��Q$	%(��-bU��2V�!�"O����٬"���3�H3o�Z�q"O��aUs~���+Q�.�D5J2"Oj� gˊ3b1`�� +W?��x	C"OV�!�'�3Q��� ��Fanb�!��ZSDհ�BT( �^Pa�n�0> !�
{�-�Qg=[���Z����?!�$#<�Ԩ(<OT5Yb�<z�!���8TM��4�3<h�Q!�^�\_!�D�?�u� R���!���xB!�Y8`xn!Rb��7�bX�ʖ=�!�D�(̴J# K9G�������V|!�$��=ؤ1cG��"�4J�G�!J!�d��������I�Z�J�.	�,/!��.V���D�E8\i�@���Y�!�*"����!� !&��E��0#�!�M����T�W/��<�t�K�+)!��"t���ʒ���i�Q�ڄ!�������O(:ij��dD��!�dφ(�.�zn�=j�D�SJ��!���V����P���gRu�P��-�!��ՙ�%�����@O�98�{�'��I�&�4l*�dM��L�
�'�>y[s@�
 �N�"`�S5ZK(�B	�'���+O7I���g�J$gh��
�' z걏Ǽ�����^M��9
�'Ll�"��8�<�B%!S�b���	�'��t�R��<:Ոű&#[�dU	�'���K�/-I��q	Q�W����'Mv ǫ
#D��ɆRǰ9�
�'JJ�y�M3�8c��J�|�VX�
�'$|�J�+��U�D��$ҷ GBT�'B0���;�������~�0m��'@�*�ͅR��샕A�6yX��'s��1g-�6�,�B�m�.�I�'���8F瀽i�@ܓ�Y�icn�A�'`�%�Щ�3��Q!�D�0hp	�'1ĈU���)��I�b� ��Щ��'hDX�6�ʬ6ɼ墱�<
\�5�'��h�Vȕ&([� ���_��j`��'%&a{$hM*	i(	�֡����'J|��"aJ�W�^ x듉yMV�0
�'�`����U�oh*�b�c�:�T�y	�'
����j*�@8�4���-;���'�`�`�S�k<� �Ñ(��2�'��yA>��m������~t��'+V �䕊c�@q���Z"�z���'��P�1�PM �b�Ck���'2vh���A�Rvh�Hdc�5m� ��'�gm��pʆ�ۂ�^@����'���� ����ǥ��j"h�	�'�ؒ��H�Z�
�.�4.�A�'�P��BW�����T�I=�J�'s��ጞ�~U��X�E	 b�"UH�'�l��L�Hj�X���$0{
�'X� ��#4���P�e�|?���	�'�����h!VHj頕�Dy5��y�'u��t�fz��(�q�� �'�2��7���NG`���Є����'���*H��}�����.н{t����'��z ̓�!o�dIF�gu���'�)�6�ǀ]8<c�o��a�P���'���Cd�p�P�ɱ�Z0a�'��1aȊ�Bքhːf̒X������ h�C����q��[֠L!?�1�5"O�U	4BX�<xz�s��P�I+�T� "O|03�������(;\����d"O��'�RN�|��z�."Oz�p�Ad�x����ǌ��Y�@"OL�y��
/I�hB�(�LHH�"O���r	�9Z�P�4��K��S"O�X���=fXS���-	r�)2�"O��S�H�a~� ���$pb��x5"O�a��2U�<�8Q�\ -S���"O�1bۀ:u*x! �e��B"O$�1 �R�.I�sUK�6v�6"O�-��:nT*P� K�/����"O-id��=*�p�R��\v ܑ�"O.�iK�r=~M���p���C��yr�\�Y�f@p�ˈK2p��ѧ��y"@�n3��	g�/lR�3Х��yr���H1[5�XZ����L�y��Ώ:��=# !��I�8h������yBXGDD�����"�d���ס�y"�ŅI��hD�!I�B�$Ɵ��y��T0-C�J���D$�Y9�f��y2�W�x�"F
9}�-B�	3�y��Ԃ)t������^�0�sFb���y�(.{�2X�%ꈬ[��	�NU7�y2�X+P��la%I�Ur&�"p����y��2o��x����\7bE16nߺ�y�ƆL�Bf��� ���+��5�yc�<W���"��L��:U��y2��%�<�"�g�A	l`���>�y��
X3�AC���	4�h������yb�Ş<� �a�S�1帹4n]��y�E��Zs�<�R�׻/�B���%�y�`J�8$�k�R��l���yr뇷 )�ĉc&�u˺ �/��y�
P����J�7�4$�����y�#R�d���z獀�/��y���y�J�7��\�w�G�O�B�f�I��y�K��$^�*q��B�R�"���y�dƢf�FD
�+ذ9�4Up6!�$�Fo�ab3,+[������f0!�D����m� A*w�}�BH�5!�Ni.\Y�&�C-2�fQ.�!�d2V;�4pSc��j(��L�!�!�$��́B�o��¶��.�!����*�KM;az��z���'�!���!�����!�$^���WF��z�!�� �|�tCC�n���2S&�x�a}r�>������pk4*��|_Ba�6�l�<���=hg!��Έz��WB�<q�dAO�x���\����P�DB�<iK[�A�D@�C�=0�x!��r�<I��({Z$�� ��G��=A�ʇW�<�0��!Җ�t��L"��sa��U�<�U��u�|�x���0G"\�P@�G�<9q�A�B� Y��ۅ �9��GJ�<Y3��	 ��&@��4=�ա%H�<��a�}�֌J!�<N�����h�<����x�Ht ):���۵i��<!B�	q�Μ(�U5BC�J���`�<I���C���sB兰X����3�BQ�<1���)'C��A	�
��1X�Ie�<�^:cr�)uʁ"S�:Yk��d�<�ਁ7%:V�Z��Ͱ$��D
��/D�� ܭ@��G�srva��^�I_8��"O����(z��pb��+-v	:E"O��2Х7!@"X;"!�1o�jM@"O��'�O�2:���o�0N:��"O4��
�; R����nfM$�á"O�H"��$�1CX!,<�Ճ�"OHdYUi�-��*e��8!^��B"O��Zc�
U,� 'n�p��"O�t�ޑ�N�B�:�~-��"O.�1g­/P1���(B�X!��"Otl�kј"*���WT^�B�"O
�F�� ��%+�=�|�Q"O�8a���t��J�?]�[�"O�LXD����ZW�X��f0	�"O �9p)��U����)}�z*3"OH�B���·(�g���y��G.v��-l��80PdYf�W��yb�+5���(6���U���y�k���S�D	`0L�E���yҁH�����.@�܉��B�y��ŎETt���V�4���v�f�<��.�	���Z��Փd���&n�~�<	�4p����Ɋ6,D�R�e�e�<ْ��2u�j�PC
A�`�����^�<1���Qv��I���b�2A��MN�<$��%F)���ʅm�<d��DJ�<�үK�_z�s ��o�u
q�I�<i@�"uy����	<Z��� F�<!t	�A(� �X�|+�0���i�<�@�͞ f�	���=��LC��Wa�<���U^�|<�c�K$U
\��!T� � c=�b���C�~����!D��'��/[U�L��I�	}���@F?D������K��� &M)
���s�<D�
���545�뀈L-!�x��9D�P�d&Z�zj�=���%��T�G�6D�X�A�֡1N4��!��Fs�t#��7D��j���.?��b
�;��Ё��5D�|�d��Y���	�,C.[|�D���4D�<��Y����quc^�hj�Z��.D�����.�9��g�d�6|B�F-D��0��W���
��Z.,ƉC�
-D���� ��W(2�z�g�)��Y��j D�Dr$��Mll�U�,^&�3��"D��{я�-ވI��vx�qA��!D��  �Y�\�X+�D����3D�pD&9J�H�b�Z uYQsN&D�h�4d�%"n(��N]�-��@H��/D��+��=������Ǜs���&�,D��x�m�!�&F�7m�cW�*D�:����,�,���Ĭ*���r0)'D��ط��K���!��K�b�{&�?D����0Js�<q�*��o|F�h� D��b���BrD�@KX/qvq(�D9D��0�EV�5�h�'X1z���Id6D��@��81�v$0aA�(v��(��3D��[ri� ���P������c.D��0d�*y��}X�%�M)r��e�9D�40��̵ud�\ȗ ��:�*4���6D����0"��{�얝K@�a�H?D��˒*��H��quDY��.�AƏ>D�\��`��o�����W�1��y2k(D�d��, XP���HT'`����G)D��@oE�:��x�m&zP�q��;D�� b��S
�>l��Ex�nE�T�� �$"O=�0*ǒh�ɫG�* ��3"O�e(	�����A��$a�(��"O ��3�+/Z��9a�QPP�H�A"O��ⴢɹ;����Y���%"O��2bą�5�Npط��%��y"Op�*!aH":?"����W&�D��C"O�=s6c�; �D�!+�5����"O�陃U��I�ɖ>�؄�3"O|�9����5.�|�����#żEI1"O�L�  �PU�e��%׮bτ!�"OU�et�AQs�QO��g�7D���k�I����&ݫuot�p�"5D�,ہO@�.��X�H!��
��4D�,r�H32�FAҶI�?gR��%D���E��;]��q�g�6b�R�ȓ)D�0����;N���@�;Lo\%��&D��9���Pl�!�����y�J$D�8��i�H������V@�����"D���
0gJm3�,S�2)Y�H;D��v���H�2ɡ��ʥD{��#7D�(�dVa 	j�䊻#��<*�g1D�(+Q�xd��Pc�������d.D�\
���XO�q��<[�J	��./D�D�cG�6Ě���(@�n�4qG�,D���3h�<tb�����&��ۤ	+D�@���ׂED�ٻaNM`ۦ�	U�'D�l�aT0BrDX���5Ϊ��#)+D��;D�**�IP7[�SŦ͡��)D�4!sn-�"�iہ5��E��h,D�@/�-eX�,O���E�@�(D��0��=1O�m�R�W?K��Tٲ�$D���K�&u�t��FF@=�����"D��2�aI���P��NN�6M�'�.ʓ�hO�*O�p�be$��I��S�/g�B�	�><� fǆ6?��i�D�	!��B�I�Fl�	@1���8�I̝W�DB�Ir��Y�T
ٞXSЈޭ~D�C�	8����T"	�8�1��_�C䉨R/���U�TS��F�C�I�+��ҷ,Y%�X���ץK��B�	�K�PP�E�Բ)�1�7�ҝ(��C�|��ʢ��Q�,����zB�ɲ6����v����(��"á*�&B�I�Z�2=�nԬtΰ(�I�:FC�I�N�f���?T�р�
!FC�I��|К��P"s:řR��i��C䉸q&x`�M
-�欈"׈`8�C�ɶv"u	ph0#��`�u�ʉ�tC�I�t\��k��mv�I��� o0B�Vj��0�.E-g�[A��t��C�ɵcԆ��Rn�y�H�P�	��.B�C�		U�*w�؍-��k�LB�vC䉜��ɇ��;%�ԍ���a�VC�	�;�x�[r��4|�!��O�R,C��,*�E������T*V�]��B�	 'Etd���J�����(��B�bU`��զ%O�U�CC�kK�B�	)p������* F�����5�&B�I�W}�M�S ��]~X%	B
�QkB�	����F|�P� Ug�(<��B䉋_����lh�i=~V�B�ɺZA&@k�� GҊ���Ɲ*B�I`/B푲/K4dvx�@ED� g�B�)� < :vg��T��q2�#T���"O�@K�/\.p���X�n�i�"Ox$aB�^�=�X��!�9�s�"O�Hd�ծ;� �0�oGgl�"O�a���03�Y5&"O���s��Gβ���B:(��t`0"O�2r�Гn����D	B��(4"O��ޞE�����)��Ї"O������jl�X�.�~�f�)P"O��ӱ��\�J(��"Y(�"S"O��s"��(#=F���dBK[.�� "O�
��Q��|Ô�ګBHD���	H�O�|���1W��$"��ì����',X���;j�q��ۈ8�ʀ2	�'p���kŨJ�^�ْKH+�x�
�'���fcϯ&$�yA��/��-	�'�uۥ~����sN�2#"rњ	�'3r�����6[t):�Fޗ��`p
�'̡3�Q�R��RbN�H�Y
�'�,��pLT#`���Q��@y(���'����UjY8�8���aFq��'�Rt�ǫ�����2�ΗX1,͘�'��ڵMȜ�xe��d0E8>y;"O�� �N��� ��]s���(A"O�D���\,Z3�\���9�xX�D"O����QRX ��FU<
��0�b"O��k��5WfpR�*S̤D`@"O8�%�I^�@��(�`d��"OL58a O�XqZp$Rp:�Yق"O�-��
�G��%�E#^�7d�e"Ot	�s<w��{TbMF�
sP"O���|��5+�Ɵ4�Z!��"O���T�/��� m�a�@�"O���ѐ@b�x�+�	��P��"O�H���
.h���2h����P"O0y��XP�Xh7�ԜNw�-q�"O$�0������<D��A���r�<�dgL`�إ"�c@+e+be)2�
Y�<1��_�u�8!{��Ţ�P��KT�<!vm�t��Р��#�8є��f�<�A�?���bJ��tM��g�<)rC��.�\�(�j�e�6���d�O�<1�`��0���$��:�AL�I�<� �љM*%�'�?jPV%�%j�H�<5�Q��i�G! DZ�HIG��Lx�dDx�#�"i/���a��33����Ê�yҎ�5(-���AF��7j�.O�y�e�J&Б%�E ڕJֈ�9�yR�י&���ZQ��>`ni��Gҹ�ybM�1r2����4��A���"�y��ַ[��"dʕ'p� �C�y� �u�!kuN-k&<� ��y�C�#�)B��ΰg���ppD[��yRV'/����ܧH]H��K/�y��Y�1=V$ɖC�:0�5�5���y"CL�m&��A�*-Y����oY��yr�Ȗw�ہm�(<�U3�yI�Nq��؆p"��V�y��W�Z�,{��Z��,�h��ǻ�yR��NDv��'�V�W��4�L��yҏC=��I+q�S�QY+̈W�x4�ȓz$� ��-2���L��!Iz���0@=��ݡ};���w�F�`|Ʌ�τL�7�˟t��a�B����S�? �؋��1���(�J!/�4u�"O,��PĔ�FO�TC1��4J�H��"O&h	�	��_+vA��(6۬۳"O����e	x��`�!4��M["O ؑԩ�1ڼ�8GQ��h�"OHDB7
 ��	�����Aj�"O��ؕ���w&���5�ΛA۪�C�"O��;7�{���5䎵h�h�v"O��4�Ŵ	�ĥ��WX��x "O�-��
#2&j=�c�7*�X@I�"O��[��-�^�z�XT�2L8�"O���ƃ1U^U�4�R;C�"�"O����
��uJ��h�(03�"O⡒�j�(UA��*>����@"O`��x�轀�׿J��E"2"O<�"��d<>����4]��rU"OnU�ѧ�)��0#���)�i�"O��2�Y���쐷	��|�����"O䥉���],P�ٖ�Ϥ��aS�"O��� ����-������]��"O�\It%��#��P�@:���U"O�|��H  E@TZ�e�)��P(�"Oڌ�@ä?�l�P��J'�5
�"O��xE�Ź1�=�DBH�|/�e�"O:q��IEy	x|�5Aӗz��L�&"O�|�g��<��	�M�=Ds����"ON`��E-ލ�M��V�$���"O�d���9Þ��Cʍg��d��"O
��2�T�v�Y��tJ5��"O�E�,�%@*�QT���d"Ol���C�(7Fmȧ��I��4��"O�-۱ώ�m�8�ѢJ�>��8ۣ"O��0�Hي}���pi�"*��9�u"O�a@%'�^���k�j�%����"O��Pfc�VL&��lٮ0�Ƙ�q"O����W�	jl�h�BӈCp�X��"O�\1���8b7����M���a"OPU`�\zT����PX2�"O�����g���d�8t˔�!�"Oč� *�����!,���b"O��"v�3Iت����V�DA"O�4*慝�l̅�"��~�Plb"O�p�爈UP
"��W?Ob���"O��#Bj�:7�~䘧H��P��[!"O΄�G	�.j���)�RiY�"O����� �ڡ����w�b3"O����K�@��-;���MN8��"O0��7J@�z$3�dLTz�C"O�����B��]���ɘK0��"O����
��tbt`̙����"O��" ���8�EI��ق6B��%"O�L+�	�$�$	�JJ-!]�:�"O�<�[� �2��%Yl[�"Op	:bN��,�P�WL�>oo���r"O�$ۥ��/VRbj_�iL �v"O8��E���H��90J����"Ob�ʓȉ�=��Dr��7
F���#"O�]��D
<F�r�H��L���w"Od��#���e%�l (@����"O�ȫ6$��g�pD�eǅر�"O�tsfI�%��-��5p8a��"OR�2��C�8�U�E�?l��H�"Ox �	��&�ZT�Bc�r]�p"O��SU�>w��C6d�4�d��`"O� ҁ%�]�p�ꁃS�th�9�"O¨t�		^+���S��)�"O���LZ�,ۦ���ˆ���u�"O���B�*T��5�3kۅT��	�U"O��
WX�d��xI�iÍvJ�"OhabR���H�0s��V4'r���"O�mI�%
)m����n|��"O�L�iz��q�$L�9@��@�T"O�\��%�m�Z�$��*M8��"O(d"Ǔ�v�T1�sK.p/�<�W"OT�#'�ʚG��b���<�95"O0в��˥Z��d{�G�S��P��"O��r�A�ʲ�kq��f�x�"Oz�P��E��xs���*t�f"O�DG�K�0qP� ��8�"O���aԵI5��@����w�3�"O��� IJ!e��s]7�T���"O�X��P���|��Ɋ?�r��4"O�a��n߽Y^��C�#̢g�"]�"O�@@��T!]���E%��j���3"O�H�dXPW���dT9Y�Ȳ�"O8)�T(L�R��s�M�:EY+�"O� C�ܡ&��P��I�R�()�"O���R�/�
�I�o�'t�x�"Of eDӼs��=Q�->;�@v"OzmJ�(9�d$K��C#<��"O��DK
��ٓeh�Em
q�"O~8����oI�]���џ<���s"O*��u&�n�(cG����D�"O��� 4w� Iz��&lî���"O�48�eY3<L���W�/D$p&"O��ҥ°?�ZuY #H�Q�&Й0"Ot��F�H��S�H� �I�"O�Y)��Z:GM��h���9���C"Ol,�ƢO�4<,ɢ�ٔ0�&��"O\ kZ%���jBB� �8@�A"O��R�bǐ&_F���f�'#�܅a2"O�\{tI�!4�2���卐=�X��"O�@�PK��3Y��sSE >�Xu��"O@��A�)^���ȂCL����"Op��M�^�Q2hٰ<��hP�"O���V�.�$�c�U��d�v"Oҍ�\r�P �h�	/=�Wjڅ�y�'ۥ<�h�DO�����f#_��y&�C�������H�7d߶�yR��G�(��w�E9m�`��.>�y��VC�n@s6�ҵs�x�����y2�դA���`1	�d��uJ%f��yR&��	��I�3 `+�{%���yR+��
<�&�Q�uB���:�y2�x�0�v��+=���r�����y����^$�R0eR�2��8ܠz�!��\�G�p�A�^-\6-9RǒL�!򄍨]ִQ�m���7\<F�!�qG�k5�U@�z@�0�Z*�!�՛0Xԝ�6N�F���Ck� 1�!���Sk4�&���p�^�#B)AY�!�d�3- �K�0r��`�Du!�$��AF��'D�U�P��
!��J����g���;)$�ԴiN!�ć�fV�S��^)����#(S�!�dã$��àb�-����˟v�!�u�P2`MA�g֤-(��Z}!��[.F0�A;G �14�����`֘u�!�� ��b�-�0 P���Bi�]��""O����&ބcW��	Z��"O��P�n��'i*��@甕J
x�"O0�B��_�j�[�*e�n%��"O~Ț�b�r��j��/F��!�"O�4�3��/}�)��Ĕ{��5:�"O�,WL�>f(E��#�<G���"O�@*֯�-@j��7M��f&`�x�"O�#�Dhf��ӡ�2�i*�"O��҇�.(Xy&P'a��0��"O`��3a�}]�9{�X4@���s"Opx��2��0��ЈO^��0d"O��0��CPF���˙1/c���"OP�PD/C �B��Ѭ�����"O��A��T}y��,̈́r:V�r�"O��&@��ڀ)RE���2"O�Q`���<~���Lz�c�"OhM!7
&��X�p�"�l�z'"OJh��j�{|�*v���p���"O|��
�Sa����H��Y�Va�"Ob�"��"�2����Gu�\H"O�y���Y`��1�G�jX�p&"O�%3�����Q����eC��	P"O�ňf�:qN���n� I�X��"O�����/RO���GlX2��'"O�P;S��K�2��*�b\�d"O�՘���������4Qy@"O�4�1hȩ? 
"���B�I"O�(R��-q�)�J�!@o*D1C"O��̟���1�)	%E��Q"O�9�P�A;�mRP�Ƀ7�i+�"O�092f<_���dS�v�d	 �"O�R�#�,#��
���^��	5"O���c�E X�*6��2u���"O,����H��ј���Mh�(��"O��SK�nO�]7"�tLx�"O����ѓm�`�va
�7��)4"O�����
0�x1���}K�ȑ�"O��rIS4
bL�� J�=|yC�"O�M��#C<��e.�e!j@�1"Oĵ(U����GM�|@�9��"O`%K6��ސ���G4D
��`�"OT�A'����: �R��.��D�"O��Tf�K�	ƥ
z��P�"O2� p슗*hٔDS�n�T�e"O�8�iH����>�vl""O.1U6k��i˳�,p���"O��3�E	�I�G��r�|�"Orq�Ð�s��L�p�E/�:a�"OrU��کG�&�0#�_?T�X̃7"O�f���"ٛ�� N�Dp�a"O�l"�W���"��_�u��\�7"O��$ݘ{�^ �V�6Ū	z�"O����Yk�"���Q�xYˁ"O�9q	��Zw�pq$E�	`��ѱ�"O�H��ۘWL�7�I8JȌШ�"O���"��]�Ӏ"�i�b�Ct"O`1���r<��B!#�	S���"OPA�.V�cVI���U禔J�"O�a#�@n�ܐ��C�,��sD"Oz�6�N�.Z�x�e�:|��J�"O���u�P�^����b�дJ�d}Ã"O����JН
��Ȱ��	N������'�'���`J��R������_ 3]�$���� �( ��Y}���B��-��u��"O���1 C64 %�7!�F,�u"O���Gk�&Z���B&��<H��]*"OB��į
�beHF��]n^= "O�|�4-��;��8�&�{V��K�"ODxb �	R��� �D/2Q�����'��OuB��
2��H�GC�"M'�4����xE{��'��'�l ZP�=2`�`i���qp�b
�'P@Y��
�e��1[��e�
�'�{L��k��QT�H8Ux@�
�'.a�VY;�h�#�4E�	�'��R���	���w�ޝ��Z	�'�]1��;@;Z����ܨ�����g�����ȷ�����O!�D]�[�`���:inz`hӁK*=c!��R�1��-�B8��0� @�V!��J!U&*#D��peI�lo!����d)C� T�u���CI�(xa|��|B�<T|���]5}w����(�yB�ݐ'B�פ�������x��'TxW���*X"�fӛ	�.��">D�aR�ͻ�ډ���-jf	[4�6D�T1R㒇��E��S�@���4�0D���a ��:��T�$R�~f �`� !D���c�x�$��
����T-!�O@�w�>�B'�ɠ��	�È�$~�.$�ȓ^�p(U �z5\bE�6��l�ȓQ3��	�(�)*!lB�@��q�j���4^��FFʕ2��%��q7�aM�m��ه�͑$����[)� �pÈ�,�	�2�ģ9����!�Ab1$+� 	� �i�$����?����˾� B�V�dD~hk����hO?版��T�&�tJ!�sȶc��G{��ܒ�'��ٺ�DHpM<P�3 @ �y���9O��q��:o�d�B�+�yb
��d�4m˅N݂mW4T�s/��yB�05r~1�Ǐަyd�ɁV/���yr��4#�$�!F�"y�b)X��Q��x"�'^����B�������âZ;Z� A�D�O>�ub��Aw���aE�
15�H�<�����%�ބqъ�dh���!��!!�Ė!L�U�'��Wܰ�@ϊh!�D�4&��`��;rxM��.W@!�$G�Lș< �@���D;x�!�T}�|*T�ٜ���W���!�!�C"���ݟt�R�����~�azB�$Ke �RDͶ�,�$Eۃ�!�W�w�����'>��8vɂ=!�d�!RTkGnJ,��1�	��!�D��f����C;sֽ`dÅ.E!�d�#���31kJ�p��x�����A�!�
|�����mD�pl0���Ƙ#�!��H.�@XB(î_���,M�W�!���O�@;�+ۻ5��d@�)�flJ�8O^�d�<�)O?K�Ǖ=��afDm���Lk�E{��)*{qb)�Caܤ$���XH��"O�q#H��4E fg�$ �P"O�p0���5kKD �ֆD&a	й�"Oz`5�ބ/ P�:R�ɋ�����"O�D�V�X�]!������>$�"O�@rC�Ʋ�t�ps�'s�UCǜ�4�'�ɧ�:\���#�P`!C��,�֡�%�!�S��y*)U�P ����$zP8�9WC�#�y
� ����ߎ3�,�k#��g��L`�"OƉ�	��be�BH���h�)�"O��@���3W�J��ȷ��8RQ"O袧!K;F�<���1Y�9�𗟠D{��	�!뺤��O�Jɰ}�5��7C�ax"�Ia�Z�Eʿ5n�:v�L-a7�B�ɏ�ŃP撎/:�<����4��C��-8�ѹfFC.��2���fB�ɉcd���W( l�Ie �N�:B��2�>]�U�	�<��}�-��]Y@C�;^�����<W5�Q�a ��I��1��4F�>�(ǂS�	��2���FD0"<����?�����{��9A�ݨ�|���� D�x:E��98�8�Tj�pwx�bC=D�$�Cm�*ڴ vhX:L�f)	��/D�p)��\�R`�2f�jv��gJ/D�ثv��%��|�QZ8Ɂ%�2�ON�O�����	�<!ȓGU8����� ��}�'����0�ŋȜ7�4�y��O�5�%H.D��A!fK�-�J��B���u�̐Q�'�I\���Or��U�P��L�y���'Ŭ5�1O�y�5�+2�@�A�Ɍ(�-`T"O�3�9��!,̟�H���"O���%�1vL��+2˾)�T�'��v�Ja��ZE�7EW�~8���'�2���p]�XG��?��#E�0+!�d_�^�]#-�Ɲ�acŕ���'��>�)T��"�eۄbY�+�P��6�<D�<�a��H����cE�) n���'D� 0,.��!�1Q�b�hr D��u�C�La0�1/ 1.�C��>D� ��+F�Z�ex�$��C@>D��Kq�8=�4��O����-�&�;D���w���|�s���D4��:�N4D�`� 	?$,���ޒRڨlw�>D�0ɂ!�	cJt�# �0}:��'0D��##'X
�mxZ�a2@PL��B��/1��؆��&=;�))���42�B��$[�\�Q�ǝ�?�`�H��^����6���^��T��	=C�B��qǝ�,/!�dL%Jdz��1���#��!�Y�@Q�h�7L�%*�FS�K�F\!�Z�/$,�{�d0R�(�I�9!�$����%EO�m�z���荚,!�DZ��8g��L�xGg�!B�!�A7S��-H��ʱڰ�C�G��!򤒉z�򠈑ĘC�,�	%��F�!򄃞g��Y����$�zѡSɉ�H+!�/bJB ��� H,����� -�!�d
X�<�b�]g���&�͘R�!��*b�X����6B�|����1.�!�$@�{��,�Eۛ9��Ty�  �!�$��İ��Ҋ/}���N�.�P��$�O��[݋Z��pK���*T�P�@`��S�����<զ�`��:KJ�Bc��!���wx���S�
"@z>`�bÊ�
\��;D������Vv�0�OU��2�÷�3D�, �L @��8B��NLgС���5D�t!�b��P:��֜=���[�.���ɪV44Z�n�
s\�;&�1g��B�I�GĨ�.T(8ZgU�:�"%��5D�D���U�J1���ߌE�͠�k0�	lyr�i>�XwaH&h X�N��_Ʋ��:D�|���Cs��p�ǎɢur:���;D�� �|i7O�;\��[�ç�^�6"Od�YE)Y =��18����?v�C������I�ۗoG�~,(`��ߩP6:Y���/D�l@�J?v���Xf�ېL6�8#(/D��{�	<d~m�cY�9KA��'-?����<�N>ͧM�<����_�~[3��R�؅� �ԍ��d�17픇Y,��@�� D�T	 �F�Tl�P2���N����=D��IC�K&�9�eK	$��02r(:?Q�o#��(jS^�<Cr�LsGtņȓ�1cq˞��0��n����'sR��ӫi��o�U�"�Y�D�h�N���>qE@E&V0�e��PR��u��ne�<�Q$�"��e��0wLN�R�EL�<��Q(�&�rD�A/.,�킰��^�<�Af�3[����n�((&�Т%a\�<�ekQ�MhN9 s�)[*�R%�^�<�Ϣu|�L��JY�Ih����]̓�hO1��a�*�59� ���'Ud��1���%�4ړbe�%�hݵ*��%� ��-����ȓ|����G�D�HKGo܅D)���ľ|��$Q#v>�}p�hJ+4؂)��t\�� ��Ͷ^K���C>4�����z�ɼDސ�{��B.*��ڄ%��DM�B䉹,�Hb%HQ>����@w?PB剗z�4�b��H�K*�,���P%f�G����.z�Q�p�
��9��&O�y�g_�5��{׋ɍy���I�y�α��(b�T#CI�Dc�6�y��ԧ@q�8VNE$|k>,��m�y�$ ,�Э"c�؂���r�h��y���o^Q5�/D����$�F��y��5�2)��ߣ
nD���yҢ�4<�t�)�~°�� aD��yrL�6]�T,A�� xQ*�� ��y"O�@�H�{��g���30/O��yB��Wf4,j!�_!�-���˭�yBʎV(x`8�➑B�`���D��yR.�>����'B��a�ӷ�yB�PѲ�ie��u�N�>]�!�%5D�ȊmI�=<i�#m��T�Y��(D�TZ�fFT�H��F�!Q>`C�@(D�8A�낑�,ac�e\1g�6PA�;D�D�p��1�gڈo��sC%D�L0�ꀉ+�P9���V>`����7D����Kͻl�y�"�&C��Y{2�4D��9��;m���j���]k�d8D�8Rf:z���Ʉ1s�]r�l5D�̛󈉬���(���u�(h8��8D�<�� E�R��@V�a�\�ag*3D� �6ƅ�b����֌%xDd`� 1�hO���n_N(ZW/O;w$��B U1C�	�0ڄ�r��_6�)bl 1Ud�B�	u��M��/U9;��Ta'�0~-TB�I�b�����!��ʅ �>gP
C�ɩ3�4S�� �
DClH��C��U�b%�"��5%ॣtlD���B�&s���؁ᘮ �jDi��1gzB�I�J�t4u��)_rR�r�F)\�C��4w�=K5��04�fþņC�ɞ;fYҲ�[<;��haR�L�B���4ړ>��$���^���ݚ3$ݥ8ɺI��m� $����]XرB ��[�|A��PWx��5$��{@`$��'#$�L���?� x����P��2fX��z�Ҧ"Onmj�ɚ4tn=�c�6cqt�x"O�r��� M��8��$׌*]N�8�"Oڠ�"�9n��;�_�<x�ం�'8�O����;`��k�kS�?N�}Q"O0,�U$".��Ъؖn�� �"O��HV`\9�j0C F��%y�"O��jUc���!^3[�ء�D;4�p;b)A�����	X�~t��J$D�hyw+��u���-�"�FX�'6D�Hu�$BŬ&(��*�x `r���I)�(���np���Ӗ�j�C�	:����q�K������B䉪+S<(2K�>?�t	2UN�`-�����O0�dۿX�䱩,*I�QY�O"^!򤊀��1 �<���A�V�yO!�ĈH�Ȅ��/^�!�\ �DÑ �!�D�P2����/zt�e �a��kZ<�lG{ʟ��W8
xR�� �N
͸6"O��8���E#ZX҃�3�iI�"O����ԾY�qJ�n��u|���q"O��2�h �v�`rM�)7�4A�"OZ*�=�¬;���_�^ň�"O4�h��ŗp����#Y�`���"O"(��[�����B��D�L�J��	N�O��)���ĞF�Ƽj0�Kb�D͠�'-|�Xb@�`�k�j
d7��'��!�~&rLkG�V�a��i{�Ov�=E�d�Ɗ;0���f+�X��)[��yR�
;=on`a�K�4]>�ի#�y���*�q+�� ��p8�.�(�y��;f��z!B�7Sd=�����y����L��E A��; X:��7���y"�іj��t��dX}*�)��ǫ�y"dʙ"0��>�����R�����O��"|���R�nr~(�f�zp�]�FV�hO?�I=A"��veU�֢$ɑ��'%ҰB�I u:1H@�ц4HZ����.j��*��2;�Z��d(A�� @�m�e
bc����S�\h`��Mzd�8{�C�(�Lc�܇�L0d��`�Py���$C�ɺY!�I	"� :
z�A@
��>B䉩|8�b`�G�)4���
U�B�	�P��{��ƢZv�y�,�Y�B��x�"�X�(��zp��=j�����&�	&���X��8�\��rf����B�� ��q�+U3.Z�r���1�b�`��I&���#�E Z��y���Z��B�Ɋ_ �˒�ȭX*�Xw��9oH">q��I��T>���SL����ç 1O ��+<O6@[��F��P�W�6�FQ"O��)%�"VF�بU Û;��4�"Oj���� c\(��bƶ����"Ol�hM�����ʌ ��z�;O���d�/<nH����.a��Z���C�!��S�4�)����pE��ysH΢E�ax���,|�����CP|��.N/5�lC�I�m9�Xʲj�}@@x�ר�=O�>C��=c�dx"!)��'{(X�����OVʓco�4�����$��0����<A���)�:.m+G�e�2�à�۾Ze�	gx�� �X?^N�e��vQd`�`+D��:�g-e;d	qAX9R��YȒh'O.�=y�ҋ/"d�&(��O��4��f�<� �H���B:,�n}�V����V"O�q!��6Vw��t*M�WRz b"O�(�!l��I`��!�eG����"O��E��uPn���m	�@V.y�"O��:'!�*L98�����|'2��"O�xY4��`���"6BB
_B�i��' ў��.лu�>��`�Q���c.-D��a�_2A�J�R�.
�P5�0D�����P�����H�2+n`��0D�HRcěXMX ��DD�k�j���-OL�=y�D�ļ� g��OG�!���U�<�s&��0�
�t�B�a78s�T�<A���jXD��^I�f�Au*@P�'>��ӌ��Ȇ`ڲQ���UA��mvB䉝5qj��ѣ\�@��ZB`X�j�lB䉃tS���Rh�fo.Ehbf�WM`B�IsS��K�'ųO�
�p���r�$B�I�@��a��aP:#(�T�Մ]��RC��=!�@�
�p���*���]�B�ɯ\C�pGAU�5��T����Z�C�I�o 0bdlF6Q��b2�./��C�	;@�D��	Sξ%��욾u>�C�	y�ڴтǚ�-z�K��#fo(C������/٤U��	QSFP3�&�E{��9O>L.4ܱy>0L:]Y!��)b�!�d�;��I�§�%/G�UY��I�c�!���/s�A���U�DW���m�6T!!�dX5Ҍ�c֩�+2��C��!�؇@�Y"�kV�/��	�$m��mH!�d�.v�%��N�6����k��.5!�Č��J�b� �d؁�W�[8!�䓰�Z� �K�J��d�O�h!�.Yg�|�4��2m���e�Z�!�d�9?�z|B�+P ;xɪ��K/�az2��8΀)��ȑ	ON�풓 _�V�!�Ċ�}�f��RɊ5v����/Tm�!��f�B�2�
E�d��L��!����yW)�8��h 3bQ&N!�^�W�ve�WNP%*�A��5!���>_ҠF��4|�#�F�[%!�$�a��I��"K�A(���6���a|�|������ڒҷ5�!�D,�	Vz��d�O}^h�� �!if��@�M�W3!�$ح�L� ��P���� ǭ %!�J���:CB̐Q���B��1`z!���Tm�D+0�O�D���⇥J �!�d�.w��A`��;#�"��)�!򤃥3{�R��Җ_��5ɳ!��V�!��aΤ��5��.����󍄤oR!�䈘Z�@Y�b��+�z�r�L�!�
TJ!�E�6�*����04�!��H##���a!R:{)�M�ug��'�!�:C�>�KbA�5������#�!���y$B\c��� Ӧ��F��t�!�DU�W-�#��X�s�>�A��52v!��W��U�G���LQ�[q!���E맊݉>A�����ʛy�!�øǅ�0C7��s�DΚ5����"O���"��,٠t���z�,�p���O��=�O�<��Ɓ�"�t�!��T"U��'-�t�d��ℊ��^<N	�'�r��U�\�0f��F���[TV]�'i��z��]�-�	˥BP�@r���'���q�؝R����%�F��m
��� , 
�I\>e��DK�	�W�lU`5"On��􁎰�p��ώ�,qXe�"OA��Z{f�#.�`|,��"O�0q�=,������H'bW��Z"O���%*S�<Ͷ<���ٝok���2"Ol�yFlLX�V�)7���.Wbx�b"O�x��
�!�����N�
�ڧ"O<À�{IV��e�E�rڦ��"O( �˕�"��<Ag�@��x0"O�@%H�<�`�rB�D�ڜH�<O��$�O؀PB��y�p�T�ג[��(��"O���ׇ�ʱz��ig>t"O���Ҿ)��%a�S b�qhR��O���/��"�K2o�}�nɀԙɂ=�ȓc�%�ִ4�r��2�,��#D�Ի�e
)a�v$�@M�^����P+!�O����O�!�4��u�j��(ŻL>���"OtM£��\]R!���
*޵�"O.��!Bxt�!q X�	J&�9��'��I�Z�H2oL<cl����|�^c�h�I'�D�����X0dH�D`��x��}�!�X��y��)�';O,��d�W4��@��i�n��ȓBt��J�-D�p��QH�����yy�'��8cǇ�<��<���6���'0�h'ũYe$�r	$�;�'RT�sd�,:K&�B�����X�'t��{��^�W��J�I°x%�d3����O�㟤�O�)�s��8:��x�`�۔x.<�@ӓ��'_L�jϬ0����_2v�*9��'�lp@��i��9�pDT-rNJ|b�'���x�g	�#}����`�����
�'/�����Ю<]j9���N��B�'�ΐ8�"ڶ#,M��������'iht�u��%*�z�1�ț7�ĩ��'��Ĉ7�܍f�#Ӯ�-oͼ�����dƫ-����NW � ��!�D��<��I�&W5B9@T��p�1O��=�|��ֱ2;�Hp�Ί�
���ҥ�`~��'zb����#Y�Y� �T�Fxڈs�'�1�'�:=���6��B=�%��'Eh����+�΀��@Κ@��Q �y��'"��
��;�m&���)F��;�'�i�g�L1n�f�U�P�1��y�'b\� C'�!<OҌE	�#t���
�'�0�)7Io��=K�����T�	�'���D�
.ou�$�փ٥�rh	�',�)�Eݱ"X����(�9 �
Y��'j�lѕ�QW�\q�ߛ��-��OF�d2�O�a�v�7K�$ Ƥ�&P�e��'�&�@��ѐ�`�ȴ΅�Gt81
�'�5��lНbwi�Bd!I�J�

�'x��	�(']$�=s�J�-�����'�@�ꔆ���!RS�E--2�C�'6bQ�@��d�T��g��)�(z�'�Y����@�J�x��>���	�':*C�oߨ-�Aw���\SR�Y	�'T�I��@)7�Ay�N��'�8��'~n���d�(�0�E��#�>�b�'B @� �2��D�����'��<��g'@���A]2L�d���'0r�!�΅>��h�􄒔H �h�']Bp��"RY~�I����p��'����� � %ZlQ�	��s�n1�'�� "�#��S���Aʋ6;Ұ��'�
� ��$$߂L� ��t���50�u�d�'n�ɂ+�L<*��G�+>Z��r�C�M6�	F�����F��a�6r
4iD.?D����B1j|�I���H�*�����<D���ٯ`��S@d�7����� D��"��:Պ�"��7(�����"D����$^
mp��F�:2�)sd�+D��Jg�K/k�p8K�l��X݊t+D�����m��tx6,����3�;D����O��h"D��0����.D�	� �| � ��Զ"}R�Ԏ:D�x�`� j��mp�e�	� Q�3#-D���� 3
	 p��Tw
�́a$)D�ē���t�ZP��œ�a؀-YDd)�[���Oy�p�AlC6�Y[��8S^���	�'��iSFG�o�Z�Z�
g�4���"O"�{u�ʐ
 d��l �B����"OL��p�� Q�l�k��204\��"O�ّ҆r��-9��(>Ń�"O�MS`��(F:JT��J�3
�
]�1"O��5K�#K�|�I^oj.=Ғ"O�9�M�.pp5�r�Y.@y�	ڐ"O�=ȥ$&6����ȶxwp�h "O6�"��W,䡴.�`iȡ��"O,؂wo\�n��IK�E+$���"O:\��A��tVpQ0
��0���"O�4�2-B�fvY��I�p����"O� �� ���ᑣǁ=�
�J�"O�x�Q���/<��p�Ȗ�20>qBg"O�!�K��S"B��
�.b�!�"OpT���ʡH����#��8��Q��"O6Y4�ΑN�<0X5���L�(�"O8Q����V$�)�rb6U�����'�'�Py���>E�1;al`yD��	�'Y�!��-��[J(-�1��^:<D��'�>�s ��V�����IT�}��'>q�4�Z T�$<�3`ɄI��i8�'&�=��k��D�3;��h�y�h8GϾ)���2i�ոG��y"̢�`�b�1?&� &M�;�0>�J>���(gZBa��L�(�:4A�C�<q�aE6?���Q�	��z�Ch@�<i#�ƙ Rn�:�DS)+�"��w�<��C�
9�m��-��c��L�#ŕL�<��O���� /�#ps��qg%Go�<�	��(���c��u
�t�u��i�<�W�)5�&���ӝa�*|2���L�<�VBR*~��IA�D�/���2���hO?�ɒ�t�����/N�8H��Ԧ�B�I�Ml�
�k�HD����e"@�C�0S�p(+�.;}�d̑�*(��C�ɞ�Z-�fɘ�-b
}s׋K|ήC�	�(�����k��#���"��s�C�I����(�:;�� d��UR�C䉤f�� b#Q�g2İ�c`��C|�B���us��F$M^��S��HV�B䉸/�2tX���+B
m<�0��'�f̀R!S����IHȷ3�0�'�D��G�%(����գZ�zq:ш�'���R�^'"��h��Z4b��ha�'�TأRK�=V� �58a����'�����L*^iB h�R�L�ri`�'�����ً[�d 'g��x� x��'3j�%/$��}aE�Ķj�9k��� �@7�&d�"h�d�0��E2p"Oru��*+N4d���ݝ��ja"O<-R��v\d#�AGf��D{�"O� IR#�p$��س���f��"ON-�ǃ�^6��u�R%p�)z��?�S�':?�$ҀK�Y?�58���L"HĆ�"R����9��!ɰ �v�ȓuw Ȫ����U��4A��X,"{ ��ȓp���G��$	||��ƛ�9N:���+����U�9y$I�p�����0��)Ct-�
5Pir!n� y�q��T����/JWgjܸΘ�$x��Y�21��-vV�Xc���А��m���+T%w�� ���uS� ��a���1���Lh(7��B�}��E�$�"CM)�)���ƽ!�8���+X������i��PmZ78��C�ɗ\,�8�a�=V�H�j����rB�ɭ!EX�"�.f�ڡ���ʸ4{FB�}J��#�,Lg��Y���.�
B�	�g(�꣣ޟe���#�B� n��C�	�����aʊ3��m�@Ր)fB��	\�UQ�� %�t���䈖w� B�ɲjf��0�=r��s!(����B�	�\(]@��$	趉��W�L5!�D��3n���bJ�3ެ��6a��!�d��u�\�P�đ�8����ף<=!򤗉"��jĄ��.�Ɋ�E6!�d�-e� �sOՀR�½A#銈�!�����=��l	�
�ؐ�ۛ!�!�䕢1�:���T�'�"��ǆG�$�!�L�S|���O&��5b�V��ax��I�yrv�1cm_r��M�,�C�&fd��)VoʮI��\� �Mo=�C䉗Q5����?/�¨�3���ZC�I�)��-���K5F�t�� �Э
�NC�I� qL|�f��cWfQ�e��2c�C�ɏ#O�L)�R�;�j�P�A��B�	��R�+�Z�`q4}y�c��W{�C�'t`���#e�:Uܥ��+��o�vC�	\�0ܪ0�Z�D��MA� �NC�	#C�,��%K�&�؍��RN��C�W�P��Rl����`��]?*[�C�	�-8ձ׈��h�xY���{9�C�I�E�N=j1l�]H��DY��B䉔7����_�rdr�%�4��C�]�T���d*��٬8>�C�IY�P[��S.1
튲�Y�h��B�I�[�M��G�hA�)$�+h��B�I6���"T��:j �L֭��B��
Մ�=j� YHs<Ћ�EKn�<��L)k��a��[�,� +FYk�<�$��`*��2ϋ�K-���D͜c�<�Ӌ��,،hRsG�4E�Z%�3H�<y�n*�8�vOB�G�h"��@�<q�b[�r�N��c�-,e$j`oE@�<A�@$A"�3ĉ�='8��Vx�<T�X�~o��cd����u����[�<Q��=6������()�$5�� VM�<Y���@�IÅ]�MV�H�D�Q�<	cLV�47�I��h׵>Y��)�M�g�<�%�N�m��I���V&i����@�f�<!U�ǥbP�����j5n`*篛i�<Y�N�	��m��̋_Ȥ	Ab�<� �8Z��>Phu���P+ph���W"O&h�r����`�R�wa��"O|���"ѕZ%���`�{:H�5"O�	3�վ���#�ǴF7�H!�"O(���V����C�DK�4ġ#""O��9pl@K8���1LIR"Oܸ3�ݩfp 0��D�5�TT�"OR 15���q�V�+�Ԝ��"O�E���X�]u~D�a
.ebBq"O���W!�73�0J௃�A�1�u"O\���:�Eh���>_�(�c"Ou���0+�����ݜ2~��a&"OZ�b�ɓ�m�Т�)�0Zc0=�"O����)��s�>��W�Z$h8��'"O�}��B;~�Uz�
-]���"O�-�ǫI7*�
B9MO��bt"O�!�� ˨I��j�"Șb6����"O`b�7^��H*Šذ(����"OJl1&F��~�!�qa/n_|I�V"O�k6/U=5o�|�m�<��q�"OֽW��#)�pz���u�x�Ѓ"O���o%7�,�Ң���Z��c�"O�y���X�r�r��*�"�
X�"O�ݚ�D�A��*��U�xl���"O�0�@��B�1�'+ o��"OZ�B��>{�>L0Ȼ|�R��d"O���(�h���1Ę�R��B�"ORiz�nXO$0�@�`�2g<���"O�|I�@���	 �W�#M�A�S"O,��`G�z^�p�S�
	q��Tau"O��8p�
�!�z��!)A�Vb�}�5"Oj��E��%����'96Vx� "O,���@
r�p��л$L�4A�"Ohl����k��x5 �	m.4�5"ObL�B��v��UZ �K*;�h �"O���'��4)��8�q�B�B���b"OV���Y+f�E�⫗�3��#"OpH�*�3�r��!�ΒD�\���"O:�
���A8�cI���̚t"O�a�j ]3X�a`�A2qDP8`�"O�d��ԛC�dD�흙C�( "OЍ�s�4z!�%s��
�R��"a"OL�iG��wӘ�Æ�թ!�.��&"OΨ S�F�$���c,�\�&hs'"O�����W���f+_f�䛔"Od��F���(�	�Y9ƤB�"O�Ih���x�PYKqhѰz�9E"OV!	�nR*39�(r�J���"Op,��n�x��l;'�{J����"O��`F ,[6��a�_3d�P�"OH��ҡR:Kp��1�ځ1��*e"Oh<{4��2~����&��T,c#"O���mUHnd���Y�D-3�"O��dT3�t�i2�X!��,A%"O8��V�B�F�|���&X�����"OX�#�ĝ��l�)d,V/0���Z�"O���]�9���� {�B�
�"O���uC" �B�
Rd<g� Tz"O�4���C�n��x�`���d��X�D"O0�a�f� K�8���ql�IR"O<�Ӣ�Ӝ�&T���X/\8�`�"O. �Gr��k���h�.�a�"O^m��3�������N��h[�"O\)�Ҧ����c�O�
t|��D"O� 00s��-.#�hR�U9q�`�:A"O0,z�f܈�\�Z0wv�]P�"OD-��i2�*;�H�!n8
�A"On�q�/�������//��"O�Iʁ	��X����G(�*QX�@"O��U!�4}���V�8@O��RA"O ᨓiV�p����&E��H��"O��[�E�ZD���-P��#"OnA��ֳ(����
c$L�"O$rW,�
N�4��A�8r:�@
�"O�1�*Fw[@�Y�y[��W�S&!�d<`_*l���e�=����R!�䋩h����s��j��(2�`@,!��$9l�I�*F5C��h�\!/!�Ď�p��$QFE�+q ��L@5f�!�d�i���2��1�������*�!���=���T%P�`=kt-�<�!�D�"H�My`��ሤ���K�U�!�	�?��'��4�:��JV!�*�"�k��H\(կ�SR!���}ϴ�;���,]�z)ү��#)!��5JȠ㬔Y���GO�>8'!�˴�Z}�d�$ Xn�9w��"$!�$GPǬ˗hA-�xypg
/!��0>�@2�L�d�8�v�[�X!��[*�r�(���w:pe[��ģ4�!�$X&;F!�U%�e��Rv"ކ*|!�d��+^�y{�εF(�C���}`!�dx�� �d�������DH!�d�J�F��0EMg�� �@� !�D�Z���g�	C�,,P���1!�DU�uJtxP��B2+�x��[�;�!�Ğ��,H����:B���� !�DħI��y���Z��a��אoi!��oz���F|�p4�"V�!N!���\�J�� ��% y8B��{!�I�%)���x{�-7f=
 "OLЦ��Kz��'�%*Ϻ"O�5� X�R*��ydL��	��j"O&��r�MdδC�[$WA�$p�"O����W�i��}[�J�$.�Ԓ�"O�\�s�Y���Z6*W�fil�$"O����%' ��C��Y,ެа"O�)���Ӳb;�	���X5J'�"O��ZWa�b������B4"O���
\��]��Ɉ�%lm��"O��T�K+]h�}qt���#�$�S�"O��g��4gx␡C�*���"O�����U5�b���4;���*�"O�0�
Ȏ�|��Q`ѷ{�h0�#"O� �ȕr�� �X'"�r�"�"O�!����+4���g��^�"O�1��R4�����HŮE�#"O���aI� ��\8n&E��"O����U�Ă�P��Ф��"OB%�h��'�P)��2	7��`�"OB���j_�h X���aȩ;6��Z�'�� ��E?���!�-�Y��'�帣h�>�yz�A��b0���'����``7�ޙj��3WI@<X�'��J�o!8в�B£M5R��'h,�	�ۑ<��U��!��G	0���'*�V�^�(�ks瑈=�.܅ʓ�Z4���r�IV�ԙ2�X���S�? R[�N���<Q�I�u:��&"O��s"0�B���
�#��!z�"O�-��F	
63�) s��P�<ũ�"OdK��[�.�0T��I���`BS"O�`�
*iҠ}RG�K�5��`I6"OX�hqÃ=�@�U�I�ZU�E"ORM�"Ҳ�n��7�	;��Z�"O���1*ȣ} �qDK�e+�q�"O� 4��,j���1T�F��S"OX����8� A�),���#"O:=���% @�H]�x��A@�*O���Eo�6��(�n`ܲ�;�'�,��4�W� ��aC	�0 �|���'o�=��c�s��e��+T�(��C�'�v�3��٨d�e��a֏&�����'*�	�uo�-#�h�e��%L,��'�dٳ6F�np�4��/]�o�n���'�uA��O x(~�S��V�mtf�	�'��22.��^*�3�AW�6R�}�
�'�޽h���&? ����? �Px	�'^�l�Q�i5`��O�'q6�[�'!޽�'�:��A3��v&L���';�D��Ɏi�8̢�h�"a��	�'��5h҄ �u���B�mO
qR�'�:�4 �������bh���'l���"/�)pC��;��#SNTC�'��(�o̍g���0��4Wv��a�'LIb ƒ';�F��w��J�p�H�'�@����==je��oD�>��'&�|�n�-ɞx�0%X�~Ty;	�'4ģ3ޒo���k N؁o�"��'�F=S@A: e��{d	+j)dU��'��rӮ��Z ��d
��bP�=[�''�}hTF�7*�0	d��T^���'z���@�(�>�6��4c&8��'�fD��kU'�^��u��%c�z�@
�'u�+�j�Id�Y�g\[����'E$�y�T�tb��C&d�T s�'�Y�d�U�Jׄ��%��Dg���	�'������=Crf����V;4`U"
�'n��7��P�P�)�k�
]���	�'���y��ƻu�0��j�6'� 
�'U��hԩE/����=�p���'�
1�fMO�w��"�I6
���'&ʴ`Ɛ*�vdxu���V��'l��#���J��DcH�ۺ�B�'{&�#T IHX��C��<�.!��'58�+",�o�����j̃���'�8��E�0�d9�`��|X����'i�p����rR��� ��^��Q��':��e�����g��DͰ�'�ĵ��hU�~K��h�1	��B�'C��yGO�T��`8t�M+L���'�ѣ�'�%9  dFߏA����')�l1�!�-��`���T�5E���'?�͓dj@�  �`C���B*=��'�P��%Y856"8A�I�M@�PI�'V��p�ɀ�6��0WS�V���'�"a�`��&L���2��%G�!��'VRM��I>j���̮5P4@��'4�! �FK��}����0eT�A�'&�h�UBξNS�55/`%
���'��!�qH��9KZ�J�cJ�W�2�
�'�6�0�#^��L���O\VT�
��� ��cCcbĽ���G,x��P�"O��h%)\��1��/��׶�r�"O<�7�݌A{�yA�-��`��b�"Ope��j�4MɌ�������]�D"O��� �P�F�dyƤN�ZxF�Â"O-BP�˲J�]K���Wb�sU"O	)��׺tQ���'BT�X�"O���`&�^^B�	UM�b4Ҁ[�"O�L��EH6s����$�B�X���"O���O�(58���Hó"8Йr"O�!��Ǌ'����fδF�v,��"OΈ�,�b�xI�%�;
5��[a"Oa�N<B�,K��K8���#"O
�Q%��?F����PD��-7R���"OXF�07�F�q�̇=+�AIa"O���Ca��`W���\�(�xH�6"Op�1cb�P/,L�#D/\Hd��F"O���() �ES�KA�Y��"O�e;�-=Öa�g�D'�@k "O�����L��Z���+2F01"O�\�����0+������"O�8�$HU$oB��Ʒ �P`P"O\SC�ļL{�IɃ#��lE�"O��(e�6s���;R���?�z�ء"O��)C�P�@ ��*:z��i"O�7$W �-kDm@�*̢\�s"O��A������𷥀��p	��"O�S�oB�B�*5ʷ�C3G(�КQ"O��ӎA�Qd��EUd�X9�"O
m�S��#��-36m�2T��"O�(:�F�|Ḥ�#c�"aq"Oh�[UˮV&�9EA'p�Z��"O̽Q�
�B�%���'Z���"O����gY [!T�ul��.<��B"Od0U��~����J�=�R"O�-�� '!�����FĻX�#F"OtU�!iL�E���`'�@�V�,8��"O�4��gT���ԑP$M2��w"O�D���P[ԣ��`���"O����U3��V�A�Zְ�(�"O�;��L3$���.Z���"O��S�/��5����tH�J��l��"OH]�5n��o��T�
�����G"O���@��)��0;$�y��p2P"ObLKQ	Q�KM����E�<X��q:�"O�]X�#�7~0R%��YS�VԒ4"O���h�'[��[eb�����"Od� %C��L��X�G�J��"O@Q9NX�A~���W�Z}��"O4���cG�.h���Ro�*b8T"O�!�Ѡ�"$�� �&��8�ʽ{ "Or��Tĕ�1:Hyr!
�tr�AZ�"O8Q�S�A6rXT� Fgٶ�4��$"O,�㤉Ѝx���J$`@im�� $"O$K��u�d%���[�w�X�`�"O|Q
ʜ�v�jq�� �`�d�j"O���
��� �GEԤr�R��5"ON��$�a�rx���T=@�X�"O��K�� �@�`���9�̕)�"O�p�R H��=�s��c(�`37"OV�q��[�Z�f� p+�(C"�Ċ#"OR����Tw�zA�
G%I�,���"Ob|�q�ɳ~'r�K��/��!k""O>(K��"{ "�LO3G`�� "O� �1�e�8n�aPƞ:L����"OP{��I�=%�Ʃ��\�|H4"O
t�P�O�;�M*A	E{C�h��"O��C��	?��`Y�!M@t��q"O�H�d���RmC5��;x�cW"O���`�-,�t����n:��څ"O*��傛�dZ>0���
��	�"O.HIB��TW�,�Wf^�F� <R��'��IC���xt@;�x�c�ҙ_לC�;���kJ]�m<AR,���=9
ç	&𙕌P�����U@��8q|]�ȓ�,|���Z�����Cxt)�ȓ
}"�Q�Ok>��3�@�B�5��K�tZ���P�SFB�;���%�s2��.4���ڂn�}"&]�ȓ1|��%�
�Px��vIX<�D���}X�pI�W�v�lJ!��6 
ȹ��8���Cf��
W�i֤ݯLr�@�ȓ/8�aEOI�%��YCB׫B9J����i�j��i��}��A¶�ȓ����]�Y� ać@�)��_g�(�%4	�90D+G����ȓ	~��r��Ld0w�����o�^��VN@h�Je��Gί~ZH��)\���E=�Xq���j(��CH�1�&ށ+�
�p�$��mk��ȓNm~aԸZ�v�<Ga��ȓ��)1�^�H8�]�&��9#����Q(-	"���3�P��ǸK���ȓ,8�e����i�0�$;|gv��E�jl� ic>T��!E��ȓ'�h\H�1�h���
��\�� ��w��l��-;O����[�URU��"кx�&DM�dz�4�f�[hF���P����E�p���C��w�P�ȓd�Q�4c81j� �;U�pȄ�H8�s� ��-sba���5Ԇ�(.�As`N�,i��I��ðKW�̆�Z
�a@凊y2�]�w�F)g)jĆ�<�L%��X�_v@�*�:r��܅ȓ��u�#kץc����T�� O��݇ȓMz���j�'��(����5{�	��I�%��BO��`Ǒ"��$�ȓc!�2����<���FѶ&
"�ȓV �8J��ޣK��؀��Έ�zL�ʓ3d(L[�� �1,��sD.l��B�,T��s��ְh)�=+��!8*B��6>��D�ƦL9�!���Z�fB�	>9�+�戥Q�p��gB�	%c;HA�%X�Ь�
3:J�C�Ɉ$� @e.��Ӣ�#D�ԡ}�C䉛 .�aC?ƀ��&�^�HC�	%W�4���D�1#@b*�^e *C�I�Ge4�H��7c|$�	�7C[RC䉫HE�bL�=) |��իg��C�ɢ za�Q�)�p9q��6��C��57O�I�AJ�q�B�2��&�PC�I�x�>�#U��:��X�$���w?PC�ɒ V�IQM!m@�Z�	��y�0C�ɦ%34t���'$�P���B�x6�B�	1��j�GT��R�B�F>�C�	�2�68����!J�q��m��C�/F#����K+$wBa#v����C�	�\G.�F U8B(�;?c�C�)� lx���k_p�h%(��aPfśQ"O���� ��t�0Q�5q$"O���W!ЬF��Ԉ����0���"O�(���+_ͺl��CD�f6���"Ozщ�C�%��$���(H] x�"O�"�#YN9�Ԡ����ċ�"O�xYC�	n" �����M���T"OzI1/Ĺ#�ܹx�K�>j�I�"O,�҅C�<&��x�q�ď S6�P�"O�2g�)��3�ۉ9ZD g"O�%�
�'$U�"Ļ>/�1�"O�:p(�r�J���Y0h��"O�rǬ�b�l�!���*b�D�+T"OHp�C% ���aF+_ƞah�"O�p0�!]5h�چ�2�.�F"O��ن��~Y��;+�F3�	y�"Ox�z��:O`b�YT��Hb�#�"O6T��/Q%}�K���.'�|y2"O��� i[&
R���[�2X�V"O�pi��	3Y<��uB�9
k
�@"O�p
G���Eو�q�Җ>c�ES�"O� ����F��ɑ��<!f>u��"O�|).��xyv�2!I���8$"O8̢!��z.�P cꀊy[\�D"O����]�!S���1)�^U�D��*O��5�H�9V�������|��'P�JaCY�~阩��*��5�5��'�I���D�)�Vyz���E����'{���%��r28�HR��;w���'�~��	(������	aI	��'�|(l5���3P*��j�n���'�y���~h1�"ϣjib��
�'���BݓP/��!ei����
�'G�5jq�ex�Ī ���e�<�
�'�Pq��
�}�q�@e/\����'j\j�AQ�K*u�����B+�lc�'��@�ohD�&I\r�y�'���*�]^а����6����'�F���G�2 �=�T⏾?P���O<��I"�S�T�T0�bM�1�H�1tc�1���ȓP��	y�[�&�>X�s�	�E	2��.X�re�����X�B�l�N)E{�Oʜq�afN����(����ȓh0�!����0���H�Q�g}�`��G7�5`%��y���p�*�Z�6��Pfp� �)�7�^� QbHz}��E|Ү�|�O��#j��!�Vlb��D�qc����'�~� ��Ct��hBkK�a�(��'|ў"~z��P�>��m#�C��.�@ć�_�'g�In�O�ɑ�i�?B�9��G�"L=h�y�'��:�Ƃ%~���k���)Q.X
�'?�E�ଏ2`�Uk�솎{u#	�'рu�`�`��Ca�ܛ ����O������=� C���]��_�w��s���i؟0Γ�>d���
zgD�(GKu�d4Y�'���z�"��yzf�+ suh��dѳ�h�ȴك��%�2!�@��F���s�"O��k�+^3iԡ�RN=Id�c��'��:c6M���ٗ������
~Z�ȓ_�T�¦�J[�9��
�<�I<	a�+lO4�i0�I W���+� �4,�)4�'��O���!-�~�<��N؀�,8�"O�P�c�*[�ZbrY2:0x��*��>iY$*�/0�jiK����zc +D�� ~좁�@;(���kBi���e3��>i��f-xԧ_�4M�
v�� �d���@}� ʷKF&�j3/u6�IS(F��:ub��	6��9ᩏ4YXjӪ�48�!�D
]�E��(S�)D�&�!���6h��g��,枅�2�l�!�>m�"%ȷ��͆a����'wʲC�IM�� T� �`��0m�:urx��%���aJ��X�W<:�a�#b�]ab���<�1KE	��%���01�^�3!
k̓�hO1�(�b���V�K@�_����E;ʈOڢ���Z%H�p��ʕ�A�XL�IM��0=���ty�x�OȃB��ӱN�H���0=�	%
)�#Kѿ@��� E`h<�F�Hu{��Rv$��oJ�1SÏ��y2YeVZ��t-N�h�:��2���<��$�+Zh-��_�"
��d� �!�J�喤�R��9��[D��!��'Pў�>5i7��	�lx�����n)��o�����RDb�)�-ˇ
�����o�k��⟈��N� �q�+Z�I�r ��Y*�ʓA����䴟<a+�=��8����"4�(D��)t F�^¬�;���M��I���O�~�j�^�8��M�<J���YG��d��g�'��O8�9r��&*�,]E�ҏ�(�&�x�)��F��H5cRyt��:Ŏ��E��7�'�S��M�B
l��P���-�$UC�IGt8�'������^��t�¯pB�u#R��>�O<��H�B%�	��Q��!�d�+G1�Dx�6�S�DB �s�.�!&-&p6�`+�E&$B�I��,Q�6��a�Uə<4Q"�PS�)��<���M`!RS�����BW��h��hO1�f�0��L�D3v RfF��	��a"OZ0���'<Yc5R=G���$S��O�ҧ�g~R��6��}{��A�e��xh#���y��1��SDN��B�â)��g Z�)�{r�i��t������|s������
�����5+���o�h&���"�B;�x��I np ��eX�=�,��A)Q�㞘�'��?U��U�i*���%tt�;Ǡ݇�y��V�O�p1� ǀ7�9r�4�(O
���C�V89�K��L�c���>�z���ka,H�v�F�=;� � A��O^ �w���d9"t:&JĞ`.v�G~��S,x:���i �t@2?����{��O2�P%�����f���Ae��h� ��y����Iaw"�ep��ش!�!kpH)� .D�d�v���`�ը�(U����+��hO��+<��)��+��sf��	D��B��cD5��*�FeP8�T�

c���y�t�=�7��
'���V8���sEI�<$�={R�]����?1��A�@��A�<9��n�����#�F��y{G�A�<Q��۪~��z���!n"�:#�^y�<�D�#6��ׄ6.� �2�&�r�<��V�3�`�ѥ��%����G�q�<�t�Ӿ6بgƗ;�0#�f~�'5xm�S2����	:{��s�|�<)�M�k�̩Sc��jb��Z�Cu��$�>��#��e�`�	�唼m ^"�	JF�'t�?i۠�g���c���F՚��p�<�1O���(������ �e���3�E�e�Y��'kў���'�x\AI��(U�D�P������*,O��W�YÄ�IN{��[v�i�J�Kش��'oў� Ƙ9�`X8N5\$���9��p3O
��I6��.� 1��1Y$�O�L�dj�¢<ى�A;4��t�\2S������D>~ !��.��xp��7C��jƫ�f����o�
#<E�`@$Y���cB �"[�*�̑��y��ø F 8(�S�������'|b,��ɨ^xX����B="�KC�g?<��>�$<ވ)E &fZ�҅#��#pt�O�m�S.K�5�^� �i��{%���v��O�<����c���  ���lU���K�����dʲ{t ���UM���y��_)U����>	�5{R��I�}�:��7�K7��}��)
���ǿcA�Aء�A2�"لȓ&��BKޣG��CU,X1y�ڵ�ȓJ�H8�g(��	���B��_1��Ն��Ti��b*bZ�q��Ȫ$":5��i�$EW��(US���7��<O�2����<)��;Q������b:��@b`B��4G�����_��h�v/T�j�\�?���	D!|f�����I��a
 #.!�D.U����A�q-r����[u!���4�.Ej �J+j+�A�Ū�Ku!�:	 �	�㚐}�~ 1ǊO$ _���>���]�3�:���$�;�F<j'�S�<)��M�H/�)
�B6�j���L�<� ���a�`���Q3�EӵeZI�<��P�2_&�I�k���L}Hc��|�<�D,s+�h��X���^u�<��䅯e�����,��H�+��h�<�PMD!u�ٛ�� �s��U�g�<٤�G1A� �K�vЈ��Oa�<"-G��P�`¤֣u}�ظ1[�<�v�]s��uC�utARb_L�<!t�͢�.��$kH� �A_L�<��c��NKf��#���&x-03�J�<Y�gA�P#N����'9aXG�D{�<1UK��CLLxrG��t�ۀ��x�<a5�[�'��iQ�86�뵣Dv�<i� D��9�s�P;C�څ`�q�<���i�����P[�|2a'�k�<A�W<<�%3h=����wM@c�<q�Dس>⪡0��H<E�MP��Ew�<�5�ͪ.��@A'���K��!��BAs�<i �W�=�z���T�sh���Wn�<���/]�>$V��l�~X�S��c�<iE�ʪ'.E"�f֬C΂�y,�a�<�3dI*+�L� �m�%>� ���D�<9V  j'���r��=� �3�d�<!�#؉bN��y7��}�H�˴'�c�<A��Ȇw4|���eF�G@&���E�[�<Ar��l�,Ip���wur�qpDTZ�<�҉Y�@���i-@�b�Q1p��T�<���*�ؤ �' 8h	����
S�<I�O�1*Č�g&�$���"l�R�<qnغ!Y�!S�G.L<@A���Q�<)��hc��`ת~�t�EGO�</A]��a���*
�dG
L�<A�̜^%B��ŝ�J
j,��`�<�S���)"���%���m��K�_�<)%/W�	?"�S���
}6��d�r�<I��J�z�b5�C���@Lu�o�<�@T�(�V��� V'��z�q�<��-��U�P��&����P	Xr�<�qF �`z��Q�"; ^4���u�<� D !�'\?2p�Ҡd�1�q"%"O%���"�B����?�\!�"O��S���lv*�����dvtQ;�"OdY���ݕ8���2�P�C�F�"Ox0٦@�*��:�E
�c���"O4l��-\P�������1tRD!��H�n_<�X����\���i���P^���%� `�ui�1���s)��L36��7#ߗT\���%�4y�Ĥ�ȓ+� ��t�ϟ?g�5҇"��!��d��#F��Ԉ�&52�!�3ax��Æ<�' #��1��c+ tԅȓpnDX	�Ꮈc��hc�hT��>����4X�V*�D��b6��w{�|�ȓ.�8�K4M�,G�Ƒ
�M��܄�=�	I4ƛZ|���BSP*P�ȓM�8���CZ�[�����^�s�$��ȓ?.x����2%�*�H o+���ȓ�e�`k�>hi�U��j�@ƚ<���
�E��4
�	���0Β0��}��*sB�T�M�c��,W�¤��U�$ ��Ϗ!Lf�ɂ#�3$ľP�ȓ>�:�(ҬҏiQ�m��/F�P3\�ȓP�~��r���^ �@2��s$ a��/������[7m����U+X�^���ȓW�Q�4b��Aܚј��M�`i�ȓ(���^�5p��p���:vw����l<��1,f�(tc��I:
��P �Ih�C�?:�z(��H �%�\��'�AK�&)������X��b���ٖ R��Zv|#�̜�1����ȓwc2���b�@1CB�)F�`)��?�ܼRѪ�2�^���U*0a ��v^��e �8[�}�# �@�,�ȓ/���W�ξ9��A�i�-�чȓo�"ԙa��>�$;@I�KbȈ�ȓl�,�W	g�8#���Q��$��;�  d-�E�!E�D�$`�y��H��n@�U�4�a��Y�0x �ȓ)ʆM8dn2�ň�1)Z��S����Oа�dYy��I�&ЦD�ȓE1�R�M�i-��@D�c�Rp��'���I�@$L��q�!j�_�D���'�R@XS救N,8tC��
?U~��A�'�.`�`��"	VeY�'ɃW�~,r�'X��hԈ	WZ�Tcr����2�'l<���i�d���1kI�C����'#J�S���^e� �>���'y�0��D�J�2xh�g^"4�qi�KBL|��#�)�K:�4�AC��j��;�!�
!L�h��'��<�0%�$f0J�i�&$�M��O$9��:�2��d��X��sd�h�͒q�N�j�|"��9�,��hV�X�'�݅f:&����� �ΐ�ȓ��9���%e��9ˣ`#W(B%Gy��Գ����`�e�O�L�0fc
�;Ɯ��G9����'@��
��1;�a� 
�9-2��+s��(�cp]ӧ��� ���Q1u�یJ��0[F�;�y��@�3L*	cħ��E�H)�	��~r��";1��7��v����ፘ�M���8�
[3w��%P�O,�Oرs7��<7�rl3fd�&2�F]� nƆ`��� ���y�%�*x_����/ϕ
qT o.�(O"�:5�)~U�����ņ_�Zd�؊A�04���?\�!�$H�`[ y ���r�z�9� H����"�E��:���>E��S˾52@�Q;h�Qˋ5mr4��0O 97 F0/����钨K��4�� 4�y(�Ŕ.M�@��� P���<�<l�	ѸY���+3�'�b�2OW-F�*]�{�
}��� {yb����U|�<��i��
>O�-HЅ�+p�԰�-ҥXf��ɨq�0���Ux�'k	`y3��_
��3&���45��x��즵�С��V>�����9*F��	+~�x��Î�r`�%�'}Ҋ�qF�A�K�_�J�r0��!�DÀz��l�OQ
_�r�0�����<G/lŚe�<A�S�Ox�����x���k�aM4��
�'B�a`No��=cƧ��Drrd1}�,�?ع`����{£���rbL�6}pW���?�C��ʁ� m��+K� ZC�ɰ �:�2��+Z�q�^���3���$�џ`��V1|�F,[��4�ޞ����`FX3gul1�h���y�Nͻe�� XG#��]�L��p��0��$]_�n]S�/�,��)�'<��থ�9P�r�Z!Ί ,6i�ȓ�d�B�I![8	l̀ ��,+��Ь[�f09t�i �HЀ�`"�ϸ'w�jm3�*� �Z�9(����
s�:��ؕ	>p�q����}�ԥ�&@��}��CW%�0��o=lOʠk��J3��+í��}��L�1O�\!k�9��'_�@C�и1����GK
5I��c�E�f���R�L�;!�D!��A�8!��ئi�y
��w�������M��I�ZN�7��u��,R�0�4�C��:��hAȟ�0��΃5�vxA��Q��[��'�0p;Ǥ����H��̎i���AE�zO�q3`�]6�����N͏V�V�	>o轻��L>���8���ҥ@�:w� �'�Ts�'���稍�VLH	�"$�Lb�j��#��!�00�l�<1K6z�!rL#\O����憡X�R yFKu�vY�c�i���`�KP	%��`�O�OX8�CtK�&���C$A"9�$����,���R���yҩ�'F,�	2�O��0������� ~��H�%Au�x̺��!��'��S�;�j�ԉ�?��c�z�Z�����(����Ї*�J|R@�^[{�b��N9��`��D�c�m��G,}b�s��H� Օ�:�1VN�G�Py�.�Iqx�0�ˊ{��?	�!���'3�,��&ϛj�6�K���8��ő7}�P��1p��6�`��|���PF$>7-6Cڈ bW��)�S�BK��t�'|EXEj�2���Hкb�xI��'�N�!�->ɞ8�ޥd�4ͩ+O�,[��F9z������=�y��{7�{��Ƚ-Oa~b�^�&7*��V����̟�ZJ���a�9�y���<:54y"'�ۋP��@�À�yH�Ё�_��4@�9�yb@U�p��	���]2J��Y�����'�I$��jy2l
w�,9$?A!gc������F+Q0�>D�!�#D�$С�Ư��FF<Bz�C
xj�I53f��#XbU�	c�O�taf�$`�\Z�H�v�d˶�'�!0���L?i$&7}�L A�H�9���%�7k "�@�'O����Ď�Wle�f�����O��h�G�~��X�bB٥Jt����R'0�i0g���4�C�>�p�OSz,��^1c�J81bH��['<t�QM�#E�=s�.S������=W��h6ϔZjJP7�B���c��'�F��e&�q�.���U��Xc��U�XhJ@gIb�ڀ�p����nW�|0�k�#D�PCU��5�p8&n^�04B��6S��|�@	 c��ur���30�Xc5�N���O>#�O"J��O�Z'��S�GC :�{��'x޵Y#�"�ֵ��}��T)s�V�c������U�2���(ϖ4[~y��'�0�	e���~��dE}�D�k�XXf�.A���"��'C��d�H�$�	�g����d\0I(���Oo���Öc+w	T	�҉�:*j��ر�X8h?>��ɰ*�<���&�L8��ʆ���`�����&F7ў$��o��j�<$ ��'jf`Ac	�����Ӄa������6О,〯�-n�"��&o�!� )�DF� � �{�Mߪi�T���&��i۟'�(�C��'Mxbr��:t{�!�拒�`�UR�$ $R�k�g\l�$�3� ��L|rb����ߴ]������� g��H�g$� ��N�'�,�q�A"D@�;O1fJ��?1B4�ȣ�z�a���D����͘ �4� kRb�(8�OE:^/܄9�'�~��O�p��'��A��#
�41�	X�_�2���_g�%��@�O����S����)^#
� �)�?�̻w��U`�T�#8(X1ǜ);$�h/O~�� ��u��,���?#<���(|q�0&)4d�ۇ�߆p�]��kx�Z��<J�e�S�?��&�(6�._}ޑ��лC�Z(9��-=��ș��P����%,O�ɩ��\�Z# 8:�4�"I���)|I���F�Rִa�,҅;X��҇�i��pc�K�2�Q⠧�W��,��]�(X6�����DAO�w Э���ws��8��.�"���a�i$ڕp�.?���q��6�� *�q�h�5A̋�UՐa%ԌY1�\p˨(jU`�<As��vO��|JE�&9�z�Bڲr���u��V#��R� 5+�vnVR�����
�65Nx�s4Ƅ�`�d=@��Z��J�X	%���[$9�j�CGi�yx��'�ป���$:t�q�ɟ�����Ћu��Jӣׯ"~����M�@��"32b�Z"G ;.nN�����w��)Sc׮�u�K�M�h�)�Ĉ�ɘ���-C3I� �����'��9sC�Ւ	��n�6V��q�D�a��1bU�V|�x�`%��cs\�
!f�.%F�;e��P��F)��'Q�Ͱ�Dޡ`\�tȥ/M�_� uՄ$�n����1�	<�?���ߘt��)�F�		T�Ћ/�2n�T1�dI�7����P��,;�1�H�K��5X���Z����Y�_�>M�@��d���Zfm�.x�����s��j��̬`��7��z��d	�&��"kX�F���b�#D:+��+s��T����*�yB�WvGĠ���̓����v'�yCpiQ'L�|�0����l|����V�uAά��P>��s�~މ���	�it���Є�����>D�@j���>غ�� �9A&\5�%��&@�hՋA-���$bՂ\;�Ab���ݲ��Xw��'l6A��Kc�^�ǑBf�0�2B�0�c��O�`����1`h�"ɉR����&ޟH�������%)/��x����rm����
<'����h�1���S�eY!2�axR��E���D�](������o�9���\�$�'"�/-% H!�O<:��;��}��� ~L��A����!:E�� Yr#BM�P��p��p�����BA�rP�S�/��s����ȓm����M߂~�r��"�Ǩe�0\�ϋ#M����W�/Qv�j,BG�'��-�c��~�,S\�-���-�+`�0��	$-YS��=�̴�ЭP���EۂI�)_���<��φE�`�[���u�)A��X{8�P���ͥE�ĕ�$�a��嫁O�/��2 �J�H�m��y�'єܹ6��v���a��
���H��k�C�,7 P1�![�8�.=���S+'��L�!��(+|�������C�ɫs� вaC�@�t����Kp����,3|M��'�
�T�8�3�dSk�Rj��	O �,�0�^�!��Z�[�$	z��'V��W��%3�|͢���!�Fe:�ᕋ�\��Ċ4	�T��w� Dt���<��yb���E|�GM�1=��Lo�!__����h�ǠDa��=`&�B�	T<%��@=�Hi��hQ
l���\s�H�6t��:��ӝ0.�|B!��$����
7�C�	=V9��i�|����ƚ9�x�[!A���'��>�I��(�)�K2?�8m�A�T6C�(%�^ݨ5�"^I��P��ζC�~B�ɻW-,lib��^�zx;�/̯:3,B�ɐv�)�����C��� �ύ�"ǤC����?<���r�Y�>G�B�	�6��mJ`gU��1
���1%�B�ɢG^y	�ǜ�a/����O�1e�B�	�	��B���;1��:RC�;T�B��*J�@�R��uH���I�jB�I -��p�$,�'"NpxF+�/�ZB�ɷq�0;e'RS"@R��+B�ɩ�H��.X*2�0�ئ�	 r��C�I�3o� �3M���h�!�%m�C�	�X��#�eZ�uK�'��czC�I�I'�Q2ʼ�@Yj5+A�WDC��>cy�
�0�lu��2C�Iu�0������*��s.^�Nb>C�	�I9r=C�R��H���\�2C�	?m�m��B����0��]�U�C�	:5 %eՆ1n�4��ƵAn�C�	��24C � 9��3�"�?�NB䉎UŸ�d�H����P'ֶU]B�ɠ��ѫ��K�N��Pkr�"y�C�ɗ� ��&���`��-�C䉲>�Y�"�&���!g�
Sr�B䉿i�� ���^�iL۴��/!�B�I�59���0��R8ND����Q��B��>}�� !.��3�p�+�KEjC䉕?'^�rdl�P
�m 0M��bO C�IX\��	`�R�|D�MP�D�V�C�)� ��!Vo��R� 'K�%��a"O�b�O�_�xt`A���-c`"OZ���oɝ4�Y��S�aD�P{�"OT��d�M�:�ЩѢK�5yO��(f"O��Q�A��@���T�H�z<w"O����y1!�+y��U�u"OT��-�g���h�-�6Ts���"O(k'ÑV3�]���5Xe0�"Oj@�wǈ�+F��Q�,���"O((v	3`Yl�PQe�26�&="O��ʗ_�Y2u�UaS�6�H�+�"O�)B�+������Q7���Ia"O��ڋE,��׮�Fܼ`�"OMk�:{��p�̕' (ް��"Ote9��<h�<%8�,O�?��yy`"O����I�(~QI�!/l�"O$)��4������^b�"O�t�4�Q8m��$)fkC�vt+�"O�5�����.@�u��*~!R��G"O{V��p:2��`�L8�9q�"O~�(R��5@X�P�� ��"O�qB�$w-�	ه�F�;	�D
w"O�����<���e�Φe��+t"O|�R��ڙ,5�(���N(9Kޘ��"O���ȠL�-*���$&�`�"Oh9 C$F��@��Ȍy+�yq"O.�#�oM�Pacg#�"Hv�\8F"O*h�SI[��B�[wE]_��v"O����KJȸ�CE���`�V"O@!�B�]�Hd��m�F�."O��Ӌ�/� {˗���#�"O�j3�	]�h��UlJ�@��*v"O��3��E�H5h��V+y��@�"O�U)rN���"δN!��Xe"O  C셲����	"t,2�"O�<	Ј��̢E��M����"O�X*m�m�ڥ�{�T��"Ot�u՟)B�Ļ��D�I�
M�%"O�x�����~����Û>�Da��"O���g�{�	��7o��%a"O2��锪.1�S�Z�hs�Ӵ"O0�A��ԝn2}k��o�0�"Ot�˥M�;����ƃH�5�b"OLA��f��u �=?7|YS$"O�	�eF̴1���bH�*� �&"O��B�M	�U�H�y��}��`�'"Ox5���W1�,8�vf.8�ɳ"O��@&"Q"$=sc�3<r2L�"O8,r��cmAFi��j�#�"O�-���, ���F��}�$���"O꤫��U+'U" %ժ.�-P"O�!#��t�FBP�_k��*�k� �?aCJ��`&�"~jc9.^�2lI�H�$4�W�ޛ�y�HH�(���c&bQ�6�Ip�[����3���(�I/\O���%ٽS2	q!��:����'9R��t
B�o�h9����qﶔz��6@x�F�	x�<���L�ܑ�ē%�앱+�z�'���Ӱ�\H���E�D�$A�b���+Xq��A�Py2�J�F��!)�2�x-����
wq��@�Ÿ��O?�$�#
9RH���|����g�A�!�d	�;��Uk#[��03V�������Ң��D`ٰ�0=F����Jʤ�A#i���C�F_8��I2�&q��Z���M�P��G�E�Is��GN�s�!���k[��a��Uh��؂g��k�Q� ��lW��A�3� |e�$�_�p��S�+�;x|]!0"O ���*S">Hy��V�zz,��B@-~�&!�U6n��S��?�㌭z)2S���2g\ب	��G{�<�u�Y�JW�$�L�$��Ց�[?�r��a�� ��.LO��P��/�j�Viʉ{5�'`�Wt<qA0!�fh�I��1fɃ�%_ܓ3��I�2�/O:�:g'���*a2w�Bt�0�`�I2z��SJ�'��͡��Q�&�`�{���;k���sL�x�]b
��5�90�aճU�D�0���>�5��bR5Ke��C+d� ��A=}��2sf`ؒ�.D+�P�� G!�$H�|<��"�һC�����>��	 I����@��S�OQp�IBF
��|�#h�$e����':*�[d�M,3<-s3c��Z�����2}��7b��{����{�].oU<����{��h�$k���?q���,i���1F(��:uVՂFˁj�1�˛�`�����O̲�;�M�(�ZU��8)yџ8�r���ْ
�E�S,z��pp��t�\X���9�C�i���޺6Vfi�m�v�R��<Ia��O���U%}���C8L�Nl��O��h���!:�!�WZ�XL��$S *���Q�͸Q�z���EmM07͛>?@:�y�j>���&^P��2���%@ƶyj��Z$7
��@�'ZZ��J�Q������0@]޼�友���!��L9YJ���;8�P ��� ���I���		����q�$ɉ������� -�����:9�lSrlT�v7� K�B��:��g>D����(�+���r�-��M��E�ჿ<��
Q��i�EoB��}��Ô|XR)�F�ħ]��Ӈ9|�ɵ�X�Z8����+T���䋴:P�H����r#N����<��Ey��12���3gԩ(t8@�|�r5#f�ؘ{�1��'4lt�N86|�da����Qkj�k���_��$�����O�h�����X ���[���P��'jb��A�ø9�����	>1,���+^Y�i���q}�6�E�:�x�+�k�!��)�	�>n����#��x"��G��!jv,ʱ��]Y.��Q"OTđ`��I��1X��̢)`�h #Q�DZD���hQ)�ƃ �`BP��d�d�|��CN�y�����^�\��%�BX��P��>ql�!ӥ~&l���#��(��+ݕ^��"<vh�O��}ΓXW�H8�k�Sc�ceM���Gzbޭ/E04�U�Gi�'1v$0�\�3�H��e��N<}�`�2������=Qg�<�Dp�bb�)LZ��p4B��}r��Q�]@x)��>�|z�Q	�����gy�Ŋ�+#d�!�B��!�$Ĭ1)�\��g
���A����5"剟(L��F��^����`A��V��dH.t���k�"�O�=�aAE����Af�
%��� �)l�p�k"O�Iy#$��Z,8�§5V���"OP��G��wh$��[�x>Y��"O�h��
�&c�6�[���nty�lpq,O�Y�d.��Kʵ�ī��pI�J�/P����R�F�bL �������J� I	�-Tl?)�@�f��T�T�*�ӑK��I�y<���݈}�:��DN�:r����$�?���P�'x8�:�@O����� �� j�Z�	�Xq�Y�Lraց='�J��O � ��Q&w�(��?r���4�䟹_�M:&e�8�s���xj���OZ���
T#6���֏S�Yf�A�U͂*�T"K�n�����E�8�0	!b�?����L�i_����'d�}�c�}�̀���$9A��ڗ=�� �Wjl��	3������sK"��T��?D�"�䏱y����H�����<�)C"�Y�_x�HF	L\05���'w������d��~�mL�s�R��ū�����
�0=������A�L�Oމ#&@��;K�}��I�2xI.�g&b���ğ��?��{J�I��(�M1�u�4��\����v��u&�|�<�&&Ms)�T�D��O�=�Ū�,ko��@��L5�U��Ì�'�����B�&Uk��X�	�~6ؘJҏ�O�`B��Z�t����DɪH�`Y� ��R�8Y���&,W���D���?!�*4kE˗��Ea�?AD��D�C&��dy�Ҧwo�tk�6����F� w%T}Q��Q������	T^�d�>(
�t�!I�ul^�¥O�.b�2 ϵ	��Z�FU�^�TY�r �)�@���/vn\��>TW����
�`ڬnB�����C��M���Q�'Pf��.��X�"a�U�Fe��?I�E�W�z���HA=g�>�*û~�b���]�6��������џ���^>�:�[��1�G�4ZE�\��T&"Yظ�gi�~�T�5$K��?)��
{���9��ZG�H�RfԦ���<��8���Y�K�9�c�_�ZJh�ɶ��<!��'yEr��Ǜs���� ���`���cA��X�T���H
 4y�d
S�lr%�ω?��D!�O��n��"O"*%(l���M$`�~�8�,�7f�Xu���"_��P�n��$�V#F�7�Q�C_���r�1/�
܊w닣/��8�[�.�oځY�~U!TY���P�僸gY��'�xڲ_7>��rT挈 �p"�����'��쨢��k{L�o�2'p�%H^����Ρ6ND��#P6-.P�UFd-
#��9M�B"X=�'|�D���T�]U��!`�*�EP�h�Ny
a5�V9r�۴	�MjbiΣ����Et���Hq>λ+ �@�aP8^l�XK G�<@-�*Oz�9���:��9��?#<	4�كu��a���4`6�B����F/�@w+�Hp�q���R�hp�S�w��I�Tǟ5b�N� ��@��S;7D���󬃏3��-�(��l�0�cS�'��9�w�B�o�4�oژQ�+���G�z��2㍵qz� �9E2��Yĭ׈/5�p���VS�CÜ�D��'qSÆC�Hh�шI�8��8���4��������?��C��6}�I��٩nh҈�� �R�`�,^�3ǎ`�CƐx<�	(&�Of0�/ۘ ��hv�Q�}@}��mF�k�`:O��PGU%.�j �^wb�*6 وG�����j��Ac*��B@�@nZ��"O�8��O<GDP�"���J~�1�6OH"��{��.�T���l�>�'m�a塟�P�-��ΕE/(�K�'�t#a-E"�ӦD�a���&A�7��qB �OVt�%�K� �.0���9��T� �'��3�TYyR�Ѓ%�z����_�)	d��O��y��-m�&t���ԁ '2 !��^&�y2g���IARO��sݺ( P� �y򋟳�^���+��1/4��FN�y�E��.{���ũ�9 ���64�y�G�:�|���+���f��/�y�k\�<�t��ծT&E��q(�8�ybj�atuH�O�G�|˅���y�+�}�F�0[�� ��y)��g����&S?aj�aaT,3�yr+�l2��@%F��7d,�C��B�I�'qxL��e۸sT��YC�%� B䉾&�49d�ʯ-.b�����p3ZC�	�WX���&@?nĘ���&�\C�	�4^&����͓!R��3A:�2C�I�onz9٦ID�$��oA���C�Ɋ(,:ms��X�4l0��i͐C䉞!����6�Q>*/,[��C4C��%4�w
�?)jP�
'^�J�<C��X��hW �%D�,���^+�B�ɍ<3,q�t���qf��ʤ'�8
�jC�IтW�Z*x�l@� Ŗ�!^C�ɶy�,RV5g�LH��?H0C�i)�c��x�!�d�$H��"O��)��K�?x�#2 �;e�����"O2��'ē�&*J���˫/�~r5"O���#_E'���E)Y�Mh
h��"OX�B��<[�iM�:'��)�"Oh����e�t�b��L�&$L��"OD �T�N!��\h1̱�4�"O�p��+g��8 hX
x�q�"OL��e����ј7
�h2~a"O4�ɑ�˗]�v4cvI�qH�h�w"O؉��&��S����h!N�*�"OJ��j;���)T'P�b�"OpKc �uH�tJ�nK���A"O -17AD:Sr1lփkt��3"O�	�!��;6��7-h�Τٔ"O�]�g�~��� �ݩ����"O����� �b0DS(�4<Y�"O@ ���++a\�R��Q�0|�"O ����x7����"�J�"O��S�ޡdK����:���f"OX�
e�*զ�I ��y�pt�W"O��X�#)L���(��B�1��"O�Lŏ\��U��M��YKs"O� B��b�V����ǫ[-$�򉊳"O��P�P*	��p5'I,�d[�"Olɩ5Ě(Ԩh�L��[8�p��"O�A1v䆋�$Qc�F##A"Oj����yv�ˢA�prL�'"O�aS�HQ:����+�E-"O�,�2+;q��Q����~7r-Y"O�l�f��t�}X���dE��"OT@�q��I��aJ�%W'=��s�"O�<�����������]!�M��"O0�@�JJ>k�.�y��\�RG0U�"O*���P�d4<t�a�G�1\8Ȗ"O�L�`�X�]�΅S���z�q�"OnX�u�X�E2P�#军�k�)�`"OH���"����)���"r����#�}�q�Z5Q�Zwo�#f�V�?�6��I0��-�=k&e3SN`�<�P
��+��y�R�I�V�YE��Q�<���3ot�)��2���DHd�<Q6��u��Hr�}�L�Z��A]�<�#RCl@ G�)+t~�S�V�<����Qj6�q���������K�<Ae�W�\?�i�G�O+�Z��%�I�<��>0��,��Rh&��p#!�J�<��M��
�x�1�i�>I	f�7�K�<Ag" �i$��h/ۺj���U�J�<�TfȥV�^mg��&Jfm�wnUF�<�!I��9�lÍ^11`$��K�~�<a ۻOa�, �)�RkT��ba}�<�@�~1TTJ�ƃ'Df֜�!�m�<�ԣ˅4��Da� P#"����i�<��*e�T���ޝR�~�#s�Tf؟�nZ�l��c�̀=At�蟆V�@pB��C*xB((�� ��ɱ�Ŭ}u�9E�_�e��[��12
ҾB��qE�D�'��kE�F'q�0d�7��l��Z��T�bd2g�C�~���P��~�֗ff̵# �3>�ҵs�6�`mI&F\: VB!ëO���؂j�4Đ�Z��24-�#��=�F�CE�˓b�\G��'-�`cœ�h��m�#�8B�q�{"�)�����Hh"!ϑ�om�1�HZ�8�!�ڭ��(R�J^�4,�[���!��[�hѸ�;�է"��chƥn�!�D�!��`H�`��}Bd3�76�!�D�$nc&E[�!X�,^�@�b�'Y\�F$W5��l�W̓'o�"�'��8J�#_r!�MW�$&�a��'�����%Q+�z-ꕮ�5���
�':�"p��!��|�e��6�a�	�'؎M��G��
�0�R�
��=�����'�*}x0��(��1����L�]R
�'�ŒDLDC� x���?��	�'6��+�V WUҠ��� F��b	�'���3��W�ZҺ����x2n���'�̌�u*A"J�.u���A�_�F��
�'���	�(Է`��885�	�Q��x:�'S�, ���9 �@�ɁM�C�E�	�'ڢ� ӫ�q� !���G:���	�'S6�$+�N��a�l�E�D s�'����N�U���S�o��r 8�'0�$Jꑯ/���DNI u���'J�i!��I�Rd�!��.��ճ�'H접�5����OF�W>���'�b�cH�C�QM�yK� r�'F�x�Í��T���b���<rƚ�x
�'-Dy��,�0DKHԈ�	U8v88Z
�'=���d^� ��Ȓ� t$H�	��� ����(0����Ф�9�4,8"OTr�G�J�`���ĵz'N�""OHZdF��r��`"�4f���6"O�l�r@�41�1����},��X�"O�
�.F�lׂd�'70��"O�$Ȓ$�!��h�F̋�6O�	I1"OB��O5d�8(���P��""O0=Kf�*9�Հ���#m��j�"ON��� �0��ɓ�f� c�y�&"O�	��.��N@��h�hH	� �C�"Od�8��7-i�i�ק��Y�J��"O�5��Aب���� f#/�t8�"Op��F����MJv$�����"O*tq*%mڨ`vb�&K�Zu� "OjM� ��``P8���Q�ՐD"O삅��=Q��e�F��+�H�"O\	sH�(>9Z�猄	���"O�D���U����Y�D���N�	�"ObmPAjۤ(!��!'�X)B��"OD��WC�(EJ��&I�@/���"O QK6",3���Y��F�(q��[W"O�9���]2����aŻhX����"Onu�E@��fH����J�U�"O�]�� Z!<h�a/T�D�NT4"ON0�Y7|�4L��mB�b�""OPUô��yw��b��1TB�H""O�����%���'*�&��p�"O�h�BG=�UT�� J��,(c"�p�<���X�T�6T� ��h=�!�Yi�<�eg��k��{"�r4D�w��p�<) ,W�.]���v���}:gj k�<����u�:�Y���r��5BB��h�<��B֯I^��R�F>�T�b�<	�,�|�p0���
�*Ű�@�x�<�a׫L`T@�c� ����O�u�<���� ����T�Քa�v)`�r�<iV`�y��D�%��x8n�pNp�<�[�R0s�A�~�ܕ37�m�<�E��<�
���lܿ�,{�o�<��,\&E�̉V�>bT��cMb�<Qҧ�U!��*@�<U�b�j�]�<���� ����-��?� d����W�<)cG��TS0w΋��0d���GT�<�E�s]z5�'���"h��1��Cg�<���Pͤ�� �Ъ:@��7k�x�<��琈<.Ļ�英F��а�Ut�<!����("OW��XF�h�<�H��`�+g�!����M�k�<yE�=>C�Qʧ�"k�:,���Do�<��(_�0H� ��ޠ ��'l�<a�ˑ�.H�A"�	��(�0��B�<��o̔���[���g?dpR�e�<�'�2o툄[�b/7��=��GH�<�C+�C���Z�EVf� @X���x�<Av�h3��8i�?Q&� ���u�<�4�;.���0(�?%9�(��u�<��u����Ɍ9Zܠ�д�i�<a���(�wΑ1F���W�o�<ɕ(λ
,�E�vl��{������m�<�B�k��ܛ�+܅*kn���LYU�<�ef��^z�@qW�@.���h�V�<��bV:�z���5e̼04��{�<��Naؽ�a�	��$l�uGu�<)���XM �Ē�lr�ږ��n�<� ��{WF���XQc��&��=zu"O�*�hˉ;(�Y�Ѝ�.��*d"O��8'�
8< �q�L�;"ƊL"OȽ���h:t!p&�
~V8 �C"O.�h�LA�4�mh�c 48֑��"Of�����@���B��H��"OHE�&�^,ɰ���BJ �Y��"O2`k����xk��R���4u��}8r"OT�*0�5`�C�vex�"OT|�d�ɖF7z�
bOy���"T2�y���>�D��'���;�~���.�yR! B�P*Qn��(�� �6�=�y�e\�(��ٺ�n���ખ+��y2�O��Y���3��c�+W��ybZ�2N�����U�����Um<�y"�ش3�=+b_�Ȩ� ��V)�y��#X��@`$쎩%,-�ӄ�yRD\�V��A祉�44�qF퍼�y���0�]��؉S�0����y��û$��3��ͫ&�=2���yR�� ���5'��!�j�y"D��G��2V�B`����!����y��Q�iU<����*�XCNR
�y2AO'R�.�k&��,���Z�y �	IR�{h&^V�+`G+�y��[�B�9����#W��Z�&O��y�K��	���Y�B����Q�iը�y2��f��(s�諅O�y�o�Y�`��
f��$>�yrA�8�j�@�eD�,k�ͺÂ�6�y�K�l�l��$J[�w�D�"	���y�L����o�>�H�L�0�y��1;)�zp��.c]���!���yb��:�F�Q���0\'\���m[��ybZ%p�PhC�k�TK^iw���yB͟�V��h�/\*]��� �y2'P!��	�ӻ)�ݢ��H��y�%��$8��N���p͟��yZX-ac]��^��O�+}�N���'�Z C�m��`�,�۰d	+a;�y�'x0��M�Ybt$�a� &^�r�
�'�4��ti�/����FW�
��8Y�'��R�����*�z��I	�'J1��7h��'P; $Y��'�ΐH��rޑ��ρA#���	�'&�ˑ�ٛ@��t�u,�"@8�y�'��AyE�S$w�$��`��,����
�'ؤ��(��g�PB�F�#��
�'H��ᦤ�<H@�ad`G+�q�'�$dY�J�4���N�3���
�'�`��R��6L	��\S䜣c(D�H���
�v���.K���@��%D��y7�Ĕ-�`�� ���K��8k�$'D��ӒdC"N	������r�$D�ВG"��?�,0o ]����&!�B�<I1`{\@�y־O��P��KZ�<��煱Q���1���;ȸ�c�,D� 𓍞<�U�`l�[�ԼS3&*D����א'�x�w�^TrpآQ�:D�d�$�O'h�L	�mܾ����9D�����#`�61�����̬蠊8D�|`�@��e���kZ�f�x�s�"D�,Zt�l�$��i��\NN`��I:D��{Aj�/�<{S��G��43&:D�� �1a���o�����-_Q��RT"OT��$bE
N�^�	B�	B52�P'"O ��Q��䣈! &mx�"O~l��K�&��`i�R�#�"OD�)F,O�Qx,)U�\��"O��9�!�}:DK�4A�]�""OѲ3m�gm��s�֝t>�� �"Ot����}Zn�yR���D.���"O�����3i��� I��]�"O4<�]X���~"B�r!B�3!�oi�=3f�fj�H��ف�!��(<5��ɽJ� s�M�R!�d8{M�Ds�L� �y@,ȏ~c!�0s�l��"k7+��8	�C�J_!���)Ll:�jw�I�)��!cE'�cP!�$�"5�౨��.G�a�C� 9!�DJ5}$���17��j�c�:!!�d?�� ��۳9�4�1���`5!�;|�����!�4W���:WC��R!���|�(Li�Ōf�ꬳU�F&Q�!���n>.<#fg�)x��Y��R8�!��+Z)���m: �F|�P��=	�!���8\���͖2un)AѭV/�!�D
�}�ņhT������"�!�D��7!PpK��+@��!�lR�\!�||>}��������vVe!�Hs�z80�߶;��U@K�
>!�$�/L�0�͘��fI�;N.!��v-,5a���!����Y>!��QJh��v��S��hriA�$,!�DE����z�'E��\�PHJ�~z!�dU*1��<]~Ĳ��em!��E�`��PN��<���H�5�!��4Hd���%�[�։0�d�B�!��Y�)DI�(I�P�s"��!�D	�	��uC*�$!��.J�=�!�dɯYb܀cplD���@�2n�rm!�dI!_�U�bk�M��� ���x!��OW��#��&!�|!s�ьzL!��i���1���M���.*A!���EP��CWD �l�~�ٰlŤ",!��,Z�w���Ѫa1b���MJ�<i���E��A�ԁ*��]�NC�<�q�*{��a��,E�p�G���<a���ԌqBDkӄ�S�Of���U�eR|	3���Oi�]�7F ����U�S���O���5��OP��HP�¬�D�2q�"�F��ɝc�2���iZ~����w�BdE���фzm|"�拴{{^h�VI������4�R�'&F���b?�1`E<D��$�ƑT4�%b#H��8�I埔&���e�?����B�yG�Q�$dH.A���E}b�}�����O�	mZc��ɺt�δK+B veRu��1Z��$�<9�	��O���'P�'7�'&l�`�O�cM�H�Bg����'�B$؏mиwB2O�� _<L�l�ãϢ(�b���
EId:%b�G��)-$�+1m4��O'�b�LsFaS�UZ��!#�V!��S c�4w���'0`�0��'nJ?��?��43��=b��ѐv) 0h�&�/Ԝ�1��)��h�/�}NE�ugrˠ��s䷟(شru�f�|�O���Y���O�6r��YC]6�Nd ����vicߴ�?a���?QH>�'�?��D�^�*���bp��K@�X"V���i9�O��z�@�-��L�-�.�@ �
R�J��m ������ԙ=⛶KY�-�ԍ�ՊT���j�_���D\Ȧ��Ipyb�'��)�I�>ԍ�ä&L���+�%��t�!��LZP�K���.g�Mr��\5,��'��&�a�j�R����ir]� ʐD�:r��[E�@��Y�	��䓕?Q�*�4�<Y����B�9б:%���|޼�# M3�ft�L���4`�}�e�?)�w���j~p`�p �WD�3�'7�	��8�	ǟ�;J?� n	���J�I�/N�P�\�+����h�IG�S�O\�X� ���J��� �#�"c-����{"1�b�Ʀ�S���A�ВY��<�A��d$a8�^�����%�M3����Oe��i�R�fN�Lu������\a&=���O�h��A�>����'�2��'�F�����]��l��H�S�p8��O�Ls���!+|���&w��E�t�O�\6f�STf�'��tɌ4��ߢ2M"�'>�7��On#}R���B<�=#G�V�(����'L@X�D�O��=�N<�u�^kh� a��YR�Ui%�Q�'F7m_�I�~2g!Sk���BWIU�0�K� �O?�/OB��i�]������IL�{,v���+_�U�Ƙ04j�9,KD��ޟ��&�=�p=�E�{���[6�W&i䊨!�ӟ`����u��x@Bο��g�g��&�ݬ���3��  -��y�a��$[s�����O�gy��'ɛ�h\��A�q��88��G,�~R�'I�ѫt��8Lq���eB�+|&� �O86��O�O8���O$��M� 晤x4����� o�4:2&�<	P!�DY,7j & �