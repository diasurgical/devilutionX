MPQ�   v�   �� �                   v�     ��     k�     �       p               9       �        @  ÈMc��[�I�μ/���)�z�:b=����Dss                ��µ&) :���0�����8�?�H���k����e��љ|��j|�   1   �{���Xq����ʫ
���.O�X�.CW �< ����V�R����2�<   �  �?   h  Ս  ^�  ��  ��  ��  � � �2 �N 
j A h����;��Àq#3{���&[�.32+Y��l!DFQF��%;doB��̲I�x��:��<�ϯ����j[\I�)��ʗ=��K����4���3�@�A&�R`������'��/�Q��6��u��6�ؼLl���!ti�kd�#�f��M��x�ݭ�=��{���z���K�۾�7N	�����n��9-93~�r:�?�6��DI3���=���1�mT�ҝ'�[Q����t�u��WϚ�5u�(��pȲ*b)��6����#�n�~��|�L}@%�e�A����n���5��쀽�L X=�fZ��:S��P�\���R`����E�<��C�V��@]M1�(� rT4�nc��c�`�0VlX+���K=�C/�d|��{g}S��ܛ;�١J	N�܋4����N{�W���jD�VN�יִ%x�H���}�<��U\0qB0/�55��oz�^�ͳ�I���V%���5`���u �6���v�����Y������!�&+0f���b����������y����Aݹ��N�z̫K�����;��οm�E�c�'t��4ÚU��MS�+Dj�Fâ�S9j?ô�0�=A	i��!�Z��������Nܢ��qW^�τ3_P�=y_���i,Z�����`�Ф�2&�n��	�zh{�GvL7%��퍦��KA��x(M�Z��n�L��)հ+|V�3Q�.���!<�xĺ�3��&~R;�[�~(�-}-_U�@���� �<������	�O��%�^�ef��U�A1��n�k�66��~��2��x׋��9&=��*[g�[o���{Փ���eš6[��ټ�������4�`����+~ǖ���$Fr���<��\q��1����/�7-q#>ֶ�.�)0`Nc�Oi1t��
���K~���}O�bR�Y�v�f��]
1��x�X��$�vo>�P~8��()�e�(�2̺r7�uS��Y)eu�V[�7N���DR���b�H���L��2-�y��vЅ3F���*ш�-m�|y�rMpv^��B1:�#��K����o�wl��$��A1O��	���D~J/�����A1u��!���X��$E:,��B���Y���h�)\�_l�5�OrP=�����X'~_����@�Ջ^�L��!��Cs�O���X%���Y)凜����D���3��Jɍ�b&��r�B8�.��O��:�||��B$��F���|)aB���Xg��?�b}����V�Ҍ���� 3�?�b;όg�Qs��弾P�q��>�1���T���8�X!�~{a��:-�37��-��S�c��a��ۃnw���V��h$��.ޛ����c���Aة��MP�IV����I/�b�<�װ[UљR�ךU�j.߷,~|�a0�4� 6,
�z%��R"�'cZzG��ES����	L���"�说��k�i�i��,nr
)���8Kͨ���)��у��k��CS>`�v���>0�#݁�t�.mސ�#��B<Co�9�U�K�50$�r�[�"��юm�:Idߣ�]���萍���ߏ?��6.����;��ZU-�J P2])���.F��!t�1�] vX/Lg��$�n}�ЮOT�Z���c�R�n{,��3���ԯ���j�.�i}���NF�}�M����l^���8�@n���3�� 0�yVU�#�:n`��4���rKĂ�܆�3?�p�����P�]Pd?�"��Ab�]7�zK�r@!�4�5<�e%㉿�)��� ��N�N�2iq�'-�*#��0m��7��~�㾃FY���a1�whz��ю_�}s��ѯ-��8�گ�)�:�D�80\`i�a�o�Q?]�����6�W����6ֹ��"���-M�[O{ĪB�W��6��h���ɑ��b��~9�f��m�e6�Ѽh2bx �lX	�T`Ƈ����W�4���4�F���_����&����pu���.Q���Q�f���k����	���3|��O��u�רH���o �?���[����"a���AG=vA�=�e�!QJ��28i���)�ui�$Ӛal>f9.���/�$i�׏T\�9���������M��_6E��ü����z!P��!K~��R��M�&�5L�S�;'01��&�������C��e��a̮�ֽ���L6Lg̶��=�[�=�؄��O��C��9e`��b6/�������u����.��B���BԹ�E�?������οv��_Ӡ�5�ኳUL����i��l��Y�*0V`�-�F矬Qμq&�l��u簕Imu�1N`���s�<P2��S��S	���_�{�ٱ��4<v-wX\�&Ϗ!�xZ�|.���kL�:0'��U=��v�90�C�DTޠ]��'��V�l1���{n��
cOx.��p1#�`���׫�^�T�8��K��x0��?Ӭ�<7:��,fT#�d�}���=M�,��q`�PZC����v���霮�ʂA�޷��t��@|(������a����?�~�[�-X���q��/���P�;��ϙ8������[ɛ��,�x�T��� 6}hx�F��t���*8�ˁɏ�sc)��V�o�&���ԙ�g��7:�?��rM�ͬ{�'�}ZC���^kxR�"��9?ꄂ�Qх�7c��{lX١%v���N�LXIE��V`�k�ݳ�{lP̫�#�g�Ӫ�l��F���G�0V�����Yz����߰y�D��)��F�S�������m���F�p��w`b�5"�����0&���Ş��<)�1��)��A��E��>P��+�U>oWC�3^z��}�Ǉ�ݥF֓l����X����f�?k��A�m�0�:D�rh���c�G\�g�IɬX�{�ד%4��Ni���.�g)��O;�_kL�*�,�z�|?���7Z���*�Z8�F���Xo_�W���i�k�A�>I��{��]4�DZ^�P,�T⫢O�eU�<���	�x�X�w���+�*�n�������
Ћe�=[6�2��ϖז'�`5p�A��>�/�P�����E����p��B`�J��:�=�<B1���#��d/(V�w=�ڪh�;	�Tz�K��{�P̓��� ��Y�~�w]�&۟��d���QH�NC>����,3��{c��|��Zg���F���nѡ�c�"A�A�y�jc#���SaN�&��1hL��ӽ�z�RXD�t�z�-)���WHP�2͊y��������+�P��1��l�Y$���5E������'��S�x+.�4�x���i?ΰB�Jќ������e�R5/��1`L��je��g����X}�p�'��1<�c�v�t-�t�A!SRn����.�(f�q�IH����R�P��lt�E{��nYG��J*q���J+f�(F��E����!>*z�͆@������K��6�1�V{�#���)`����o$�1�����z?�ܤڟ�R1-�F�_\1��9LX�iLґ���V�M*����Ǧ9b(�I�*�)��np����M[J��>��}R�UoV�jih�Z�Y� Ţ
f;��:]���I�P���=���tE��\���oׯ]�:�=Q�'�E`}��o��A� �X�;���8���*r�������4����4+=a�</M�|���� �w�Li�r�������G� }��\vg!�x�X:=����p粠�+�C��-��������m�Z��C�t:n�:BV�ge�]�:�]*���Z�B��%`l��`��;���s���=Y!¾f�zPL�PD�j���e�'a�ᵪ�VrP�,�s�8;����ဌ�̶dG$+�izԃ����x�yQ��T_(})7'2a??�����s#VP�/{���P��Ƽ��,��~CQnA���~�� Æ1&`ZG���҃��|���~���6F�`��1@Ӑ]P0�6`�[d��~��K��ʇ�}D�}紪�)����͙\]
��B�n�z��}l~��FB
��M7�ڕ�t��L'nO1�mD8�ǩ��C�e�k~#���ʑ�2̈́�#5�L`Oc-�3JQԼ���=�RSw�ҠX��%s��o�5���Ab}���X��]53�vb�(�H���Z��� U���ж k~*�DӞ�۴'�W��B�N��jm�K��&LLq��<�w�"�B�t��$���5�������{�ؘm�����^�bq����f�4Iވ�2F�qBPlD[��÷f��s��#%V(�����˖�=��zO�V}:w�kI	��{"aS�_�5X-JV��zh1��XW��5�/�.) �#�_C�۲�qh���O��#���ڵj����m_��K���>^{aPݣ�����h?�[(A�� GA�K,�"ۙ�ӓS�x��B�*�@9���t-��A��S���|�`.˕��0dM�v!u�c�O�cs��͟�
�6�П�P��Z�:ұ^���Q���=��5��gI�Z��wR��m)oA�fY�W��V{t��[UJ�HP솖C(w�S��M�U�e:�&1u(�����z��Z���%ib3�w�4�m`�M��DM�-�.�V㫄�j�pL�G����]e�� 7̃���AmCr06`��1�ϩ�&�ʰ(�.]]Y��\@��b(��}���d�cF՛
Wr���X�R$O�,v;a��Ǚ�	W�hA1B�'d+��D|5�Zn���Q8�fq�t��O���h>%t�N���럒f݈�p�:`$�<���xKЀ�x]�����W�A�i���X�~� ٧��l��H*�z��ױK�"d�`%����!�b��}gP��چ&C��o4�DMڂb�Z]?����M�6�㜒9����v�+��^	\�s�7�s�6�Ō�84�P��g�ʀq��?]���J�۶���u�	���g�tP̕�{<a��o��Ճ
>ÑbB(�!Ο�I��4��m�J��[�(��%x	1�3Ux����p3�w;�]5U����0���[n����+Xc����ߋ��?�~m���G�k���޷�h�m�W+�|��k�b��(�dV9��b�qݹ�4��P,��;8w�F5^&�-`S��z���Śj6�=�P�������4�[�ν�6E��/�G<��tJ�R0a�⾊E�KW�#���ÆDp웈��E�M��ý4ɲ��d8�N	F���ٜ�
�����5b\�j߄�+-@���X��d��~&ɛ
4$1⍥�B1��iR>^!���<:�!^�~uP,imMY�8�ǃ���Z�c�jO�	V�NWeBe���������!l�3� X�wܣv�� ����D~���*sqT�!_F*>��|o�\��3�M�7E��mC�k�����*!�5 �'�,���[{ϼW��E��]�}���W6(����-���s�L�U�kϵJ#�����y�M�O��xs�Nw�KKa=�ЬH�0�i +��:�b^Qi�Z1�kO�P~���@��b����^�ܮMU-g�ߊ}�[�>�]6_Kr��q*�xB���L��m��ć�,��1K�$6I]�b�8�(����8��4�S�|��D`��Q�>�ς�N�.�;~$����%m^�c�����Ԅ:�o�$�m���{��.P��|�f>Y�\�[mk�m֝�m(Vn��Af��˨"�G�[��)ȿ����y'�!�䪯S�f	��Cn?�	f3�ƥx�d?���Hϼ%VW��36�u7��f9���E9ܪ��J"Y
�X�i=����7u���1��_�1P�nT���]\�݋�ܬ=�1��P��^�O;��
��mn~5(St7���/��Xs_��<�H���p�����ȟK��K�YL&��<���*��Y�p�:~`���1�.�[���G��
��RL�R�gB1��y��$Tȉs-]Y��2�؃�p^��n��A���e��XT��⾪�����&&L<{#{�Pl,��mk��,���Y}lO���q;����R.�EX���[��a��Ckm��,�)�����le�#��
�0��PJ�b����%C%�-��)
h��ɡXY�a�
�o�sC+w�O_�}	����~tY�������k��������L��f�E����� r8�����r�����3E)�,�>����:��^�b#�1	`6G����-����������T�g�kC��W:ג$��Fz�搘��A�>�U��d���o}�x(I+H��P, ?����6]� ���/*�BOi.��w���7�U���+|8g�B�FӐ��uEۄ{�\��{+mW�L����^��Vl�4&j�ci�M����-�w|� G��8zH�#l?!C3l�w��/k�DIx�V$��+޸o[WGn�������Ҥ؋o���6I)���C?��V�tK�[1�bW�P4���������,��N�#0�?�p��ĩ������
��sx��PL2v-��m}�%��ݳ�P�ا��	JB�]�3��f&(���PD��Cmj��k|7��?�B1�*�5��jձ�����-u��*t����h�
�}TH��K�c�x�6�70w`10�O�l�ڑ�J�OX:�^�s����1����o~�7<�3���_P�:WR.�1��|�0���37QG�������fKFm��ӜK�ؚ��^;	^�D�mbq�藠�K`�R�1�3����v�QoH��W�g�r/6��FcE�����2U�ZZi�����ۮQ��S��O�J㐛�p{�?����7W(��c�QK�zh�-G�h^D�c(v�%�m����Em�j{�Ug&�SZ�;`9#��pH|J#Vx����#T��+�sy�:w�7xO�7pV��w=����������Ә�������Ԯ%m�.d4(�;�)��ٗ�5h�p�(kw��'%�Dh���w8�߀q3%��"{e�^ٛ��B٤�(;++e����쑬̬RfBe��.�z��9��<��ǿ�뾅�ls8KB��ZsJ������-
���M����N��Mh�N4+����0���^ێs	w���p�5'i�cƗn��� ��&�6�I�\2��[m�3�4ڭ�$�Swd;�x�Nsfә���󴻱�7�����^1�ؗ�<%˷�,/˄�`vҬќ7O\��n̳��vY�ǚ�|�*�����(c�����",�J�m��4�%&"���ʼ[�.�]�°u��M����}	���G�1<��c�ۍ��>�j"A�U�]aY\�^����9a���3�q>���$�����ƚF�L^���I%3�y�5�KhJs7�x�B��-:��f��7s�t�u�1,�}g�*��߲�^ܯG���x��|��W�
��a7���ul6���s��o��tm�w��Sշ��~�U�9��9�d���5���X���|�7��i*��/MB�]���f��߾��&�	�b���i�v��v� ��Ks��L
��_K�'_�.ͮ��d��&�ԙ�??2�ʨ{�P�u�Ձի��e`�`6�ŰrJ.��IT�N��<5�d��77���|%t��<�&g|�`��Ȭ��n�>��\�tWkv����Sl>�1a��ҞJ���f��J���r���?�E�ݕ�;T�aZ�R:kz�O�j�9N�n7D7�	��6I�����d,	D�L���vc���CkUy���*\h���R3�ݍ�Q���}3M�m��g����wm�wco>��o�.~zR#ttcW�M��Xnm�]��jy��7�ɥ<C��7BYU�߶���ɬ�yq,�e�:����(�6�B0�bH�{�ҡa�rF$��"l�pt
e�J��Ee�~�%�,x�q�4�v8`�"��7�X���>�S��7"iXe�!���=_ʮ�[���9a�t����d�WU=o��=R�񛦳Q/Eu?�Y�e�Dp�^Ho�֚�z�wo'[2d�;��I���J�x���$?�V�1�u�Q�E�+l�[;�������l�%��!��������:��Ɲ���M��p�&w��'$(�-��aV`T�:��{�GG�	�e�ݤ�'�.-��X���OAR7������Q����ԝ��e+�6��n:j1եѐ֪�0�lJ���8�8�e0�����%&��G&ܗE�y2��Vl	�v�X*�W�at��F�a�E����L����T��Ƽ�;��?}L}�h�"����Yt{�sWH_B��vҽ�f��F���nY�`�`!`�o��	1wˊk� �A�M��\��R?Y>�D]������}@X�;Va���1��� ���[r�݅��ۆyk5�ho�����>Q��c(}��|*���i�ëO�{o;H=�����m����V���V-��tȀ��M�H�T��^���hF32@@�?Q焇3֍�6��G���ASO+�	:��n��,�%�y��Qj�m�nX��W&.������8o������=
b{���K`O���P6V��=�qp��RwcӸ��Կ ������&b�S3�k��Mn�%;��RJ�A�R$&'�7��z���̩�-Q����-Gѧ��>�0"v��~b��P�mY�{��HyB���y�}y��`L;ر�̳�|R/4�|��=SNo���ӭ��~{e��R;��lV���Wt�*1�neH6�C�r�ə�d�	&��|���.��ܷYA���K��me`Y`�`�x�z���J9�_��#�uDsR�q|�`� ��#嬬1j�a'K�0q�WnV
�o�9�O�V,b��[R#��}�
_�%w��w`R`���A�3bχ4�
�4�\�F�1i\}n�^+{�˯.	=��ɱ ���e���|Xj�%����F3�z��PF[�bLf4Sv� F�vL�F��B$B�>C���n�l>ɗs`�B��<Zez��8��錗����"���$0��E[?�g�(�f��x7�L�!�K���s�C��m8����X���w}��lV�nQ��N�tXw�Ta��
�����F[��u��=�]L~��f�؍1;y���W�t��2*�X��D1���߹�~�1���q|=��&���l�˚��A��)t�`|`0,hC&�2ن�с��*c#o*�7�vcE�՟oc�g�|j��ژ��O�ߍ6E/8/�������c��M.����ɯ�+�+ėn��d$M>T#ߍi�y�H�Ey�|9dG�؝l��o۩�qz]|2 k�B���OkgB��s�U{�Ӛ�Ղ�c�_]��e.~M�1U����qW(�x��Ƣ�Cl�%�Ԛ��wX�Ѩ9G��j�)���|�,c,�m,�?�i7VS{��)���޳�?�^�}A����H���S�?���o�~�V�0e��6�vga��H���e�(���8IP�;��G�4p|+ư�`%`�?�9|/�l��]�ܹ�C'����	Vn�n�������dny����{H��z��������S{z��d�t��`t`]G#qpŬaλ�kC�?oe&N���m����܁�e�V�g)ٲ�r�z��1RL�&��2KJG��sA2n<�%�	�۶E�,�,f[�m��9���o������-/�h��/k�f=\���߾
������\�A��6�3Ȥ���f�0;��=_g.�H�W�N��Hd�‶@�-s'6;ᰭC��B���B�+yGzS��NǞ�1��u�E����PL���z��
�S�9�.vSʛ�z��`��s|�̈́m���N�*8�1�&M�v�z�ҭ�����
�,70�>�cM��rK�J_���Ͳ���u.���4:������ѩ����,5����(wq��� �K�d���cuA�L:x��c�WF�>i�������)W[9�
���\ҝ;��@J
.V'���9����1�z�o�!�Cu�z�?�� 	Yƃ�I��Ɔn�،qcT�/D��Q&H���Cj�w��x�q.�Ub_7$t�s{��=�ŖE�^A�C�>�u�-�zF�N�$a��@ӈE~�gQX���f�}܁�{���^79=M��u7�a�-/�,Rԥ�0�M���C�`1`GQ�Z��bP�+��-�g��GG����Ƽ��c��f���`�f���ܷuw�=�~����w0&W��>�wť������]�7UO��C�j�e]R=�'m�wc�v�=�ڛ��띄L���^?��� 2���k�ĳGb���T�1��ƻ�g�zVg\���M��
��؃l��ܶ�bn�u�ٖ�K�1r,.Q�$v��%�*�E���x�1��Y���I��u�I�:23����)};��c�s��X{���'仱���d�S�+M$�ދ�v�*����xԋ����p��)N�<T���
��ł͂�+��Мq��+X�cT��k���L��m`+`�`%`�`�`�`�`�`�`j�m�#1�b��V����Ի$�α�U���Y�=��k��vsēLyE�����	5��k\]�-x�x�i�񀍁��	�����vL�RՓ����#ڤ�JZ����(�������l
LlL���}9'{�5ۆU,�k+7N%Mߗ� � ��
f�l���ǫn��H����>�#�>�[���f&V6�	����{���W�<ߍY>��lˤ~�Nc����2G�"0f0U�%0�|��`O������Sb38Z����%b"�7��������\0=0�N��`��������\��[U��l�퐰ps�H��W��!�_`G�R��T������XZ�O�.e�p�0n�\�8�u�k=m�� �]��`$`��������-զhUjJ�~L����M�98+�6E,�4��S0C�`0-0]�20��@'c��}�Y�k��k����`�����.�����2��x�p^����cl�#g��&;�z�)���,~��*�T�N�ON*5yQ/W�}ӿ���ƅ2v0�m]��/��պ:ז�ԑO��+��K�s� X#M�Ӯ4�#�K"n��;`���,u�T���A�ؙ�0Z�Iꁭd��]*�
4ؼ=D���Y��I�]��=0[��b�Sӿ��`ֲ�j���-?"�U/����fG�F�La{QݩJ�/׮�Rj�I���A�q��e��H��]	6��1:;�C�W�̫9�X-�j��K"$��}��'��P��c�n�ht(�
G&��=�T�2���{��	��P�I�Cyl�)Bw�)�9���-���;�J�
��E#���Z��lHU�"m�vѭ�A��iaq�����(_�YIe16	�,�e!�]8��x�9s��J'<l��T�m>�B٥%�����c[�gl�[@(8��e4����RZ�~]����a&wUZ��}W\U�+b-��4{��G�ָj<���}��v��>�쪷��N�6}���\1S����z��	"M���m��
�,��b�-۹��-�����fk(�{L�p�6nkL���~��/r��r���tc�?L�(��B�50ʶt]S�7���_D�A�o_�B�w�Oꎸ͒���2`�V�b�
�,���l�W]��(ih�u�!Üo�A0~�*�����	�6�܊Ŵ�f�%|������

їWWW0l��X0I�T�F� �VZ3�'�~J�Ҧ��'|�Zx�#t;�n`tˎa5����NF������|M���K�f+�HK��EwKL���Z!~N�u����d��Q�~i�`�`*��{��T(>��RX�:��y���jNoK6]
}}QݐBٖ�aؠ[�Q�;&�Lt�oM/ќ��/����X��,O��/�5_�8gh��~�����R���͚�����w��
O)����3N�z�\g��_y6Bṟm��`&�N3�ka�`l�ڪfݠ�9��2��Jm^q�&��&�xE_N sGY2X7X�(� �t��-�B�^=��[�f`��E���F�X?FZ��܍�+e:�?6�uĪ?�����S˃u�M`XFG.;TC��e�'��p����t�����U�G`Ka���i淌 �.�lX
X��y��B׫:'˔��2Z�!��,,,e�LHK,�+���uT��%/��Y�۬l�Z����c��X^��Ɖ�Ժ7�\��=�͏2]��#G�I�yOG�atT�r[Ƈ0%�1�)M�2s�
b��`�``�`�`N;t2���8��G�U�s��7��˖x��*�f��s#�f�1BW�?��q`���H�B�T��q�W�����L�n�(��CE�����h;��bi���fO���T�|�C'�Fe76S���Q�L,��+�0��w9s�dՔ˗�oD<�z��ɂ2�a�u�1����at�`v	ꌷ��U�(/�ws��f���*i��N��`���k�����h�j��29�GLh�fŗsc����HH��W����5��̩*���P������~@����_>��;0b0�	0�Q�!m�v��E�vi���y��)%�7Y�8`gTJ+��Y�6҂���F2�&\iR6����KJ����j�+G�F��p��$���r,^,�iR}������=�����`A`�`-`�`�``g�wL��峂jj��~4�ʰ�U���}��4Tw�<��=��Wd0�r:>c�6�E��;��l�ހŀ����a�g��mU�Y�W��o���|G��l��&�l/8U���>��-���M�N\| H.:4ޛ�5�C�%�X)�D_"e�`���t���ˊ6�.״K|XD=��Q� ���\0m�����������[R�ה�
��?��8K�ĥz�����-��0���M��=��ޅ�E���kDX�����������rP6~l���}�����Y�����לK��鷽�s�� M
�7޳$��m��o���=��-�hM������5�3�h����-��V�ݥ����ӎ�]�Xփi��p�C�`�(��;vL��;�;1a�k9��czWrM�{���g��Ҹ�V���`t�`�4=�+��.�MM�%���ɽ�]C���7���at+��$kڸ[&�����T��=҃C8F`Gm�-����0g�р͂i�����ɝh�r�y�/��He �,Ll	�eI�H[ ���OU��Bj�*}���C�..V��Y�3�ޥ�����l�S�c����5kޤV����c�R�L��#�)�7Q���@�FG�F6�0�(��u������y������X+�8�X��7��G��5�����_f��|�5v�-�H�����D�m�Q��i�d�*�Y������$:m��+�V�\�wc�cҏЕs?;��V'�'�I��;ܷO�@W�8-�� M`�����1�e�`�`X`�`�`G��/��Hٸ�{'�F=N�#�8R�2F;�E�=s���J�b��ƬYUM>�/��T���0����i�`�`]������<��T���<���^k��="�7XTE�ᶔh#���юM�e�֊�����ZnԳq�D%��HMIJ�#{��22�E���R$
��r���s��.�%i.l*"f��6#C�S�i����*%MR.�B>�yVR�[c �j$i���}c��N�W7�x�G&��7*��>'/�k�S�#0�c ��s � ���1S�NxLD�UK�&�t��c0� XX>�����j=�������4�o�f��[�uj�jbXX!�"���87J�Ѧ�D��L����o�\S,����8A)o�4K��,�TP������������d��W(Ֆj6x��~�F�2�y�遑�����;j?y�K׎��)�H�/q�u�P���C``
��sHa~��* ��̝�yz�����$:�1��St�5�,�J��-#°�U�հ�^��T���e$��o���S{f��[EY�0AI˸����?c���	�I���b�F�$^�fCKH���a�c�<Ja6���?z�7���,�ylwq�h8�X')��+mu�����j����.�R���\�q;05�)�E�񃹁�s[Dw*����٥�(śOX����"�LLL�� {�֎Ga�r�S�Yz��oqD��0~ F֋aݜ���O5ƶ���������$��%�)|H�D��,�VF�L�P&� ���L�K����+%U'<���(=�� �f�2�N�-�逭�i���$<����)��#�mg��n3��HK k�������%ŊpH<YBή�8}��^D��oHk���'�C�݇
90�Cۘ�+��������{��~�V� �>�o`�`;t=�I�S����pY�|,ׇ���I=��sH��c6H��f-�Mh�Kn�89�f��Ȳ�"©r)(�>�䰘��b�"���9*�6��:�Y��:CwXR���ʫ>-`_�%^{�HUWM��a�(����c�Ӑx&�r��g8uBD�Q\l��o>�VB�F��
6���q
������>�Ī�I���}13Ji{��*�N�����0�/�����5Q���R�"�W3�����8��p�VsU��t��7�LPŘh,)wE){~��&��g��(!�#`w�R���p��QL�4l06V��j�˗8O���$(H~{Px̘��%�mVʀ�Ǥ՝�Ǚ�4�X+�{��'��E�3;�Ա��mg���j7Bw�_]7�U����9�HH���X��+�/�
����-�����%n�J�6�\}ޯ~��e@]��(7����������8�s	��q�Գ�1z��l4۟Ayo��{ ��/�~��hK^7�gȾRݰ��淜C���6��,E�Y^�˿0���Y�`�`�~�ޕ
�X�!��_��x�I���ai2`e`�`�莖_�Nc8�bC��ô�����'�P����0:~aJMCw�a.rAi��{��I%lCJ7v�phE�$�G�t�w���`���5C<��嗼���=��)o6f
&Ƌ�}D���=6y���'6���:~�W:�������e���n���H��&��1֠��q��ޞ���7��BŹ�٦�St���>#�6cY��y*j�L��eU��s?U���	:O~��0�a�уŁт�;	����7"F�����~/���4�I�A��U��a�q����ɛ���|,�&��>I{q5U�)�H���^վLb/��e�W:=ڳ��3��Itl���
�DIxtq!a�0l	e�N�fCf��[��Q�w���q�|d`�`�`K`f(����0��`��Ѥ���E�}��4/��:.o3n3�i�\_�^�_ѓ���F�|��~��M;��(IKT+XXp�*�ғ7�T$���(�n�Q+Xw���j��2m���JwOb9}vLis;&�C�0k��'|�"R.�:�ߺ+�:��i�`���,jj�Y&t�����ܬ$�]{!�h bg���KX/�'�~�m���ڸ�[ �
ʾe<���Y7�2�(�	m�0!�5���}�����st�ϕ3�ʫɍ����Q�H��0�0����ė��D5�=����e�"s3I?~EZ>��װ�Y|�?���[��/0Մ�_٧�DQz����A��WLτ�F���>�o?X�P�=AY=�~����e�`�w�+{d�C�����p�$���JQv�1�*����<�͸Wx�+mvf�%J�80lƽ'�ٌ7�΁���"�t(���)�7������9o�8��6X��Im,yC��e�uy���N�����c�C��F���{85�$�L���L��(�t�w	���/�3K5Y��'�5�P�Kc�G��b�&����J��5��P���k��0%��v�j�)�}y�&�N�R�h]��x����Eίǥ9����Pd°R�!:;�6�0�{���ft�d0���!�K��8	Le%�HS# ��Aw��)d'���-uK�
�<���AY�E��M���?]b�@s�EQ|=����C����B�L�=���C[(t4&�[&�a���d��\��9�3�w72-	,L�	,���CY����P��h�m�w<��ۀq�Pv�V����Y�
Ye���0�2�e=J*!+#[2Z�Ȟ!�앬�����t��Ͽ��q���+���\3�Ga�ϖ=����r`�`O����w��4�.���?���JU�P�}�S�O��#��,x��u�O��8��M��T����f̤V��u��QJ^��z
����� �[;f��V��ސd0q�}/IQ��!-��s`7��P��H�ƶR6�_0ͬ�7��X��k��A�:��,[t��1��>��~�����wc��`j�a�
`�FQ6�����A��ѧ����S�re�?��h�6����#FV��a�,�`l�}f,hj����;hy�CT�w�?��Y��������l��|.Г<�d�M�_B���}�%}ɠ���%T��a�6���7��Q)q�1�۳"9i�e,�'���r�r�n����nco{�hu.�і庠���B�]k�����U�.1�25��q���ݺ2��-9����¼|�&��9XX1Q]��=NA�Kqj��B��QK��X�:�*��۪S��k�g�Q��/0�r0�K``*5#��m/�3/1�H�w;�!V��5G�|�C`���X^�o�5��ӬI���
��cm�le��ò�L�T�-�����:�������z^��:����`9��(�D�E�#,2���HJ5�m�u.j�l��L���$������3`�y�6<�9��9k&~��~��ف'8s�=��+X(X+Ƅ�Z�+_���������7Sgӂ��+���}����N'���1o��kޫ�_H�ytG����T*�ـ}���S ���]|&>j����_!7#��Ï�Y��`�`�X�	6&�ᯐ��I󜁂E�����=�g��㉲i�	��`����������⼀i�	�����.�����2�ʙE�(�d� ��L}�����q�e��➲*	0����!Ftk`�`�`�����l�??gK@��e�e���k�X�� cCٿ]�9���r1�I��k)oHH�|������'�<g���{H�c�QF������>�@�ʂ���Wc�~�p0Z��`�N1�x����72%����ݚ�iқ=l��X�ϴ��]�wkD`I�s�!>���܋�$��Oq�쒅F_M\gάB6� ����O�G#�������<{�160:0z0B��`�`渮�s(�oே=���EӮ�6���c-�	�,�a�i��Hd�,dN��)s���3�Й@�*�(0|�q�сI����lr&0c'�~i�T��)dq�L���r)!�3���رm��@ө�y�J��v��6N^5�YV-+@fF� ֊��9�����q�9\���hEd��!����u>�\tk���a����^BKhM��%>���1��Bt^��^��������4ɟ�J��8<��Z���1�yT�	�7	����8c���)�*0r0e�E�z����16tP�*i���?�����WnS&�Z5X ����A�]6 �4{2��Q����ٕ�^d�/�����(�^T�zٞ�&aO����f/F��E�67s�P�a@!fŸp�9�.��#����FF�j��;�F�=��)A͡�6_��>����}cGuo�N-��(�}�D�\�+ٹLr?;U�%�����Α���sﯡ;�EA����L��W���Ԛu��e���3��L[==Z��50���� V(��Ql>y��鞡v����>9�W`S`$`,`z`�`��bm�r�p~>W@D�i�?	4os�bϗ�]*�
���*�F��"�Y��)}�����V�qL<A�d'GYH��,��NP�9t���5c^=����4QӒc�Z����Ky`�`z`,``�������>�����&Ͳ�<\��������`Z``O��Ll4ӶSm#^m,�܌$?���i�Ӗ��k�j����ϡ�qa����8{22�F�|��B�k;� 9.n�x�z��\h�^ڙ��b����;0��?7����h�N�Q&����-����A�(k�`�����p�I�4���ĨR:?ָ$)jC��Yļ*��	�f���/���=&�ҥ�R/P�iRj��ҷx�nXw��"�nCǗyǞ�����Vn�N�i���J�ߦ�XX4�Y�4��{�.��^�؃{k���;4�����f 쒼
�0	0�a�7����}�O��w�K�M�e�*]�b*�&����]#��k��
{��o�1/�W�%��TӶ�I�W���+Cl,	,ll�9�(��ٴ�7[Õ$wS��A�P����tk��:�d��wui�;j��\}L~�Q������`���P����}~�����������s�:��^2�O��T��}���e!�cj(�F��I��%�Q�.�aX^���=�)��i�"�C�U2`��XXV��w5��j��)U����	�����ߗN����k��w���y�����2F.�x�^x�Fv��&�?B����K	���֏�_㿈T6����|cm󾦴@ڶ&�
f v,�?�z�Ek*�S�,��LP�����i X#1������b4�vY0tu&?�?�||H�3�1��%[�	�a���2��g }2.�@J���2�)�}Ow�<x����C���f_G�V>'�*ދ�76A�Č�������Ղi�]X�cx�|��B��+�����{��5N0S0��]ݟ<�gѹ�E���F�:=:�nma-�b�y�S�[�_�tY�IC�hE�g|J�(�.;=ٳ����:�E�TKR;�í�AL�$e���R��~�d�a<�nw�!��5�s�a0^0+�'`q`وݹ���t���7C������-.a��`�Cٗv����}u	�:A`=G�𡜵����S$�T��V��f(��VQ�Δ�D}�5C��܂�z1��;��W9	���#����2{V����X���խ-s0����}�
>��Y����e����ZX��}�ښD6^����b�;q���A��^9(�&���߿u���a��4l�"e.��йd���I9�x�O5	�9��1g�C`�`q`uy7�Y%e���C%	-�y2�3����#�h�5e0#00?\�ͥyw4���&��(K:�Z�m�8`-
,�e�v�:+$�$�t&6W�")������Zx�t�����H���5�F��ޢL(�S��)<����#��=�,�q�-0Tg�X��j�����e��ݧ��m5ֽv���Ɑ�]&��5>�
#�ʫR66�Q�3�J��i'䴪�J�����.�<UR��,�E�~u�ʽ#p���S2⺕~B56�rS�Yo^�F����#�	�v\�P7SX$8u��>�:)_ߙ���cm�,Lՙ��O�u���O�؛ů��p�����)�C>��7�fq&�_��N��������1�(�O��D��+J|}�X�� ��o-b�T
��23��΁��~�H>�j_3� ��M$�l��,����CX�	f�
6x?���+�A�+�g��$5JrD��v��t�Z�2����E��F���D������\g8��m_DL����pFm�8Q����7�윌2ƬRfr����TI��oԏ�2�ut�� s#����"Ƃ�Y��?myk�Op�+_N���`��XA�|X3�.k���W�˝�����3V�os�Y�<�������������
9c��c�@�,�)l��Ha���jkK۶���N��~#FVV	���V ���uX��V���BV��a�4�b��X3��Cu�p>��?q#�Қ��N��\a{��^�M����i��(�L�p;V�I�B�6۬w��(�g����}�%�}u��y���ۧ�<������{(��	ѱ�����F
��&�u֒�NM�'�_�"v����6^[��x��ʺ�.����mO���r7q�Y���b-�۟팄&���5�zq�o�^�B���.��w�B��?�m�+��~Z�G.W�xd���m�g(�X&XX-)�����JV�cgR߹*���G�"f	���|�+�L�Ee��C��-w
J����{LR��Q���,�U��;E>Ό)�%T/�~��v��+3FR�����T�u�
ޱt��"����N�����q�<�n�0qp�B~���[gq�J�\��ǱV��L�9��=r}�'�{$O"��@w�5bb���2L'��r� �߸�eV�|�Z�̞�%�->�G��͊������`B~�P�����vb�v���!)����ԃɂ����Š�$�B��\��W{<�h8�c��Q�K�@X-X��#�ǋ�,�k-`���(&�q*�S{.�%\�א�F��N~p��g�AJ�;�.�ۖ^�эv��Їg�?l�aK����:�M�j0O02�����݉S�Q���L������sY'��b��d0T�v��u�e��u�N'����,٪�Ű
�1ʌQ�J�}3�����YY��tv�CO�4�Ε�n�4�ʼ]g�Q��1*�`&�����Y��$�.>B�<�|`�����@l�ֶ�����)6r��:��Idt������T�l-k`s`}(ˡ�ɣ��'�f��]]b��{�f?b3l���:ן�޺C��;�vl�ڝg�2�-����~� "�%�7�S�k`n`�`����bL�En۞�*����߲W��ƚ�k0��]�x8A�A�rB�j���T��{��+�ɀ9�т�r�ˣ'p����[�͝��#+e��G'5����K�ӢP��X$��5�3�1�Z0N����fz�~���������Z7�X5��s��S��b���$��/���������֎2t�4�i����:s]ɢb�����_��Eٗ5"����eq�բ��:�_��,��u{�t��\���Y9�偵��S;���U7���Ҳ/r/{Q4�[��R�Ys���N�ړ�9b�mxaM�Lc{4�4~k9r��v�i��7�O�]i��!��Z��U�ѥ���SǼ/�y.*G/�f�L�'�q�� ��++���twwM��wbq���Z�uX�y��,�5�;`�a��D�'�ٚ,^�����J7��V�[��q)�Qf6
Fv�gm��J�c�`b�ċ7D��^u���"�6+�0�w�Ŏ��L1LG 6���Q~N��$��烴��G�O�y�5 ��k^���=�ud[���S���D�ޯWM窨D�w/�>�i�5��߮�٩^����j���
�kW�WN��8n]M�řt3��&��[h�T	��*��;SLL��U���1�`~�D��]�k>z�K����jc{��$�υ]VɎ�F��c�RGnP~~"�hpIl�|��47X����Bb��0�L����{'���0�/ť�iz�՟����mdЏ����)���͂������]zmZ��6^�3�p2&omJƚb��vwIV�{Z�M���R�G��)m[:���``�P֌��f>��0ܱO�F�Q���/}��öW�r�^��uE��g�ر(�A�=K	���c��+��j�vD�lA��X�*�0�j$����n�3�k��Xe���:�'����e�ױv��+>r~�}�m��Z��w6�}r���mʝ[q�dVm���Du�j�l�0&�$�K��n�F�K������+#��Nc�ˬ{C�u�-~����=I?Ɯ��0{���eV�]��TK�s����$+��+ej�!iJ7���c�G���w,��=�ȿ�*�r g�K\j^AϠkϞ�F�p�������^E�Ӷ�CPV�X0-��d0�0�>�������F��"�畾��؏v�I����@u�`�>n�����	���"�CY��5��� ��
*
⿆銡���S�ϟ4�v/���y"����(���ѧ�m�BlXщr.B���%ʖ{A�ę/%j]���vwQ�w1=�5X'��9X1��#ļ�&������'�l��L�d�"#���(�����.=��Q00>�Y}p;9�Ǯ��-���ӎ�b	O�y��E����S�XB�O;=�#ż��"K	O�N~b�w��k�I6[[;���添˼��;K/�Aݐ�X'}�h���0�������F놮���]ַB�#�m\$�Rן
��E�4�>0?�q��7�G�pv���Y�ވ�׍���SG�>�~�bb�d�c�(3C��,�L���0�!���n����$)U��5!v�k$`��*���:�wAm�qO_��8����k-[��4X� c��2L�6f��]~~O�ɯga_�IR���[����(��j��19�4	�X(ʴ��\�~�a��=��VU]H>5�y��`���P�bb�`�
�BZߍO�^kՍ޾SVl�&
�&����zu�f �� ��w�PѴ'gb�o�#��,	�~����[~q��7]�`ֵ���:
c��e��1ncs!����`������Ƀ������)��Z��h��\��`�7�ȷ�Ҏ5g0I0]0KTw���o�:��ƇQ/_��o��^��UI��q���M�y�s:�DU�c��������:���g]�>3����P|,�ܨ	6二2-�0��K���`�Xcm��:�� ��=g�"������B,(	kk`^`�`�rd�������3fQIfw&��vY�M��K�a��9f"#b�3'�N[�*�;�_��_F�g��էeR��C�˨��]l�r	c����a��C���M��t�`O�(�x������ǘ�+u���dbë$�Z9dQ�9`FCX�F���J]s�=�N��ȑ��r��.�}�bf�`�`�`�7��c�N�D�+��܍�v6>A��I�Y>O�>g+�-��|Z33��yje[���M�-�}K��z;����msU�P�M#w_Σ��sa�>X4���sQ>x�*��jzzt�eö�ˠy��"M���h�Vq�k���_��~n���n	
ٵ^u����� �Q��z>y��} !r�z��hc�i�I��@�07�2�K�$0q0iĪ<�vL��ǆJ_��<�Xй/�/�{ؼ���$%w�>����n`�QМ�ZLId�1������ٞlZ+j�%�ŶFʪ|��5�M��{l3?��g���_�+���%XX<��	�A0_����@]�ɉ��QG��ċ/9<a�3��M k�y�Q�E����]F�e{�-L����5OU�ـ���y�%���"��8Y��ܷ纸�;DH��@[b���w����,�t6`�`z`����|3��r��-��w5���F��k4`k`�`������������g����}1U���6���Z�dP�og��t�k���	q���K�U����&�ϕ|<{���F�F�$w�e?D���e��.LJ��>��8�AN��)#X(3��G�� س��r�z�6#m��iR��!�ssp�g�e	6XSsU4� �$�}xuC7X�/��I��s`�\O�]����N��}tek�c@�8�p�p���M��� ��I��`z�y�]+#{���V&�U&�R��kt;=@e�A:��'`_����Q]ئ~R5�$��O�����!0�6���I�{`��bPF��lY��Vē��MY�	>�#��X��P��4�M�Q�����K��c�(�C�2��ꩽ$�#�q�����4��:u
�	ll�1�$����������9ɬ��o��e�[^���ۀ]�뇵ۗ���lu>�k����.�+�"�7�>w���1�c^i���n:����J	*0�����p�y�6,������3��������Q�M�GW�1�s�O�m4�ܝ��<�t3��4֨�&���:��B7�(��H��Fӡ*MX���~ĩ��-X>1؁�mu9��8�S��]~�:1��>���]���[�6�F'�X���l�^0O� ��f�H0�G��M��wNrM�:=�.n�"���`�łU�]GuU`���]yE�ִnn[C�I�}5���v
,e�N���ڜ�����G���6fY=��-$�w�Κ���bn�3ʢsr�oz�_��NHʟ'�N���L��4�b��X;��xv���,mE ���d�}K���I������k'���	`��g-_��^g_���P�-ٶ�Qs��!�V%E�>��N�6�^�gg��)���Ŕ�q'S9��1�I0A0�V�S�;#�&3���7��=��s�d9/�Y�U�9jam�
����h���|�����}K��q��-5v3(3#�[m��q�~/�&�6�2�0�i�3d���ϑ����5l��e_�t�``��t�EG�Q�9�[�v˞�TE~d<b�
,1:A�рE����Ẏbݙg�V�=�O���x�ol!V���`�`S(��{"Y�n�*re��)ZEҒX�C�O
��_��w�'�Ơ[�����O���}���}rcH��,��e!���`��N��=�Fu.��S#�8�{�A�Ȕ���.�����_`|`�`���v�5]���]�>�н0�<Roa�|���/�c�`�`�J4���Gq6����`ݡ��H��J�ȹ��#��+�7\hSDlLl���)?����t�!IY��5����Fm�� ��= �V���F?i��cL�N��V���4�y�ə���XR00:��Bur��c�ż;�e�@�]Փ����7���+`�Du��o��M}�F�b���n�U��`��O��އ�b}$4��E��;f�X�3�$�,����Lynr��>P�?a�Ԟ����.3L���4�Wj���&�f�*�pL��qa]&���m��&K;*����[�8���r.�[���w�cW��B:�9�,���6�4�w��{&6 ��?� �=�'��ݾ�N2"����eǨ7������=N�'��e��Y|��`���pǷ�N���M'���-m�z�n�Dm�h�
���8���,(G������-�5Os�̚p$���[_SG�)bj`w�V��ـQ��k�+��v�<Q��>����v��wXk���Au�����l��i�$��+���7�ĳ3�b��������L�=���Lۮ��v.���Z�#�N��^<���R�nĬ;��km��ZQV�X�/��V����D�4,��Nmg�ك�����-�9!楀�E0��'��b2x(�$&X^���;����
`-Llc��->ˍ~g̮�r�`Ri17'�g�+8N�+V���5������({A���LV��!�K`C`�`&`�`�`�`��R�MϼT%�Xg����D�+�`7������f
v,T1�Yme�ߍ��c�l�ti�Ҿ�c�)�k�ݚ�/����Y��-/�����F��w�c}"�1�{�MT����^��[�M�2�������l�������>���X�,��L�LeFf��x�(��Z���R�x�Q������\�F��gk�`�`)(�������:���oK^�fy{����e�e����~�8S��7i�Ѣ�O`�c2z�n6s7oA�s�2�%I���1�选�:R�ND�q�L��&k�o��Q�;�)�6	FV>�|t�i�c��5i߁�?ܯ��l	���ѩ���E�N?ȫ�k��:s\;w�t��X�.-�5��<�bF���M��n���-�A�Y�V02�S�N+*��m���=��I
��&ze�rX�#�[@u�`-���0�oH+4��쟍����'�)sm����l�I��i�HI�c��+��㛎������@�5&�֎�2Z�t�e�a�y�;����&~d �v�1�FDH�C�&�S0q0a�B�JB�v,l��g������
Ĥ�:/i���rb���b-�)�!���i��Z7���e�1�bh�X��=�>��,�xn#�A�|'��6�(>��H��Ft��e��=Q���`N`�`�``��mcL�h1�<���`8�x^ܦQ�Xh&�L�6����w�$t��2*'	���1,U���Mw������u���%�-TZ����n+C2~���d�Ol���۟�\���l�}`m`��z���D�2�!�4h���w<
߀qB	!Qff�I$�D6Ɉ�2"+2RT��#���
eo);+YI��>nO��������s]B��<�7L%�������i��Оm��0��`_P:E���̮[Ƅ;��]�������{�(��!%�q��/C�x5�0����]��|/YNwt���p�ܾ��_.�3	V"W�b�H����Ԙ0k����)�A�B�'��\�D�s`M`��VN�g���p��~��[�����쏱f�i�|��7���g�I����������dь��ěW�.vR<�;Y.�c�L��};!�����t4�#��K�,��w��3�76n�3������=�;Fv��n�"����Nqi�,Cvw����������*�-X�J�D5��J*�}
X���a'�`)}��$�b�`|`"`L�������&�ʬh�B)X�ɀ��,3�|V����ݠ���]EX�3�E��L�����g���e��"��j�� -�a�*�������;���J�r��Jz��w�$�T!-qw�X����P�?]w�S@&�E�WCA�!��;�����N�=��S�^NHÂ���Qo��[E����Im�9��GC������追�%��|ʾ�qdR���q�&&�ȋm���s��O|����j�v����wwJ"��=�Q75}��km�K\��n��vMZ����z�����+�X�zի׽��c�THLLg\���j��-	��A���p�(�-�����G�*���wّ�3�:t��)1r���nyD�^�4�+�$k���bY-�'�0_�;����Ԉ��-��!~�G4�����ֻ�MÕF�K+M��s>�Q�t�:��mnK�7���=��Lr4$�^�����5�r:Z�+X�o�-�E[�9Dοblr�����Ø~��6��;2�.�_t�q.�n�����?mr�ňY�q��y[��R�4U�V[����ӻR�T�OM���������*0�T���c��7�[{���1��)J�S�i��D��4^^4]<�۫��H�5+�e��A9��ٛ1*�]���LK�B���`�ȱ4}�f��s��#��^0+�g8;�υ�U�6	t	����<�E��%�9�Ѫ���e>�2�67�ˋ����c�`n�	tJ)F�/?�4�J���י���ت�<-��� �?�j����	��!��
&���&��-/��Y*z4�"����8�-�&�X���m�af�u%`�����ng8�|��:[v�;{x�$��m���5 �C�qDD��)Br5��)�3���F5�;`���e#kK�V&����NE�]Z���T�P����jN�)���-\1���@��n���[�����gBZ��_sZ�=Ï�y���z����;���gH���(�{���͸z,׎�G�!`��~�Bd'����^P��&�:M�=�,������Vh<�,�a0J0y01��{F���`w�p�&s[�����(q�.��;C9?��P�t���.�
F]��� ^R��h�7󇱓��r���U�P������M��#`�(����at�雺RQ�Y���Z��>֘�;��F��l�W`3`s��������7�;~|=�	�k���5�i�`M(f
���g1w��&��t���~�3���G�ۦ����`�`�`�(�i%�Ұ1�������[���8�6Ɔ�e�+[��{0������8�Ϭ�z�>cv�c2��� ��V��	��uy`���!��_�}֪>��w)y���kC1W� 0�^��b��}�Eˎ�`���Ү�>���z��,�����$��u�`�`�`�R�X��1^b��25K$P_�&�b���Z�ǬJ3ID��o�u�Ė�Ib͛��n��؃%.b"�,&�8�,�lL�`ϒ��͒m��X&R��e�_�>���
VM�ʍߌٵ?|����&�S��wr���$'�0��E0)0r�A�3`B`
`�`�'�_�������?o�K_r�I�Oc;Ƌb�����a�`I��p��9�,�e�g����
W
�3+�%X��/����/'#D���z��!
ݯ��`�`�(�PX�a�`2`�`yf�F�+{^i�y�D�͏��X=���/��P�;���S^�3��0�pMg�Ã���sǳط]d���9�$|�ދ�ߣә�m���o�i����~��`��y�D1��9��\�+}v��X�"����}�{ �脑��|��p4t<]�j�ƛ�8�6
���7�AZ�S��Q	WcM�Q�AҕAǝ��7�d�^�V�l:#�-#�m0��%��ܶ�A���R��
7���~�b�r��.����g2M���)��7e�r�������4Ҙ��9�W�`�;2"�I�?7�\Uc�:��gB�U�!ͪk��wz~���-Yq�p��������X�`a�E�k��J���WG���x���ŵ�R�$��ARٟ����v,�KDvbe�+������Tu�Rm��Ө���U�q����D�~�(��:�"��7E�hʹ+�I�	�D.�k�n��,^ľqK�e^�U�pe��")���b�K ��C�~�o��82Ca?T�[cS��|�-η�;��w����a�`V`n`�[��<�[Nf��},_�k�g� V�W���;�U�~?V����٧��RI����5�����B���i����w��ʾ�1����6x�Z�NL��/� �3x��a����q����$_�v�;���@;�vB��c���L�����IDG�+_��[#��5*E2Y>�>���`Z�Y<�6�X?_+�a��`p7�n]H���ט��BO�9���i�̀�E��u�`glR�g��7����I&�����Q6��b�����������L7�O0�e��J��L�̩*���D��%�r�j5��[`�`_o�����E� ��뮹�F��sPLi�`=`�(¶���M���5��x,��5�"z���#�v�/:�7L��� 
i���	���D�O�8}B0�.�D����P:Qdg���̾�c]-��ͷ�a*�6��My��``21�TB`
``x`�{&�4K��e�-V3�4��+�V`f�����Hd���2���Q;v�Iڏ��"L�N�M{�� z=v=l��!�|�}F��w���L�,������h���#�&��ά�sS�T�Gtm`�`�`i�Z~�6=F%�S�&GN6��B�6 g�gLH+�G3�%��_�I��4�<j�}=p�I�,�d6��v㮊4X?5�Xt[,0���K}Y��ΪӨerBLybϚ��v	io���x���G����Ƅ����W������	��6㺪\vL���Bv��Н)��A�m����F��D
�Ky[`HK�F�;0B�T0&2�E�u�����t߶��
��<��U���:�,� X�$t���-b�[@�/يfK7G�E24��=q�/�=�@�?�عQ����/�;6��e��^ݲ�:o���h,��1���q-�uB`�`�`oO�sv�j�ļ4y[��$C4���.�]�V=�a�(��7z)GI?3KY���p�~I1� �}��¸��>+&z�1�-�]�]�3v�3�)�E�d�����¥b���������[
�(�]����Tl��/�Ǧ���E	c�ow2*�E�m|z?GVv�;�Ԟ�#-R�0��4.e�����OY#?��$�X,gL���4md7H��\�<�6M��U�Կ��@w铍�D��Ӧ.0-0>�G`B�{���0N����,q��Űn���:0��بC�
��w�"���l�l}3��s�-Ik���C]ݱ��`l`1`J��i?�� ��*�Yh��zLl��Y��%2�E��[�r���~?
�6v,:�Y��h:���X��*����֩�K`�N{F�4Z0u�т=��wTh�Jm� �V@~�V� !��K�!#��[DY#l��;�J'���=.�	&S��#oe�^��{f��`eH��� ku�KG�K���ޮ���q�s�����}���rWz �.X�s�:dg�j��Ղ�vK�I����r$uʈ�~kV��bu`g�L,���睿R����z药���9`w������o",,�|�s � kS���{y�T���Tq��ѷ�d3��6�N2ŒǑ+h+̛�hd~jj��L��E���A�&�ާ��]0=�H��)��x��E�_?4�3����x���S0��`��(����β؅/MO��W/&����_f/|2n�+��u�X�<��M��W�4��K��m��C��Y��ۺ��1��Q��1�$�EX"��DO��R�|H����'�w�M8��{�����N���L�2
0+��5=�vXIOf��%XK�*?̐4f�b�5��|���v�����YV���}�o�8M���b���f�����X��B���:���5A�<O���ΥGر�RE���+B����'5'���G�ucἭ� ��eh`#`~(�6��p��5�5r�+"iQ.�K��op.(�-V�5",��
��;� ���#�~d;�U��|�7�v�AZ���L�������f����k�_��r�U�����D�?�j���xQ�S�{�#���ܞڷi'Ю⥖s��>��E1\�j�}�qX�޷0EOM���ԧ��)N_>CEa�p��lz�za�`�{�%��,��
�OKE>��2�%'B����(Vv�
SX a�(����&o��-��4�)��5T�K#}"�a`mzJy`d`�`o�x�V,Ua�,���z��C�3��,
,B��a(���zeJ%��vGv.=��f��tF��J�(�(�5y�m0A�W`�7����N^�e�i�3V�?X�_�e��^�GX�y";C�~_�q�v�p��jܯп���c�0�F�f�v����� a։�\���O舚y刼��9Ƌb���D`��O� L����4ut	� ���b�6�Q����`.`ڒ��	�n�X�u�ܥ��Oj
ǚ�
�D1~����[3;&�ߝ5���s�_����!q�I�~*���2j0�?>�z9����:�=�@�D�4��j�y��3�4�r�X���v�cFvĈ��,���Oh�Gω���D#�=���EY�����lb�N=紺fQ��!c���E:��E�B����[���,�Nƒ�,��:�̓��͖o���z�{��{Ώ��5��\;l��&
&p~_	�L�LL�G�Gh����Ƴ��e.U��$2(�ƃ�~N�[s_���S�F˝�F'��������x�u���{v�im`�`�`~��$v�Od]��ǒS���l�3�]�u�y�^�����lŮLf���La�U�����99a30���^q``�`[`4^{6���,��I���m�$��;��e��>�l���o&���;3��Ћ�o�*,e�l/��lT�����D�4�����`߲db�����yj������VY����
tZ~�H[p�xgy-"�&��x�|<���ƅV1�{�]D�9�ﾦkS�ݔbԊ��x��S�ԲPvLL�#�&�������|�/���=a�s��{
F!���y�=;ƶo��x��qi4t\�$���R�O�_`��\`�>zߜv�Ak,a�!�ۃJl����:$7�ۊ~	X�yq��<{�i�;����U!~L��m7��e�݅v#Cb�;f�H��+�pɛ�
Z�����Lt!��}�\�ԙe����`8�&�tB�I��Z�>o��ڗ��g�2��w1Ȩ�'+�)(�E��'h'*<�J����G�p��xg�?ĩ���dp6�s6)n���'���P��fW���C����.<�ْZt����*~���\��͋�O�ߣ�T�w�,IH����{�45�z��������FXwkJ�/��.�z��>杯S$�����Gb_���a�#J�,u�.�`#�رޡ�4h7�թ�,��5RY��^���jʦG(Wr_��[��ę�'L�V6E�������2_!�� /leo&���n�.���~��q�(��y�
����"M����=��4WK���Y+���&�Τ��M���4�/A�ŭg���Ƒ� ����Y��լ׹���g�0�� �qn��C����f	��Y�M�Ja=>��d�hד��
��j��i��&*�ߐ���mIG��,����<�MU�g9�L�+�c�ם�a/��ͅ+�Y��!}�x��>�$э�X��u&�>{c|�Φ�ن�o�O�w��3m�%[i�;>�3'��_�ψ�"{�>K�b��٥�XRE0]0t��c�,��^����)�vy��<�S��h�ϥ��4�F����OcN����f}z�n�}�l��*�h���ua���3LH�*m��y��ݴ���?�;Vv���֯t$&��u����ң���+�|��͛�0���(MZ� �r-&����k���ft�ɪ:��->T�\��B��E��*�}S�}�Ll��� s��8�Jj�g�V���hG�����:P,s����,s,���i�����e]M�ka�M��Zޘ��,t�ݞ5th&����$S��*�3{�av�@�$X4X����kh�������^P�p��Gc����$�M��`���>}t#�I�h�Z��->��8��%M��b���[����НO�K�w 9ݭ�p�ն��m�B�V�
X��u��m�I�~��`^H�6/� ��^��J�ke�<��>O<�U�E.]ӻ��r=����S���2��C�q�4�x�V$�X|�!���|,�e�f��ҁ�Tn���m`�Tơ�+
Z4�����e�zt�7d�x$��^O����|,�U�wW�J��Y�*~����6T����1w��O��c��kK�>;�I?��n� Lf��ZdZ���V���D�Qf��:iTc��r#v��f�����K.Q�w;�Q�(]&i&<���M�h7�r�ɤ��]M�P{1//��C���~��X$��b��&��R�\�$��2YK��v� F��@��觴��Qu\é���1�1��!8_���5����al:�|b'Lo���I���e`_��?�mw?��u��Yf�F��ׅ��x;� ��u�/�l�G�Z4jΐ��Al�J�)����K6$o�g�v��:��D�����|��x���Ń��í�bn윓�W����rd/����.v��o1͋��$���:�=:]ߵ�~OЈ���B���ޕ� &V�V�]��*|��(2����<12�AUݮ�\�8�l��o�a1��Z�̫zIq%�#�����8b�c��N\��L�QR�ӷ�Ⳏ��r��^�	�T%�l'_^?�q[��kb�	����"'eHg��A,��M��q�OJe�H������bm�jF	ɉ�Jk*OVR:��%޳�����]�؂Ly�}H}?A��'+��{܃�������|����S���5�b�W��/�8���苣�4�����S�e!={U	� �бd�����#b�L�����೽3Y�[�y?�nyO�r�O��x���hVa9�o���h�������
]Ec=���q���'��.6�\�t�﹯+.F���ɊQ����嬿�O]���|�U���r����M2
�b��R�-���������+��r�L�����jX�y�+����?�,E�j��������:Xke��,�n�o�U��\�G��	L]�$r�%l�[](ʔ����w�q��_��~�ܫҾ���GV���M��f{x�����o��mJ����z]3�Q�#�>k�`?�^�b� &�1V�TbxS����cY�\����V�U�_�ue�U�͡Fw��S�����	y)�oa6f��{g��� �1�2gcN��V?aѕLb.dL����4ggF-�Բpk$����Y�f�d.<��
�S�F�o}��q���x�����`Kͅ�.>��$�)��2!��-�qI��6�����@E�ؿ��95��?ȗ0���L�۹��阉�^3ߍ�Imӱ�S�ڄ)����;�C���0�n�%�"�V)��W�yü��6fc�{�6��%��[��#buN���nX�Q�����\�����#̑<e�h�g��,>��뜓!V��A�]������|2������N�fm���k��X�=w~���z#Цq{�O����㐞mc����7���b;\1�_[O�U�}」=��(��&�i��o�����?�$�IcK&��"���7��L��ls�r�uY{�Y6�d]�ߌ�F�M�o�Sl�IߋT�����;��DI�����\����)��6b��.����%�C%~6��.8�_p�x���T�����aiD�ױ�O��l�c��׭�D�,�8.����z��-�R͎�F��� �q��0lKF��J'Fҙ��x�=LƁ���O�r�v�U�o�q��S�ߵ[��F�&�dc?�aj�O��ҵ:��F^�=&������'�q��L�;�Oi�c�	h��,��/�X/M	����)$�E2M�u���\��a��D��|YM�|�	����\�A��l�W�����ݨ�r}C,��N�f�<�8:$[[qD��FX���?u��l��M�[8:;'�B�7��b�2�u�XԜ�����$�-��Ȼo������i��4�W�Q%�s"H���sJgU��g?��g繆dUȈ&������v�49x�g�/�8����׌�|�+ۤ���F7~��A,V�c�I�]�X����ә���Z���C������;2��J��Gb�_F�X��>xy��`
NX5?^(?�	p�B6��੖���[��!��o}#s\{S��h��M*��̒~|��Y!�<���y���[�(����ػ�G�\o`�8��yj_����A�n�맄�JI�b�M���ރ�BqM4���N�>]���t�ƃXg�9�W���~��ᯬ�Q��<�=��Υ�R�v$���뫹>j�q��=��ْ���������7U��1ڹ�w�7�z	_�����g/x�/���6͝��$nSZ���({ɱ}b���ʓ��q�P�,Ŭ G���A�A4���]S@n@�s$�O]����{f����B����E=�����)�j���<ʱ��X�����\l����W,��)��L�F��Gq�Q��������HӼ��7=�Q?,������5J�Y�d�G�/gJjl[�;+�Q�!a��.UA�����*�	�X������6dy���Nn���$�i�"{�@�\*|��ש��s?N�5� ���u$��٧=��T�����D�6�����]2�k&v]��4>)_?qu��D�KS�gܮ:�1��6O���p��"ªy��Gm��'�J�ס4yE��{�0ݤg�����t��B�h���UX���aJ�N��[��P@�K$�A�D)�n���ؔ�&$�[�uGF�������Rs2�0���8�%"��'+!���}�ǿ��TA���Ԡ�;2�����r��[Aʰ.R�rf�L䷸=t*����x(#[q����0���i���}�k��p��g~�L�E~������:�1B=�C�lBx�u�����Q�f3�=}Z�7ؐ�+�5��k��.�P�iv�҉d��V'�J���`�O�̕}�]�?����c:a����Ʋ�p�kܼ�������)Ȟ5�X��3˜�u_,�h�u�.��(���/ШH`��ZZ�kuktaci����h�j<��*�+�"���IÃ���~u=��u�9ش=x�>�ڷ̍����h������W�t���Be�3���7D�C�.���&G��80�����&|�\!G�y�`������C
��a>�&ϖ����Z
D� �`F]4s�`�=ܤ@c#�o�f�&�r���#t9@�{zRq��W�z�n;d����:��A�W�aڏ�Տ���:{�����TW���czp�.�59n����|3����0�:����v5a[��l��7@�GMG��r����;��yn7�5]��z��w�����'lT���e�*5��t��>�D�a�*���M����~`}�m"��[Ϝ۹7�t���(�8힄6�.�j�Ȱ�!�
����8�\q��a�ﯽC3�U���X"	���Z��3wG�.�"_4Ǝ��|Xl����f@�����w�k�B���T�֪~_t�rS��Ma]��vgؤ�/���AX�������Igg�U"(��Qk��m��`zXU�B${�-لg�2S������B�-}��V �u}�7`L�)+�#�@����f�-��r�E���r4�*;qu���eޣ3-���a�jŕ�~�}=���e,��j%�s�J`�%֮��X12�{�������H�V���1yD�w�E�T����V�o�2�z�^���vc�:y���x�*��d�G�7��1����?v��R��{���a!ͦ���} �ܐ�Ę��g��9��a���ZS"q�`@�Do��]2o+�Xb&!y4,���|�?&\��Q��Zb��:���gK���_ujH����f��*\�&}A���e�-�`��yvCY*{���Ei��nik#�p3���JH�ASd�2.�Fߧ��NpT�u���ZX�Y�ݙ��5�bG��V������=�����x�����0�/"����FY>IU=�Te��[+�Bm6��*��F]=���ݔ6��&)�]���2	9Л�#o(���|!ќ�aI�X��|N�i���eF�dYW��0��.x�Ú��7����6kl7u"tW�s1�cSc�u�k����c7���v�-w�<���J�.�Ы//
GW�\�:I�Z���V�C:����T�n+	R{�P�]����6�Բ����]4���[�w,N����FƜ~CW5�y7	��VC�ϙ�n;rZU�s��x�2S]�۹�W0xT�߀���1�9�ŀJ�ϗ�OPAa�1�,���A�ֲŉ��-��)Z����bf�[��*9O(Dc�"�z�3X?�2�h���N^؜��)�d.֧FCq����r�O��*��FXn|{e�ϭ�c���`ۯ�'�>;>&Zȯ�`_ɆE�v��/�Yo��$\0<9���E�	JSO�'a��6�@L�-!:���j�������K	���
�|���!M�t������x�sߴ:�6��
oi6��	��#X3L�_n���E�LoH�����i��I�HS�
\b�u�9�#��ݳkZ�,W3JN�4����*�bvW0��;������>�3������A$��m���.���[��g�S�D/�;�}��ҺkA]+֢��)V�R���h�u����zI�m!�O����w�����D^_�g�����`�Nz|��Yӈ�0J�FS &�lH�燲��$��4#;�T'��P�R;'��&T�d/���k6t���5-�#���F����f�I#Pp�6�����}�(YD?�e����k�q,rEc�Hƹ���{F�-�]D�{��K��}�g�sJ�b�ɡN�1��;�׍���k� ��+�=G$�ٰRZ�jɄ�{��7��u��߻��n�t�Hf�JA������_�2/�(F�r��a���3J�r4K����K��b$|T�K�Py���2T�iDC̶�ɳ_�����l�vYg�M��c��^��Hem�N�+�wc	�.�hG���_��(|b^��t���)����E�]�.�U4�G������dį�Um�,�팡����`�e��d��c�V�]���w��8#W�e��Z������f4��
���陡u_?/���{�GV�}��_��cӱ���� �]�T�M�"�,1���\L��id�\uf��tS���ܗt���u�*o��\9�P�%��������j{>o��D���N�g>�0�bk�[�����|;Um��D��� oݨ�U�Y����*FS�ِ��䣹ΰPe�����XmAW0b��h����p�f����_��^f9c�D��֕6�=X�˜�&C�Q��-����`��@lvn��mH���e�JY'vOR�/+y螲^ԃJ���q���;^o�W��"�)���Mٸ��yٌ�+�od�����/�v�"w�?����� ���MR>�`�,��k��G@L-#j���u���<�8|�à%���[�u�㤎F̮?��b=�U�g��J���<�V+�������}�]
�:�T���:�#_�8��9�X�9!}��-r��"�55 Ʋ9i���x�&$�Z2���%��`'��B��p��r�_��/b��'���TC^b-�Q�1i��&	�me��j�In��9at�� ���\#O�}!����}G#�aEQx�|�2�� �`�} &����\Y��47b��f��4��
V-^�fr܌.�'V},��8��S��:�3�|C�{y���O���X����><����v��Ej;Hʀ�1�D%^0���~�v5L�Zd :�&�~ ���^�'����rTI��$�?W!�<�����2��ֆ��zݚƨ�NƬۄ=��N��j��[�,q�Z�m4 ��U��@Y��Ϸ����k���Ï!}��Hww���.S ��f���2݆d�lc�]V����mO���9��b�?��c���F�O��7� �OF|�ܐ���1%��a��7�8�n*��@���8���@�:�U���ԝ���Cbo2��3 e����m\1�6��d�O^������哫c�V9+�cz�L�\�W#��C�Ѫ�Ӄgm�'�}�j)���6�{��]P�
����N��U��Du�|���i�a�L������A0�nR����5R�
���;#I�"�:W1���i�v�pC������h�ρ�����v㫉�Mq�\Q1k|�d���դ�q'o�~�O
��tyq�R�{��E�M
�:iZ� f�V��?1rpv�E�P��������sN��C&�
�w���p�g1�E���ƨ���
�j2�79��@̿ ��s�t�0�_���U͋�. 6kY�z޾_8���NO�!�(�u���3?jj&��Gt[���Hbw�)�V�g�5Vܘ�I�o�U��1�kBH����娱�td��C@�	��6Gr����]3�#0���c�ݣ�<Ϲ�u6��y<������u'A��=�R˂#b��.g,�8li�h�O?����`1m�V����A�-�ZvV�*0@l�qΒJ���)}�˖[vu���@��Ij����L2RJ���83Ձ��6��PHV&�N��6��^dӍ�"��}4�X��_��) I'�#C����ŰӀ؞��XVd]Y��T�)N��@,z���������P�}F#���@쓔V)S�g��6H	�Y(ʙ���6(���6��i�R/�t��Ń�
;~ �J��iFj`Z�76,ݞj���̀$��bu}�8��j`����9t�UƖ�m����@�Ż˼��#�{�n	E��<}]������[@l�:_�d�V��(~E�7#r+��J������6σ(_{��># R�Tf���d�t(�N�%eǝ���!��>j3�M���KTrB�/�&�_���n�fe����Sp���=]���usW�~r7��,�HG�~pZ�[),Y�%:��AH[�8�Mc��b�d¿�����#��<������DMJ�`O����xꉏT�[�J�rr��8λ�P;"���L�k��30b�rE�����B�l��'����ުS_��8�f rU�k��2X/s������#XD��\���E��"����������Ů�c�ܪ���W3$�r��;�yA���h0�du��~�<ͻ�	�m
"��G��Kw!��`����0��K�0]�Y��=���Z���ᙛ���̤"�f�f�o(u�F,��?r,����-��Yu<�OH����Dˮ�[����`9�@0q��>����$ز=���&2��R�X�	���h���-iBg���_��P�nZ���ڟ^�Ox��W��'^3sr�u0��N"�0���M��R|�Kb�Z��Fe�c�h��:�7���Lr2�Gw��	X}����{ۑuq{�^��׸ߦg1�n�;����(���U����4� ���z��[/l�(�e����Y���͊%����NId��J�sc?����jeO'���MS 1�����w�׶�<jb�};}��e��/��_Ih�{�����|fɪ�D����$� �n��,�c~}V��U��08���d>(�s�!���Х�w���}��U��-՝Q��"�.5�2��W��Q�d����5b�F����P�t�0�r���uD��^8�/!L���4L��W6�S�2?:/�d� 3�l,e]9}fP��-��lyy�>|p�w&_�n8ἳ��b�9P^�BQ����	����ܨ�7���`�j`��8���7nZJK�<G�,\��,���ه��J�Ӣr4�3>�_)˶=ϭo�&��VH �����SÐ@��# ��J�<�A���($k��Z*�C�l1u������t&׮g�SV��~3�v���Ǖ��o _�p��wϦ^��P����\���3��CYl:i�VME��KkB��$��P�o�_T�I��^v3)���C��Q͍?�m�$��Hb�B��<��1��k���?�9A������3�S@,�C
��I���2i%�������~��67{ã��F�
�����Є�d��A��c�x���! f�yS�x�rk_��B�3-���'�b��4z�uxH��ï�7��P�n���'M�7/A��d�ϥ�i���kD=���ƥ��� E��ɸe=f	r����zn�7�#���u=ó�0|u�/e�(�g+k�9}���3����m�֑l�ވz�q�Mm;6�E�A��?,4�[��rE!1@L��2֬$ǺW�����4�z�=���]�`o���	�w�3`�>۹5(��^���}e�������P)�RrP��w�{@ލ������o�AR�\�uo���η
#P�Ĵ�L*�)�J������n���6����="��^ƛ�Y�ؿ� �/��eџ]iK�S|�o�,�(,�����~�n	�[Hqp��U͡[�Y���X�[:���	t64���M~�3E7�F������䭯�x5�n?�e��h�x��믦�We�X����@�Le�KB��'s(~���Y�8��k���Z�R��C1kZ�݌3�3����KZS��}6֪o�o�|�- a��u�}E�5���^WF~�2��0�U��H���D:�28U��mn�ȱ�����J��?-���|�_�����C,�}iË���
������K�I4ogT�Y �K4��韬�	ɴ�,�VcF�6���ͥs�n�^�|o���*�}_e}=��OV!��tL~;����^{\o��νs�ҫ7�__=�܀��/i�xn��ꤾ(�Yz�d���GM	�ɪ�e��l׫�>��S Ѩ>�9��Y�;�����o�3�{�|�]D2K���������Y#�ڕ��ލ:6?BjѫX[g�g�ۇqj�w�1��n�J��40�gZ���eg!�[�\WJb�gV���<{0���Y�_�֙aOS'�O�ً�:{����[6]9��2]2י6|i�<Ր�l��2^b���V�ں����{�A������+�-��[��^e$�ȍ�2�̞W.���QnR֢���"G�95�_-����P�q����e��@���Cݶ��e�w�pzڤ$�m��V��h��Z��nb�����	���C����iV&
�����f����x�������38��Z9Fu�����m�QK�ɰr���7Ϸt.+�㑋�X�P%����n9'�&l]T��%�¢��f��S(�n�3o���e��X��(�B��h+��iARZ%�䣷Z�t����i��m+v����Ś9~���Hͫ� ���kZ����2�A�T��d�{��^AA�1�&ӥ��*���3
%^��lF�i=��-��l�a�rsd5<Z&��~�Ԑ�x�<R�ˈq��
��H��Jӕ��[!��,�˓�^W1�1c�S�JQ�9���>y���|�L�P5�/�ٵ��oY���z٠7;��uqu���@��K�A���׼��#d�=�O�E2+
�C䗕�)�C�}�A<�k
�P���7�!�6����-�L3��jnU�翙X(��Ko7�"5~����@?�ǯ�-qyP�iu���viã�#3��Ly�?L����'vϠ�������������|��٨��ك�6k^8���W���6d�2�u�	��?��W�h��>�m+En�?7Tf��9))�RnDW�>j>��:�����t�Ȇ�'^;6ωUJ�r������d�Ч`T���\���],!��o�>��܁�m�Fb��vP�Q⸜5��DR��6Dv�R�P욍6 ��"��;�Ҍi1���S�ݢ��v��P��]Y= ��SNw���~�z�C�k���5qE��i��]�U��H8&	���	�l�UGH�C�*B^sS��ȖD�S�%�����B�$���^�E���˺Q������1�7��){6�&@l+bV7+�*�:�^酨y{���ÄՋV_/��{��DM�nh^^x�⏿<�l�P��)�){<Q�1���UP�_�)���{����*f^���9�$���ٞb�Sy��_v��\r�H��h�+����F��'B<yyk�P�qe"Z��$��Io5�t�ML��\����CCR<�uO�R���|�fÍ�|̂9�@�B7=B��{�� �\�]�W�ƪ�	M�����O�,T�0x���u�8���3Q��'@L����{�����8����{�+��@L�(�D�)��=�����=�b F��J>�LE�f{@�LP.I�Ĭ
��Z"n�����B~�FJb;ޥ}�f]��0R�0�Hj��������������O��;��:@̏<��I�Tǵn�T��h�Aw ����gd�i�0im;���zIGM��&Fo��A�29���q�`&�>������S�<�#^���R�AZb���(Lh���eT� `�F�F@R�[D		A	$%��;�A/� ��n���A�S��=�gfg��3��}�#�Ha�b�ޟ�8X��F�q�*�H�*�8T���Y�e��#����zF&Yi4n���H��a�_M�{�T���ȭ�ŀ����81����Riӵ�'��������'4��{�v�����/cr���27U����O?`_����I�W��_3>|��uM :�ʟ���1~>/g�Wo����0�+��_�Wz���J�#�$	Y����3|&c��rx��?��1�?�_��e��3nvSv��f����T>���vQ̓'3�a����"��� ��FaAT��{�˴�E3+b��{^F�V,/�N�"��-������q�l2���Fu�����XT$�3O~�/Q�5^QÚE]k��ڶ_NP?��/*\�J$��'��w���3��N���zT-$?��7��s챚��^r�CA�����ۑ���ƾ�9q[f�������}�/���nYc;����v"n��ll=��[ڠ6��>��,Q��;¹�y'�e��Zd��������!�˾��¸�n���mdGm�5t5�CC�c�l$��tm�Č��2�����m��o��W�5�N�jw�������׋�O��=�6�2`���bd�<�S{q�b�}Wh/�ό�q-���4��F@��_�!�jl$v+$R�`��sb��4�\���gj?�0�S���B�����mrR,,gB."�N�L��\ufo�:g�a������f;��un_r�Z�B�h��ZB��s���U�|�pG�e���������oFa�YL1��'��W]0Al'�#��OY�~�`[z�l��Č�͇m��t|>GO��=����4�"W0}��I�c�8�! ���Y��'�`�W�����_�V��]�<=vr���K��1]a����)���:Y=nm�A{vJ�7	���{�ߚ,�LT�����&�!&ڤB�#�v�?�[�Z�n#�t�bd������\����~�B�&�In���2�Z����eSټ�B�2!��5s���1]$A��:։�O�7]\Bkӹ)��Kn�w�v}>����>4u�i8B��<� Db0?�{��ʄ#�5Rb,�'�,���s�������!&j�~e�������Ӛ��`�=7Ģر�%}�n�9�}�!��F1��&�X�1���dX\%y������F��[�����Ky�.�s5�t6��q�/Ζ||4Jkݐ���
1�:񊫅�r�6f�����Ԧm�1�����da���qhi^���)A,3�J��T'�IrQy�rV�����"��O,4=�p�	����(1�0B��:��6ec�4[�t��
Cr�r��r��HnN��E�g�M@̆$3�&��[���Ŷ/�)�����>:Yq�����4J�nu�r��LM�\�؛]�.c��܂X3�Ԭ��B��׼���Q�ta3��z��)��~��D^�8���J�*E�%l�����!l?��B�3&GJڣ�F�@!GUB� �"�������/|��`�?efȨb�*�4���腎:й$K &����%oIUv	���Z���aĂ"�p��>W�k�F����Aߠ�ۂ>�#n�rC�2Z��9�f�lC�����
�gN��읚�C��B���yw���O�8�}nۧ[��s\~ ��a����Brb�U�v{�;~a�ދ�S�e�<$K%r�����
�.m�V�X�F�́�1vߗOQŲ��(@��\�*�&���F���K`L��!�^���2|�s�heE��j>ݝb�پ���y�r�:����W�{N!��%�R@���˔hsF���.�Z��7�/�FJ'\?�1MB��?�hVRZ`�����2�|��bq~k�,���_�z���jqi��-�hL3��hvo�Sn�MB��� �ک��r���t�W�ʲ�<wY�!vx���G��^1�p<Q�o��/���!��9h{�u�u�����1����O�1*,�v�o��HG��L�CL��*���wh����Wޙ~zT[j��Cvi͔���R"p��{��\�.0��;$~���SM��4s��M�_��V�(�qc'�#!vE�A��[����{��*�"bY/۩�܌}{�Q��'}��=���2ӌO'u�lk��J"�f���E��������ޞ�SJ�?�fEa��H��u��WFu6xM&}^I���3�݃]���/x���ԗ��oC�]�v<Nq�����Bd�nw�����E��"ϛ��ٿ	�׳�]nAl'�Řʹ"�>��{і:�(D�;��j��������W	��c�Jy�1]s���V���@^�SA��l��]��l���Y�b.�\P^̣@@l	�Bc�B��'nd��z��� vզXב���@��͒�ؾ���X�P��+�'f����A
K��ZC�7P�0u���^�5?����:�<�F�Q�Y�nrYD�8��IC�ۥ�W~Fj��2�B�}>͈����]zx^�]�!��j�ݩǆ�^ѕ;�����$� �R���J��[A���w�u�G?(?�1X���/?��[�I�k���gt���{�d1�x���+R+K�V������;;�q}��ȻK=b�t~:�%�����&���cY��N��3��d�y��`�L��w��ce|�X�cW`��Ӂ���O��� �Q�C?�G�г�l>0�O@��g�SQ'�ܥ�����oW��\��F��<���/=�M��~1�n;��[wP	�v��?��=���xq�Dv�z=��T�U���P�Q)�|���GX"���8�q�����'�媅o�w]���U�6w���2���!z2=��TIR�@��A�m�D�����Ҡ��(+�b�O�Ui?8��z^�����bE�t��z�������֝8�ؓ�QV�4I�zҨ��E[�aI$k�]�3��t�@�&M�iNl)>��w�	�H��G��Z7Xb�!�$%��8�i������7.�G�	���%���о��������w�۱�l����p�v�WXh�\FJob~��J��_/��߸"�8�2u@�WOãN3꠵&�e���"O�
 v�1�1�P��A%$�Wp�o1�����39�b|�ڕ?�w�>�ػm�Ө�>(O���|\c#9gP���T�ߦ�,Ǡ�Zf]Y?�CA??Ę;n�]0a�Ϲ��韻4B,�{����q�c��E�>^,��#�����-��USx��c ���f�r�F��Y:⫻U�\	��|TSC0n�{oF*W�)տ͇�Qޔ�~hn̋�N�� s��2!����W
$�;�
fGEɸ�c�A,Ʒ��q9zV�]t~��TW��&�N����X�`�K]�%�ෆ���͐��MS�{yL�XJt[_��!��u��bM��ߓ, ?���1i��/���x�����4a�"���j_N�&���0�n�JW�X�˄)��yN�Is�(;޹�a&״����axJ�T>f�ۗ��Ƈ͌�,���\�<�VB8`J	b!�=Xz'#JY�\�<,�F��c�")1r�l�^�3��
]�@Qb����o�s���ޭ�ʏ�!V�Ľb�(2na��z9���,bo�0Sbw?C7|%;6��c"����b���컃f�c?�l��dS��>��(��d�e�H}�6���|1�Dj���t��Y/��|�
�5�K�X�����Eڛ�,*f잖�ÌK��t�K�3��NNd�$��n�A��=�9�#�њ��]]K��A31ĺI���OJ��ѧ��~���S�����\���f%�!�oh!v���iLASԀ�t����6E����M����4ekjΐ�-S�1�$-6�F������ϙjA����r�|&'��@��Kz�cb/�Z��Q�y�p�Z�b);-k�Pz(��A G��\9�bAwE�Y���|�^�QZ�!�P(l� 1�!�n�����,de���(�˝�_Ҿ~#�s�J6�#�Eb�����\ף�`���hG�1�� ���(&]�V�p�R5v���)(B0J�w�QU,)l%U�Ă�Q��W���,O�Er���n�8�8fN���;�Q3�J��\�A;�j�h�3��|Hۻ���rbXd�+�x�i�x�(D�0W~�l��.UŃG�C���t�z�d1�9����0.C��=�����{�P.7b��'(�i��=�=�V�9��OKAl� �8��[n)�f%>k�
�/&�U~�5�ƳS<��4�Ms��i��O���'_��Ŭ�G�#��B�X�����aF�31\��v(Ğ۬U?�|�A}�s.�+����	1JR��eR�F���B�U��?@�GI�R�{`���e��k)�X��$I�e�E�8�_F_�O���k{�k���z�E������Sͤ�P�'N���}kd�b�6z��S��>�ˬD(O4@�㒶�n@�>��u��M_�[�:�nc�������$�_�,"ڧ#boZ�:�k���.��y�2Ã�������jK8�B	�)��7!�s�U���隄�5A�U-��V"��]c=ܕE�xa�X��-ǣ���̨G�+i?���n)�JPc���B,p�e>ޫ�����8����7I�!�vg��C9��V�ۯ-W�P#�[bTÁ.��Ѫn�u���.����S�6�.
G�iqUmK�x��j#+�F� ����-Y��)(������6���5��]Y�Ȫ����C�CMY�Q�C�q<�}��۷��!����hf*��bp.���t�.=��B%����~f��Ê���I���M}'��DD�x�9�G8��Q��z[�9>A��t�On1���%��T�>�'�
���D�Cs} �8�i0��艈n��<�F���X�����{�S]�`dt�#���_^�����x�a�E���?�X�������e����E[nwT$-!�b�o�����Y-w���}W��e�%�Fqc'I��}�H�Z�BGb�.Ą����(.X%C��Ki�xbr�!vI\�#<��5���`����ti�v{J�5j���P��?h1��V�������RAUq��R fo���%'ҙ�ЕTo���2[�1*�5\�֚�J�p��Z��\�R��`��-�R3?���v���iuļ�\1�to4�I���|��eu�1�1�*��sz���*�Eil%��%!Vm�IҫN2�+,S�����b���B)܊��淜?��󢥯0B�U������O�lԚ�\F�!����ܨ��Ý�Q��vj���t��p�;fٺw���YSx��6�ɮ-�P,:�k0?rV���V�ڃ�u��>i6k���7f)���";�Z��a��M:��W6���1�k�S=^��u\Ig����>+B\s���~��R��3ɷ?��!6��'����k��0�Oy�-{;m%X�Y�����c?�NDc4�Z9��t�^�x��ؔ�C�3]��Kh��M�:Gz����6������&�Ã�gx�;�'�wBLu��#<�_
����s�7C��b�X܋=p!C��4�3��YR����k�[��G�9�\~BL�NNZN�u��G�����Sk����㑊�
��c~�ga{�1m�xe��7q�Ĺ*Њ����B�-�c��A�E�^���.V_�1��sj<h���UT �(PRRA�;		�F�K:$������N)��9 -%�ҍ���{f͚Y��72�ͅM� [ހ�⯺�J��[}$����|Dq��?�_Ц��,�}9�cL�F� _����2�6~}ȹ�U$���)x��z�hjl<��U���+Ê�������Y��r�!�O7,�f@�х'v�q�-�K��~j��VN�4�u?vg�.�=9E���>���ʝ
T�������N����]�ɽ�}#G��9�utTf�F�����\���O!W���P�����A�������������6��P���D�sl3��Y��{�ǹ�͖)��#1�1�y ��>�aY�ڥ�OUЧxͽ���K� ���?�>��o���[�	��z��sAEϩ���g<�|dc�[�=P"!YP栚�^����c���w�ÌT�������c�US%0��iO%t�zr�mֲ��9���2i�R^�k��mZ/!�D�ih���X��m�'�Ѓ��G_.3N��R�邲�c�S���^���S��N{zJjD֟4&
�ٷW�=���V�I��&�	��\��	s����%�q��1��G�;#��t���
n��<�	_^��Y����O*���2]R�U� G�����S��V���X��g,6�.�U��B[����5��;�	'U���E	����w��:?:�]�ʁ�z�g�pmq�{$^�b�*��<o!���!!�'�N���E�.���j��2�Κ5����r=��DBK�m�tF�K��KSW�:�R�a�B��|��F���i,���-�K��sД2���#c��y3v�2���
���TL�:��4��#�v���t�;j��C���Q����K�k3�\���l9������?CJƃ*ڐsnǒ��F����Q�ؑ�P���9�\�+o�%����2L��B���>B9�z�}m����q��r�6Zn�~��M�����7�i�!W�϶�؃(�8~�?�2�=�Хr]��¯0�#cƼY[��NT��� �uؕ���H����<pe}E�r&�1'�tI�q���\>���{�9�i�}��w?��c�}K�W�{��ǒu�.�\MD9�,�,TI�?9��w^�.��
�^c��	��_�B��h�H4;ڔJ�MՑ	���Z��C/�<���*�7�}��p��r�
f�u�$�_�IJ�V1�cE��&�K&�#���V�A�ş@ȭ��1[T�pu�c5����9��U�.Q%��؄��l�
�� w�,A�+�,0ȟ�V`v�i'�&��n]�S��)|�g����8�ۅ&b��e�}�L�+������&&�ɻ�l�1��5ʠ�L�9��8d��d�PwC�з[4,�[�ї`�.���[=��Y�S�������8U��$�j!�_!��9nS�;A1��N�QT��|rr#^�G�#�I�F^
�b?�RZ ��iK���F�����f#��Ӧ����$��4���r����ۏ�]ւ\;�nP��@�w�4g�Q��E���QE�IшEp��Σ���51�+@n:��c�5-R��h��"Y�w�%�x��Jַ'�T��"\R��b��ANm�3�e�U��!)��sI��5�u|ԭ
��|�p9�#��*t ��E��_�>�V���6LQ��c�'`��ZC��<����\j��
��h /��Zi�m���W�k� 'J��ki��Ԗ��j�MJڟrV͒#��z�����i�(l��sB�5e���˞5u�!�ɇ���a�o�w��f�6�c�[+����P�]��^LD߬D풪d��
�#�����p�-�|��;�C.S�s�r<�!saрG;�[�r��T��3R{o+v��Sl�m�@��b�Q��93>ͮʳ�=�J��*�0%����łR�1]����r|_,>�_��Ռ^�����@���'��f�wL豣oq^����Z��<�%Ã�����/���yI���& �Q��z�_�$�E���a0�$�\��c~��Gk��/B��j'A�l���<�Z5��a�eN>�U�-�X�N���b�PIX�75�H�ls��>7gT�@C����W��\����>�:do*Uݖ������.�K�r�q/lp�/��q���J����\�]����v_�!�^�w[�y�� �rj���i.ߚ!5\{8�irF��|���&,���*ߞ�"!W-�<Gj(O�ӓ~�����z� rY"�%�zVI�qY�)��{�k$�a:EH��c�wU��ǜ��u%�[e&�Еb�C
��J��M�v��JX~S���n�a[a\9,����b���1e��_��@.N���N(�C��y� ����u�u�y4n������=�/��U�6�-|������ZѮk�u�!G���})ؚ���ޜq)���$r%÷��4*Yɟ�<u��h��e������ڦ��Ľ ���Å����!���J�1������t9���h0��-��u5�mV��%֕.��5�ǋ�5_߹�e��Sp�.=r �-9c���z����tϢr׹���[��M�ʼA��؍kP�2w�h
9��f���5���P��S|�B�J�ܿ���2OȈaN�q"7�(o1�/�	/�0��yK9��"�!���,�o�q%k��������ծ!3�93Ј�p�K�7v7c�9��r��\9ʶ���W����fhĐ��(�"5�@l�De��[��Ȇ��Vˁf�T�R�k��/tg�X�%����q��C,�u���@N~1#�/G����aD��| �rTʟ{��(i�v�G��92�D�����~���QW���j�>.A_���Us~���x}��Ą�[�E
r�-#��)�hy_B�&�k+G�!7/?U"Q��&�ui�s���fȱ�'#u�Kw��4��n����@.g��)��ᾙն��D�!�?C<39��@���~�-����t� L�>OV7�K9B���|��5�Y��+��� �?ӈ�#�=b�!'+�!��wKt�硎�(�������[@�3D\�y$w�luF�^����7�@��&���~y�瓼_��E�����?�6e�̓����]=+�mH�O�7��H�v�Jm[�
Y��;�u=��J����kz���E;�����R�EA�m�P�����+R�d����?�Y���b��0W�q����r������5:"S�˷���?<Ѕ\o��q��xR���u���
��K�2�SrlѲ<�Te��vd�\dA�C/IT���f��I�֟��s�.��[��@{I� �͞-�^
�d�eI�j�7�[�q1��y���Z#U(��,B��n����~X�]+9�#�9�dH/�	=� ��{��<�#wD�_r'A��rr�Z.ӱ�)�ř'�g���\쐛y<Yx��\ňI?=��|��7��s�;�u*��k[�/h�{3�����*�L��b��Yu{���4�.���
T�oX"��z�����6CNx3��� ��Fz}�k��YĲ��6ڭun���.�O�Bn��[��ꂪԟ�R~�}��C�"�#��R)!�a';�;������r�bL�n�.�+YE�ӑ����AN����hܨ�������F�lʝ����B�(�&;�{�c���yfnZ��x{M+&4��dbTY�O�!��~�"B�{84�H[��!�J>��Ņ��R�؞��D��M�C�?c~���px�����`]�Qȩ���!j�����{|<������\����r�}Ί���atM6L5���Y�c|�b�`c�R���Kȡ������f�K�U{!�4��9��
ʗ.��bV��Y���!�K$L��<�Ww�t7'�v�K�#�v���o":�I�Y��Xl!gS�����T��5��k/��]�U��-t���M����V,��kb�����<K�2�Ȳ�_�/�E-(��� �_�!��y^���쑎�9/��7�)�FJ��3��>�	����K(�k����ϰh����@�)�Ŕ{bJ�ⱊ�`䲖]����Q/�%�ɘ�/@3_�Wc=D��x�����H��*n�p�i�b�7v���lE��@N���S�]��u��-|�$]*qy��2}9MhQ��Ѡ�L\f媺:r�P�;*���l.u�&""kh9� WЈ�+fP��!�8��֠�r����&�+]����������C.3��d�k��C����XC���}\����@���i�����CYL�	9���n�s[��8�bF�U^=�9�4��٩��~��m��Xơ�՟/D�e�Ri��޶�l��%m�@�D&���FZa��x�3�IZ-*��9�L3�~���̺?���C)B9}�qy~���1z6b�����OE�!�h�4ș�f��=.�6�:m�r�E72��w0�<��F��y=nIA�'�wMVM�̥��AyVT��U���R�:��2��	������Ҝ��~i�{Q��h1CN��M^H�����N������bY ��H5>�a��e�HW��k���9�tG	6)\���;���9DN� �D��X �ÎYR��]^H��kKrѩ�A�~*�U�{&��Ν5���5W�z1~����e$���cE�r|1�8e-x��	���m���FC�uzD�i�	�J5�E�� .�P$�ZZ�m?��5��n3�J��s��#7��:m�%&�$��Iӧ�1�=�UMsn0^dA�L/vn��8o�ܟ>3]�A%�v�St׮Q��;!�j�㝝8�\�<�c-�\P�bbGViai�����2z���m%͘�
��*BY���|rz��ت��y��\U>���]��{Q(�ǹ��>��M6~1�xe	���h%Y)vUd���{V�S!�x}��!>�U|�iomr��ɐ��/��ڦY[�t�|d��s$r�wvFbª���b�Z5Wr-͆��������V����G��?�}N3�(�������hB�Er'�.�;��F��~z|�U�Q�K��vD4^�h8��=�������B+��6�L��H,�<=S�a�þ��C�$~������z�wȥ�	a��7�>��0E=�*S�\�P��i��L���U�N��� ���RL[8��.5q[���g�i!7[�D�]�4D-�==s<-�ar����_/i%��$6{%�R�c*A.��ڝ�m�7a�m�H�\/�_��8y�*��]����o���w-
��������j��zq�!W�,_�b��4zq�O
�r�I�s�6��>��z{�??�������l����N�~�r[�{���ӎ2�Z[��I8��`��c�{��r=#����}?�䙉���$i�yʗ/�%��5!�3]p��%��B���}!�%E2��ף$�q2���{CN��Bw��"�9I�_����x9�%\~�WWs�,f��+��
R]�GN�]򳰽?uV�l\�ʨ��K�S=�M�ǭ��"g\��;`��\��v��A=��Ji�E�$K�-��5�I&�y�#b�4�zm2��&'u�%�Z��+�o����D�r./�����J��q"�y�gQo�- w����m���D(�����+�7�;�j3~�b�f6�n�_�H-U?��<;h���eP��a��ЍԡA���%E��9t�H7��R�
J����qݙ��q���}������]e7�$�.�wa��tM@'��d�7��L�&��C􏯜{AW��zg0����
���q%�q��I�I%u.Ψ��Y�`����ټ���g��Z�F@��a��}�N���vAO�4e�I�b1'2�gי�\6c&��\����]1�s�V�^\���n�A���m���J~+7�j%�Δ���1m���.�M��P�h٨���`s{�0�(P���Յ��K+w�Ab�Xk4
:���C�^߱!��� ��}��p�?��>�	RJ�4�鮵+E@����s]�U�Gm@��X����a_�@`��1rt��Aq����$�s�fY(xR�	6�XE[[�y���y����a�{�������B;�h�ڬf�-b�����11|F�b�����r��b	��,9���¡7�	�x%�;VgFne�G_���ʅ�!�� d�,�J�=��Y�e�"T�� &ۚ�>�~F���x��,YJ��X�@�Nl�F*'@M�{�|)�j���8oM̱ˊ�O��g�)�56i��ew��S�U!�ôu+'�Kw{��FoǓF�ƙRM'bOȖᓋ�?�s��m�@�uYA�m�1��>�/��j�s��ݾJ+������o)ͮ�/3	��j \�qS�J�=ь�f��$!��d��4�tN�KA�t�Rd���(;ءd[�4�n���Ѥ�5�:�	ltE�a:0R���*�f9k֗�ؗ�L��S�qKs�q`!��o�A�QmO�r�J`�n,�a�S ��)��/#��r����/2?�}	b�[͖�=t,�������ƃX�uaȹ�I�J�γdAle6O����C|�8��W/�{�2����2��ZE++&��k/Q�#'1��g�s�%����S{P��$�?�MDS���%4x%�����C��t$�\b�#����٨O�G��Al$�ѓ������� �SU�-i�;��Wi��@}���6fI���B�=�9��Ρ��h�}>EaP�� 1��NP�(��I���9�ɐ΂"�-w$W�"��b\ <��>f>�11рuM�qń��8%�%�C�[8� &�D�ϳ���j:�s��2�M��b��1�϶]"�k�>��$pm�����(�2�\{����w�gw)�A���b��M��~vÆ[��3u�3�K��_#�DKŕ�?q���)rb�D�Ҟa�蝱6�>���?���Ö~2�T��\6���ث�\��^!o{�q��d1$��i1T�M2db�%���X��K�|��&
���#��|	����a����]Q� ���c�9O/O��*t�Yr��@��:�{�[��}3�C_P��:���Q�j�8x̷a4�������d11�U验y͝�U�P�*�����gN�J��ݞ��)�b(�_�X��`2Wr~p��JxbWj;�s�<�=�&;�S["H]틎�2b%|�ˤR�����N>lU����WF��].Z־�s<� F��9<�>��B�=�*���)�<X��
�ʚ��D%=^�a�/���Ȋ#�?,�1}Z]�>�)ܧ��4~2�/�*j�"��6���fZG�5��.��U�0BhK�����Xql7:iF:�kUܛ3��ຸA�n5y��++�w�OfĬp[s�S�2�l���4��<��c֌o��i��+���E����V��Q�s�	"�~)O��Wz�#��W���02ѿmq����BQ�i:^\ݞET��ug����YƑ�1����~��Kao�tQ��T�"�=������|1���OM��b��?�������D(W�\����i�	ߪ��f������8oSwY.k�OT���#��9�m3�d���R���&r4ʆ�ѐ~g{��)>��@�.@�Ϭ�ZM��Z̉ bqCC�%�
���(��GOݣ�@l)���+�(z�!?t��F�	b�M�d��I\%��2BJ�S�5@̽�SO��F�a|Ks�Hj8,�4�ƨ+�z,���i]֓�l�ݽ�AL�(B��ݦKe8B%�i�ƚ��d���o���
�VU8U*����x�;���_���5X��F������v��*�w�7�QV]�,3'��q<�<{9��Უz��N#�|{_�"�P�]5�U%��$�x����{Y��C��7��W��~KS�['���=Ǔ���S��}��Ğ��H�� ��?�Y`rQ�����"��f��gvX��{ޡ�W4X�&>1�*�S=��J�~�K�p׃��"�~�.q�⦮0#��˝t��y���TQ����	G�!�/]A,���w��%>�`��a�F������F��j��mU[�0��?��M�9�7�%���N��E|M�����F�fW�L�;�{�nF΃�&���!��\2�1��7�{�ۗ=np'v�U�X�,��&qFb �J�ù@ub��4u\�!)�&�Ue�u�!' �32���45ƬES���sez=�����T�r�O4#r�����;��X״I� �7z�����PC��?f���QkzTc7�7ݡ�ŗS�	�e����P�[��}w+[���1V"Q����yĻ7b������l�,�
��	kFZ~%J��Ԉ��3��ާ��iD[�\�Qb2?���ϳ8}��MS�R�4�)(����1���u�hy��+s���q�|	��f���X�m��Ʊ��>�]o1��S�S����61w�↠: ���θAǢ�غ�;�M���%_	_3Utbd9�w��
�]����K/x��]�Yw��{,AL���c`7���O]�����d�
��&>X�B#<��F�������˶~c����!A})�
8hY�\���g V=�	����[�0�9�^9��İ�J��-V�|&�0PyC*�vAL7WLAUa�>����g*Q�4�ici���z��$�g�'��Zy'`߹m�PU�\�xʍs1��J6
�A�C�kk��N�3˞��k��GT��S��&���I^�|�v ���Hc��ñv��)���y��t�1��x6${횛sO�S�xZV>I:����`a�D Ҕ�JQ�`�ʉ 6sp��{�l�O�6F�ֺ���Y�0�?0��`��?�1�I̧ m�ݶ�g ?핱
́O���]����1�2�W��v�a�7H䕺���A�H`�3���Jz�ܑ��"^�tľ6�<��f�6Ѣ=�9[1dAŤ�r�ߝu�1���b;G@L齟5�ꋖ=���7oIB���Y�Ƙ.3c����7�96O]�U�@�-v�
9� ��$�E '[j)Fb��B7�T�ĵ�<n]Z��� �p�@�)�AG"/����ބ��*���L�q���gib���$}�nуX��\��CcV�w4�xsNJ���2�hLX�����d:�*d$�]�
�c'�����Y�XZ���j���f��wgb��\��7�0��C\@���ʤ�6�̾e{lǘ��t�`��U�x�aKP�չ.Mv-*{�C���WO�/�o_�y�p�S���G��\��`���m�CƇG��'���A$D"n��_N��G^j�G�g���wf�/�V���������FV[>o&�X��Ks0�_�Qm|�x��FOG��yˇ��X][�>����j��Y��y������f��5�E$%;�&	LCy7:�룳u����^a�b�bN^�t�${Q������'������x8�0�)O�ؾ���N��'&��(𿮮�B&���6���K"�d�X�oD�}�_��AL���h&���g�1���QY�����x������W_�{6
��K2�D^��t6\72l_��Xs��4ƛ���Lȶ`�U�_�\AL�Z	��ʴ��[��8�W�̎ ���B�Ñ�>k5���/ݰvbmL����f*9}؉OƢGY/'75�o�N�;F'\��r���𸢫�m_#�]w���F�-Lf޷mx�Z}�Ĳ��K)Zv�[�q�4�T������Ro���6J�Ʋ3�{�Ĉ�S�My���|�������>rf��q�����y��z/̌�
�˜��\e3Q��NҜ�NFi�<�q�����'���~��,���.�(e�0<b{����0�ݯz�Z�+�)��� V�BirS��Гm��@I`���6��Ď|��� �q] �!�j=�g���7�,2�5>��B�ڰh�6��ˊ� �Ҁ�����5�vם/PIh�NO�#��d�f9�_�y���~�q5��M4*��Ytc7�Xr��"��-
i�������[w����9���ᖃXM(���Y�G���v��q�?|�i2'���c�5w��_=zu����Ϻ����ek;��2�
�XШ��!/�\v2!*�y]O{<�Y��S��P��x���N�=���KE���5�>V���#�R�l3�,��_!�Cz�(��G��e�}#������	&�C�M"�������{K�~�Om����.;�@��R`��z.��Ȝ����r���O&3,�l`��Qs��Т��@�~d�1"I�N�3n�x�'�P�����XKz�w!e�lax���&Tg����C��Y��]�L��[,1�WD�����z� dS�g���@�&�i�y:Fd�-w��EV_s�uo�Xfm�M0��An�Fv�����7����n��P�v�D7����yI(Ib��i�Ũy��d�WN�鐽�@�3���G�΅#�����8�* Vɣ: x]�6����-�&��� v������M��W䡪,X�5�&�`:�4a�Z��e�c�qg��0t���Q5b��y�Ɲ�4���/�����߼�3��'Sc���Dg��GF�|go�7Z��!��1�3*X0)a�I��}���<�\�Yc�^(N�UgH��4�[�bW	b��
�ry��e���Ѱ��e	S&��ܯ<�s�_��foG'�b���fU��������eg�AlEZ���7��������FVKh%0��l|$twJ�2��۴�Fkl�u��=�cQ&�j~��]�b��G�����Tp����=A�v��6��2�T�~��:����S[�9�(�S�g��z�=���|�珲��ic$V]h�ۊu��@)���Õ�W-֭��qN��?��>.|~ɉF�4�=�*)�bK����Rc�Lpbo���
ALΉ�����%���]���b.ks�H}7���������~Sf��>#g���(��e�]j�q�e1������k��
�odģn�"8 &�E����9w�L�� �B�7��"��a|�O����,f5�b�rQツR[*��3ٚ�p� ��G&�>�̎��.��d^��ĞJ�̗>{H���mm܍Ԯ��Uf�Y9a��]�RRh��,/�b�{�d"e�0����n[�m:�&ր��JCOO�<�����(Qh 67��	�#=��{�VW�)�<�l�����7�����\����˃�	+��4�[,��P��V��r�����K�H�Y(���!���$W���x`�|���v��	k�5�8���������XZ���v���D
I�P�)8��� 6�E}ucn!�����.zJb����Vh���ePh�a�KJ	iA�[Y$�)%Ρ[R������	�A�I?�Yg��v߿�ܿ�y<]�>��ﶞf���T�2/>&�0�
��<F�g�3y� 
_H���~ݙ;�{�Y�.��ckF�qKh++'݀3�y�l``���FV�[��C�-{{��/�'	���%�2��>����7r���^FvkB�@̬�k]B^ك��:�;�gX$EĢ�6�-B�h,���C���"As�&θH!3�eW�9�������)٩�zz��M?B�������{LZ;{K���	Cݛ�F�hpV���Z1��P|��0�ݯ�>�(bṷBbVH���g�
�7�v�-���(.mi>�z��3^�_oq��
���DKR���G��7.���| �=ؕ�o:j�٤�9b6�sLb�Z�e��;rl�u�\�~u��i� :%���'>HSތ���΅3!��#A�=j��JM|��'p),�d|��?���.!��ј�$r~t���2�m��XĿZ6@P�%L����V�����G$���zt;�7�9�1dA�����Ӈ��!��P�^{4ء\p�;����.�˧:c�N~�a���9\��*#n��@��bg����$�������6�bkoeU&OYܒu���`��2�g��CT���K��)X��1A�Ltf������B�x�>��]8#�m"ϲv�/��9-��21��.����X�7�e�ٞ�Ղ���d,W�
�ynSq_��F\İ���X���zO�`�a��@�u��z�����$=�ƈ]_Lbĥ�cG\?�f&�m������MA�S3�z��ː��&�X<�+_b��8���1
��[S�u�j#���nm����S��o��c�Uv$3R�UIff<c��wi�|�O��b���<��,D�?�g�o���8��T��|�|_������id99CW)y+}V���~���s�y !S��
��#���<[B8�,�=٨bi�Q��w�e�'�=�1h������%;,?4�^m��N��$�$��"Cw���.��0G��i	bKT�T���%<�����x)�gCF2{1z�ը{�4ǀ�)���5�A88�rs��8i�+��G|1�O�0���x��2��3/%;N���R��&Q���ş�T��l v�U�Z��\���D��bJ��*�i�苑iÂ�S�X����Iٸ�f����1���� �������Ud��)-��*��V�A�-6��V�IA�%E�kY�P�6�@E;�x?T���Hl�́XH��'ɼ	m���A˙�]�G� 6K�j�?� ��y|�]eOt?���<A��nbbnTo:����G���y�`~L�_�l�7�?ä�y�Xo�����/r�A���"�>����_,{��{�ɳє�BD�;�O��:���oT��&10MVeix���s��=�zI��|�jC�-$��@,�d�2a�2?3��4CW5�B5���hi���%�YIe��$��~ b���D���G;�0��[	Ai�e�3��~�}�g�>�C2���al�b���XZ�M�u9F��geCg����%�=�G�=E�o8@lB3�Fe}�Bݞo52x��ʻ� � )��<\�y����f2]n<"Ą����4�4�Z�7�.�����i��vb=����4��k�1�=��֒/>=W��&p��gb���{����������r��A�F�!�%c	ͺY)G��G"��W� vl+H���Rx�N�1�$h�x��^cW;}���G1�B�m��a��K2�m�,����ِ���!�wsR���n�s^���^��L?1�\{��h�����!��9�Bg V�!��Fr�A%|t�x�n�
bC�JC���Vq�b�wX�vO8��AlX�>�n��̫;���+��?��9_��]��QE����7uu��K.�T �_�z����äl��[?A�l� ����ȗ�/�4z����� f�ݔw��mo �j�.ޙ�b�z��+^�*sjr,���rP�qC�9����L���I!��E�h�� �Q�)"GF
�K�Kj�7��m6��u]y81�xRp_�!_ʚ:�YZe<��E$��fX,�Gt��J�(A��Z����qZ:���zS��s�����4�J�HK��Z� V���K�uv��t2&9y�hĚ����*�2�b�OK�J��I���;w��tc�Q�j$I��6�X��1��z��H��e��HAL���S��9|�1�ׁ��%����X��>�\�I�8'{�SwK��(~<m`6���AW�Ӡ�Rw[���>����^����4����Ć ��y�{�f$}��c:m�%@���_Zȸ�>���:��/#X����5v��/��c�#�� r�J|�xH�b�i�~]�)��Y�O�E<�T$@,��C����t-�I�G��PNs�l�l�Z3\Ś�/���ߠ�l��#j�Sl��h�!-ⲛ��Q fA�2����vjO^�jIF@j��2Ϋ}o��m6��|T����qپ]c�;i"-8ͷ��e|<��o��� s�\]a�4�%l�@��3�Ĥ?����ȕ��qv�x�rf��b'Έ�Ш��J��v}���/ ��OjD|O֓gݓ����X��^Z�i6���K��H{cׂ��n	�]9�!/M��Q
�o����_cW��T�3������l�	��]@l��q�I�Z̨i�F�/^����Ҫ����a&�M$i�#�Y������Á�~@D���o�ܒ� ��~!Y���t�vChxgէ۫@���>ɏ�J��j���#�zc)�@���(^��5�Smӿg�Q�������.wQt�C���4�ɖ�	��)�� ��8w�ܗ�uLS�W%so9a<�B>���hfp?�1R����01ՠ'{���":�-���� �1�O�?ܷ�N��v<�8W����8�<���_%��A���1d��Oڟf�b��\�W�����ËD�-)�(�*��d��p^D�ئ�g��	mmM6��xF���V.�q�sߣ����������R�0�)ŏ�"��̔@T����=��m��%��wӜE��������y\���<�0�X��cRF�<<�g�4�b�w��'�2n+��!�P��SM���`�0�COg:��J7�x�
��	���b�Rl-I�M7D���1c���>���m��8�lLA�	�����%�z����})ؖ�aĶ���ބak�)JH0(d<�P�b��w��rtĘpF����_S!}1����D�h:Rst��p��7Db��?t�)�k-�z�����Ny�p_g���J�Re�7.k���;4>շ�� ����N�;��*Xu�ҏ%����|�{�1�	m~���r�F1y��=ߛ�������,�e6A"��38��n�����A�����*5n��<�U��|lR��OFt�-1gI ���p��O#.jV)���>Rh/´��S��&ZAS)��Cg�t�^S:���0�9�b靄�U��[t�8�N�!�����2kn��y��</^�J��sك��+=��H)J%S�T=No�rH57��#6�!�0xq�FO�B)�ZM�_��o[�$�ދ�ǉ�M�fz�IlMu��u
��ksi�z��[Ƣ?l堀ذ��J��(�Aur��%�a����~��+��Ef�kjS�@��qdl�X�.ak#�*YmҐ�:�����F��Dx�X���{^����5^b�C�)�I�ӷ��6�e���͎.Y�몵��������Z� V�5,�W�6r��!wK�[�u������]��}�|�9팵`�3�_bN����'K�)�:h���͋@l7�|���Ŝ��)�njm.��/E�9V�}3�i��J�1.g��ݟ����*����uRU�f�,�e��T8�l���P�7[�x�!���D~�,2�3�)��_� �e�������"S���-^֞�Ai�bQO&,v�m�C�3l(A�c�,�l-��xb?���U��aP%�2u�g$-���KvM��qc�HF��8��w��Z+�]�s����sWw��
�Z[^B#�����"U�J�@�8�U��0D�����znA�o+��8���G���ܹ�"�(�q惤+�#����f�8��`=!L�3w*6�v��b	���s��r������R� %�7^�Rե�i�����Y��� y�����.mj9<�&�6�iUH�m�"5J#�{N�b�a��e%$�y?i�|�tS��5����M+i��_3��I��f4|���:Y����VMB���"��pX�Ć�H��d���j�z#�-* ?j���"�X�n���M���>���1�*�UT�@x��S %�����#N�M�03{ר	����2�0�P.�X'b�	�ޠ�ʢ��8��=������F)�r�u�<�G�^z�c����NW�V���`E<MhM{z�ی��y�ٽ ��8P��R��ys���q�h�Ç<����*6Q����X�`1�$mCf#���'Z�w�#��ވV����e�F�<���>��6,HA�_5�+�w�G�3�@�JV��,z��/���5W�RO���U����e�j/��b��D#1B��<t~�4�*��*�[jF�f׵c{�r�q Ll��&[�Qǳ�Ģ�3�d
�	V�~ȫ�p��4 ����;�N��w&���������Y���¡���wv�ş��I�?3�b?�v*���Y���yO�}UY�j������������u�"�,0�bt"&��C���o<($L7�yM@�0����T�V�`j�'\JD}�Xl^���ͪHpiI4"�1�O7u�w������2}~-�(��/c�<�
i`�A��R�c��`ӗ�Og����-�p�p���W�,b�E�?�̓s�<ލ0��Z!�_c�u�m��ؔS�M\�I�,�-�p���2T�*P�zHNKA�^8̀͙�8Ml�n�z�V:�,L��u4�qX�ĩ����`F���X��7z���DXW�T���A
����ucU�v��J�[EG���]��k�r���Аks@B�'�����(�PVc���e4rB��F"��ރ f{W'pp4��p�r:ruH�5�_v�<���о��/$S{q����<��C8�CBY0I�jw���/��5v�[̨���c��xqF�c⟜���Ġ�;������2���Φa#�f~Y��6ї��ج�+�$�"�×6��㮵���#�Yud�����M��o� 3����ڰo�����~�Q���
gݐZ72�2��v�?Z�H��f������G�]�|z'���;D;�}��,�|��/>͸�F#�{��<fV�!�9��Vw��i�u��]��߿NU��?n�&W��%} 1ڊ��̔3�`=G}�������<�l�d@\����!�>AV
+��t���\=7�A��s��(��4lr��7[��&�'�?�}�_��&���z;�N��99�>�e5�I�f�� ��ޞy����Q����,!�d�]\2�+�NEeB���KcU:墱ځ*C��kʌK�%�%{�/�X���@��3�5O%�1B���iA�S$���U�L��w��bϷ	�Z·<X53�uo<�H�����۔��\2�������B���(���~]6� �?Ӷ)�h���uPx� `^�DJ��N�n�[@�C�.��n�;�D���vov������3�ӈn7L*R��]��ꏝ]i�?�����&�`�1&K�:${���nT�:��Z���<~��@�B�㓳0b0M�B�2j�(2GN�"��|���_Q頙�H��@�e��w�+H vEJ^.ˈ�8�k6$����7�0�/M���{#5S�����4t�֡���S�G#��n%��r� /�Q���1�%;T*�(���n��:��=�d f��^��X�z�I�p��_����s��io����#f��1�B��lvi���H��4o~<��k���k5��h��p���]F<�)lۿo�D�[��2��Y���V��a��i�i�X �^)y�G>&���e�-�߭�?�4Z���bJ����9ܽ܀ں:���
�vXTw��`gM�m��ŀ!6���ܠ��`}�D�,�IS
=?QN�W�CE�.d=]1Vז;�}����)N���� v���|��M�у��,F+���7v�A�X2�+�YdX�lJ�]���X�z�Y)"Ƙ�ʰ�n��.� �iJ�=���*���PS���{%�	b�B���/^��ŝ�a�x�ؙ!s�/���Ϗdҡ���A��>f�����k)q����a�x��y���I#��n��1�(��IW}6?h��k����� �T֐0p�Ni-?�0���b��<�,�9�+�/�p�3���X��Fd���-�^+NA����2�@��i��`8�A,f���݈�� ����'�mO�U0W0Mv�Gb1��\���BK)h}ψ(0A�EZǵ�����m�AҢ&N�bξ�l���i��3�Ux� G�fw����;/m�GXs�gľ��W�o��ŝٙ�b���Y4�m嶘�Ĝa�D'��T�X���g�ø����',�m~�>6�,W&p����Uf�b�h��d9c�9.���TC, ���Sn���O��{ksf��Xb�@L�:6Q����l�pD�`݃�頼���$�!qC�^�ث�D��я+	@��I��B��������~hlY0��7�G��-�=��Z f᳂G�D��,3i~0�������0����o�;"H�=�fOl��+�X���b1��_ԟ�����gi��AL]��"ҁ�Q����?�w]��Ć�E��K�SB5�m���ًm@����ˑR������z)U��
���� !<M��[�%�vO-�A�cwA󲕎gY��\ƫ����?����e،����Et�j�'9�w ��>I���e���b�r�Gi's b	+�jD���*H2}����_A���K��#�t�ࡽ�����v�>_��ܒ���L�G�1���n�ʙ���&���Ju�v��r׾a�#(��$htm{�V����ap����~�ϫp�د�s�zu54�>��b1$,~�)C}�?��Y�eO
�5r���M��+�)�u���0���z~����!�A��y,�%�Z,��?o|}���!��o��;50���G٩���d����F���<�� 1_����ׯ̧ܴ�O�3�/A��|�y?$�uZ�y�� �d��èDHB��X��#��MQqAL�=9'�F��:�8��.��ݽ�A��%�C�ؔ�l�
 �~��=�K�H�J|+O�� &r��uM�3ƈ��#�ހ<m� ���}�䓇d�[I6���L�;���2����O˄Upb,�&���ɓ'��AT�u��tԠ�!b/���k��*�F%�p�-�|����VaYOs���b��_�u Ƣ+<�=&]^ݞzq��lb-�DC$ƍ+�qV��ᦱh
�}@l��G̅��#�S���ȟS�4_�ڽ�ng��30� 5��g9g��;$K崮ӰWAئ�q< 6����'��O?7�$�Lk2b}���8��Y���V�k��c ��r�V�?ۻ�M��5m9�(��u���M�҂��ۡS� 9��Y�ছ�+��9��3�8 �R�d}�{h9g%��V���5�HA�G5�K0D�y�!�ە��(��)�w�<�,��������ޢ��<�95ӕ�l��)����NO
O�6�$5
�
���%��� �,Ǖ<@��[��V�&��e��=�������p0�q	�y6
b�n�H������u~�y]*V f��,|m�	�)�:�־�� ��/��I���^9����&���U���d�Z8J�K,^�����;l+�:�y�a�t:�L?<@ V�J�`�ez�
��Ơ}�}l�� 6�FQ�����V��V�v����Ʒ�JH��u�*n��F��@}7Y��1=�*N��v-���JBĆ�$��m��+f�v���>6$�X���.�������,4�p&����eӚFG��^�ŔB���Ĉ�8�ئ��b�\�=�!�k1���.���(�%����b0q�l�p�oI-i䎠�,)"� �:���Y��s��%��/�I,P1k�	���o��^�7�li1��-[���qc�9��[�E ��j{F�k�r���oxW�|�!���v�G���4G�������1*	d��nl�X��D�nWҼ�C ���[�{$�--�k�['� 1���Rm� �Ԫ����9σCs�~�����;��LIr�餗� ��`B�q��FyѼ]8��0�( bk�Y5��!�EU�<�HG5&A�fq��y����"�CÜa���p�sY��\nQ<!�E�-�`���L/�i5��o���B� &oJ߾,|��O�{1�{�Xq�
��^IZ|9��L.���r�=(;Ė�E�2���tڙ�P���skmAl������j4�Ǉ�i�L3�v�P���9���⑅{���>L�*o2[�����6����XH��'�V��~�rs�,=/�m����ê�.9���K��" ��Z�ߗ~֧�-nOp�=X@,ޠ������C|_����rVj�3�EW�a�Z�EVp�v7���1��饓�R�-�Ӳ��(#�/�K@���{�rCv��oY�d龂7G| V���:�s1�=��Ѱ�4 �ɦ��b��k��\v���a���o�{�*<a�mv�G�Ǡ��biVA�{u"?�o٬��%Uv���@l��[���k�nT^�Fi��]C_f�/x O �x�JJ���b��xC�y0���ӟ�Ӹ��,@���LB�"�P��/c���Vs����ŝM�Ih|�b����bZPO������V�H��x���� �I�|6��"�Ac����Į]����!�zQ�������A�i�� �t�h�](��qR����5<WbA���p�u36W�V���߀$G e^�4���l�|��tof[�Q�w�By�w��(uu��y~	byEc|�LՌ�gK���jy� &e�_"���[���b���z��mMR��~V�X�Wt����������#�^ZD�.��G�i��5�MJ�&���_c���
b��ӷ����+r�,p9A*� fX��&�<������Pp �^Zb�ة(^�$��RL�H.sEg�h����1�x�^�xY�W/�:b3Vv���標�IO/+�A,lݹ���PQZ�!f�������L��RAƺ]�����Bo1���̴����c�zJK�d�bd�~\�Y_�&9!�'��5��� �70���&��l7ӦClbޛ1������~�����;,���b��Ǒ:�i�I�V�=���@,��R�d����L�T(�9�<t�haU���d�ڰ%�z�l��vq����\������Iꇞ��L/��=�6��u�n�4C-�N��#����Ҋ�.d̾���%
�ĸ"�01��!V��F��h�c��MK���n��U�z{]�y�db�w�����%���Mz�z ���)M����M�Ǐ��H����WG��pM�C��,�kb��^b��^k���F����$h�CA��䙅�<�k1��pr2/z��<��2����dD:O�C��O#Lrb0�o�#^�b�Y6]L�-����v��r��T�Ѓs�ļS�}]EM��e�* �@��}R�<V��~B�5�O"P^T�x���%X7 �z/|����{t�_/ʱ�X�P1�JR�wl0\ث3D�`O�Y�$;�6:������z��nЂX��[�s�����f������ f��}8w�A�c������Q�حBo��+ܹ�A��Es<%�ux8 �/�K��]�O���7����ӯ�Z<Q+���0�l�m��A��	��'ާf�ŅM�jL��� �9�0yz=���8�PN��-�	�zLI�1/F�����t�s�W��� e�j�2�f�ͥ���J#�E;��r�ey[���|�m[�҉90b�%e5ύ��]�gF�F�6��@L�G+���n�v'��X7J�!3���D��`BdF-+L=�HCz<b��{�:�گ�f~�*��qMd�N �D�T���*��Л�x�X|���(�YF��6_���ڷ�L�A���}�[=�5i��7��VY*#{��G�9�_�y�@��y��	b�����co��fo@lViUY�ń�@K�әT�<#Ĵp?ͭÆ�O �D������&�Y�g����)o�ƌN����A�Z:	/lg\���B��g�b87�f���B�(�� 
��,�C��:����D���$=2w1gV���M���K��"��	K��M�e`5�"b�����Z�lb�ւ����!a�=�B�M�(�& &]�x�T��'-��,�ۃ���Y#w:`�r��Ȕ>vfEg̗�
b�Oj�aW�J$q��)��,ALV=��	��i��[ɵ�T�r=�,5�0U�a}��K�4n��a���|��kGE�
f{=�ic�J�]dD�B(!���kJ3�1��܉�Qm�/�i�qL"KTa�b9Y<[�pYjt��b�S�1$e�a���_ͩ�t�A�� �^,A�������IOi�%��v�Ǒ�S��^w�w��C��'ƫ��I�n4'�a�}P2��I@�6Í]�ˋ�Q'eL�:�S) Ĭj��x\�@�m3Y<Z_ɠ��v����D7�w{\��Yx�� �&^p5�yY������,ap bG�'}o ?_�D�ݘ�t���|���a%���$=��#*Į_<��H�FP̠@9-��_Y�{���Z�(F�Pv;s�o��^~��� �w����S�:�uuI7#?��%Z�0_&]]�>�1Q������XE�q���=(^�pJھn��-�-	y�-7�e[�I$�z�Q7��_�'�yK�2�9H�Is�;σ��ʩ(�;�Z���'��ʑa+)��A�m�n����Q�r5���k�7�9�>��6�C�
���_��l��)��}�d~H�.�bLG�uF�_�؛ɦv*�ᤃX"l���e���a�ո/�����ˬ�c�$�9y���%�q��_[���W�Q��nrR�ĪY�����b�Q��ЁU�m7q8/nI����-�?��>e_h���eX�a�R@�;$AJ�A:$���a� H�4H���t(�J�C`æS���&�̜od�������ZB�k�oY������ɭ�h�0lk��Ʊqe�5�Y��d$ݭq f�+:ܽ-D������cm��bDu���B���Dl��4�U��AL0���nv���:���Un��B;[�U�9�CѧV-���)&���X�GMH�B�$��뻮��տZY
�vU�K��؎D^Q�*�tg���C�,��5��f)�1���Z<�����۳*]�k��?�0���EVǥ�O�|Y���.�T�4"ͮ��F�� F#�Q)�ڗ8\���t������*�����:�zT����iL�i+(r���3m>���#t���\�u��j�z~����8�5!d�</X˷�cj]E�@lp ��Y[H0��| ��P�A��7KJKO���ܦRy��2ċa�$�/����o��Li�j���pYkGg#�g�c�f9�jP<��O_^܉��e�_��{��F{������Q�t3ݑa���>� vK����h`��u������'V�&�+!|���������gw��5:���y�%�����Q�-������{���$��(�\�Q!�� &�r�S���臀��0���|"�J4��!��)jX�Ӊ��1�x����
cS�`�0�6�;�����@l����3�nxe!�����.;�Mˮ�}��A�X�(����zNb�w��8��^B�姲��?��������"�w#O�m���ǿ���}x	b(���ݒ�a>�{��,�Fpp@,0�<� ���Ao�=+i��d̫��ʎ��B"����pyÂ8Q�CE�W��{�o4�OY{Қr)�����\!?�U6�P�
�Yoz+��]�q�'�43���B0��ds!2���Pc3V�����8|g棒ƤI@��.~>d�����*��^�5�鄪����S]XtzaW��m�\io���|C�N�Ҋs6h���2.[�1�@Y�qhn$�Yú�����C����E=[n!��.�p���������!����Ts�P0h�A���/(:�U�򼼅[}��b�^ƞ,Q0Ѹ���G\:�Ifq{ &]ؚ�&'��U���`�ƅ�ר��ԟ�Z�Z	��Vo)�@�Jf;�b|/?>�!�q�p;+�]�42ņZ4���F�o���	Tm�A�+r��30��S��i���	b�۸��<�yT-��IdT�rĊ�c^�_��9�r�`wl�������V�%���R���"�����VL����5v�oOJ��0A�hʕ�c
��ōI�w�؉k!ĐϜK	�/9��5bP	���6|@�cΣg&[�Ń�s�Z�W�� &ѠB�����BJ����9	��mx��]a�v�j4i��E�X�v�X:j��W�H���o�R� F�@!\����%�A��X�M�����""��?���A,,�4�P�n19�ˇ4��&��٤�cj�o�U Vk�b @��}ap/��to-�$�Ė}��o!R2L�ȍ)��@�xA�qp��<$��߳|V�@ͯ�	����������)�b�0@l�_��ϲ�sw`�v��W�9�����l�7�?������2�߬x�n3:N���Z�!���ȗ�����D�Ù旃�l�:�A�C��^�g�h��Vs�{J�'YbK ��ST%�ؗ�mxߠd?�.�\~�ߨg�kXY�Q�Ս���p#��Ϩ��U\����E���'�� �D��f]�	e[�&��a�C�1m���K��֧V2�LY��I��R"�Y�>ؗ�[|=�(����jr����&D����&] ��#���$�ίd$��[���AL���æ� ��
�rs�[ѭ>8�`��c�C���4<N�+$Z�@���v����I9<������{ziKSi��D	xx�8�5�`b׺��P���[�OYkJ~���Pb3a}��˟}���#&�%s׏�,�W��xi�֭t�pl���
�ps�5������&ǜ���g�	b׿�}l���3:K�:�ľ�چb�?�۲�Ԟq��'��� 6�b^��H��+>�c���J�q���@X�Rўj/;�q`�?���r�fiR%/�S�ƛ>F;��1��Gz�ymtpS�������lC�W0]	M�m�jw�~����
b��f�Y�ů�"0���;׼�@l�����Z�Rhk ��5ã�f��-�pBv�&�YM;�j��1m�>�]��������w��{�A잉�����;c	�#!m�Y�5y �]u\�m���ί7�`ʀ��bP����6�;x��ßߡ1��Xŧ!�T_���Mq��u*R2 �ƨ�$��eߝ4>=�^S�.�|Co�ݓ�@��u��D��b�h�n�H�5�&��!��b8 ���R�U���YX���b�$��AX?y�����X�1���M����{��q�s
)�!dVx�U3�l	|0L��؋��&^�KIFFAlgM�k�۰W�6���n)�Zf���}�;�'m�}��p[ f�.�'�e;��DbR���5�H�Η����S��.�'��3�W���rA�cI[B��cP�w�;SG����9 f��<X߉��F�Z���|��.��n�,S�Zr�<��!(;o��X��{�Մt~���]r#�A���|���h�vfɥu�K��k�!�_���|<��e�V�y�T�/�L�v�'ZR��0�&3L�V@�^ k%
���0�L�ɑ<b�ܹ�f<��&�|J�\(OֆA���Mm�dq�
~Џ����Ă�,�S�g��p/I�$n#Jd;N�A��
P����-�d�5��!#҂�~qs�\@���٭!� 1�Ҙ��a���}�[řڕ&_�KA,��Hn�����m�݈Ύ���=|�e�-,��c�����p3!�e�1(�ۂ��!O���CA�8|�����g��]��?�GZ1�M[:XwE.�������l8�Y�0�a��vL<ʆy�,���X��޳ -C/�����v����+;���(����gS��q��U��^Ę�b#<�ݨEAL��8%��48�(�s�Y8�z'$��<��|�GKPf�ތU��)�9�T5��Ge�*���ɀ��B[ų� !�k��t��r��P<��E�t��=�1�i'Y������R�'�
j�-�]��]3� �P�E��A0��\_-�?sn� b��Y����""�7M��)ꎃX%gƵe�D&z���DG�1�2� ֿ�ǳU�S!x2[�I̎1�b��(�m�jã��G�u��My�b�:�g�I�5�:P��K\�,��A�:;��CbFk����槭�� Əj�Ŭ[���i��ԏ��y��(��ɌJ�����&h^��X���O%sd�����U]/]:�*��z̍�̣�����4��	�؈5A���5������Ҿ�F���H��� �;@���������ݎ�w��y��󛡕� f�WfM��"ш/�W�z�F&1��.��]`�ec�:l�t[�m�V�%�J��Q�S���K�as;�0�	<���pa9��2	K��l� b��_Ӝyn�>���n�}0`�u����������bF�S�w}@,J�qf��(Mg��g�R�ӹ�����ԯ�(��cd�՞�R��F�}A9�{�72�ɒ�4U.(�����G�����aBwf���/Qf@,o��:)�{w��+�)'du&�<�;޹S��@C׫߶�Z�{bo�H�2��Sgu�o� ,V��@̼C,�J�";��g0��Tn�b�!Pd%�؞ֵAυ��g8ܺ ����b)��J�����5IL7zQ�o�\mЄoZ�Q�2z-�|�-�5!-�#
��X��/�c����2?�N�i)�-�Ρ2��+.; �ʬ_}P��B=f�z'>f:^�bz������˿V^�U�)����r���/���0&j�C�%_��a�}��M�!�Rq���u�r}s�*��Q�U]a?vų*4�O]<����{��Ă��h�E����7$���<��џ��
�e�
�i���tA�`��5��,l$d==�m(7�0�UG؞X/bp{Q]��p+�-��ża>#��da::�S!Ԥ�"`�ƓL
b�g5r[�
�%����'zU+ۋ@���ƣ�5�1�٥�����z[���L>�^W�7��i^��w���,·?1�9֥�)g�S��������A���~5�6
Z�ymT����B��-�-
b��g%C��1��Lrr��)�R���O�AӃ�O�\�n��\$v'Q.T����O�?���f�٥)�>M.y�T5/���\a?vo��@����\�_�~�c�1�Rr�am7Y�S����r��P, #����#�))!��<��i�&�/[��-���f��eS3���׸Yi_�pbC'��:���F_}�}�-p:�����+���zX's��B��f�f�g b|��5�7��/D7��JSI��+j��D����A�[:��h)� 櫰W�t�S��+su?���b�?3�×%��)��n_��9
3��3�\ǋNн@���	��ވ������4��*��^*�o�r����%��CY<V�������PA�x4�m��C��p�$��ɓ�kA�RW�mM"��܆�s�/�u@Cq*3N2����wi$�P#K��f���dCqR�V��c���Đ��|N�������e>�b�����'���Z��uăE��B~47�Q;����xb�8_�sU��@,'�A'�D釋�kn��S�{e Ƅ�z�1�{���t#wA-)�F-�|Yr������.X_��=��ey�b��l��(�"glg7���/f�@Qϱ�)t�k��%\6Z�쑞�-v���rp��w��G�S����#�*<g��Q+����
�~�/W��o��Yf���cy=�,j+�"����ʍ�%g��/\5�3���f��`�E�bvn�2Mv:t�/=l�Z�U֞P����B@,9��^����J%� m�LkD�H��\�D��Ȭ��{�6tyb��x�hf�9׬�(O=R��0�����B� �n�Bf��V���AL��kUqSV@�{?��U>����T��9�YB�1V�;|��̌�Wڪ\o�g�Y��d99AK#�:�N�/f�_����jp�.M`p`��F�Mv��r<�9֠��ص�l̈́*\�q[���z��m_�7�r����4 ��P��C<��}���C�4�U��|�ǲ~]M��3���������%	^ah�+������ٮ��֪ ���d6��@@���܌f�d�L�W#��0��e_a
�$���.������DR�V �+�a%*T&��r��3���μ�F�wC�Ѳc��/�.�h�O��X�B�@�)�ڔ��6�gub33SPAI�o�z^ȃr���K!�Bx��OvS2�zC�S��_��V��,����C�8�÷�+��b������z޷�ˉ���~�����`����q]���ř�,^�d{�(���������$���aڙ�ck�W�̽���K�FO�+��m#kt�w|_
b�U��1d����f���ďp�.w@������AVb
���@��k� ����{�ɆXw���PF�eb�km������� 	�T��M ���Ҵ��܃N�%����1���5�k�g+��zP��髐�p����Ȕc�9�d�����$v��*�4�l��!�ک��J�a�����'M�h���eXU�@QB)	A�S��[D������	i���+���Q�0r��oo!8Zd�ڊJ�m?"K2��dm!�KL�����+��:��M��>E*x���x`!6պ�>���W"Xd�����b&��w5-_��!�D��\:���(��H�8�_iz�����k�k� �&��W��-��V�\. �l �?@���7��$S1M�4���!Q�:c;�+.MJS�u�C�6�bB�yi�3.�\��D��[R��@��S��^|��̖u�bl�:+�SK��7�<��LV.�F�b�/d��Ҙ�Z���|c��%��˄����a�\ҫ�З�0c����By��ԁ�Zo�GdW���h>f��>ſ�����:��N
e�:�[�auc�6�P59^�j�P񣭐[¥F?����4��m��/˫pOԉ�(��gG���Kr^&1�WH���9t�=�Qo b���ʨ<�c���6Q�T�av$ӗ����	�3�3n��q��~~	�D�3��i&!���(��5ݸw���a�>��#�	���ߨ�f�܌�b����
�Z�M��F)έ`�Sl�أ��/��F��m�q�)д��U����BU�!g��(vU.B�qV%���
5�d�����P*��,�jv?����2w�~�V�f����y�~[\D��R���x�v�5�&x�ZT�gBG�`�gX%?��7#�j[�w6��7Z�oE7�@����a�ʹ�|7�K����7��I�E��H�F�n�՞��ab���;�֠���wkKd\f�?���]oh���}�j,�K��^:d��@��0��S��.h�}��.����c�o�v�����7>AB�#t{�<����M��	�s5l�yO0������˩~3�K�W7Kԗ����@�*&M2�(�pz�柶{����Ֆ`Н�����WI��g5�a7]b�u�l=\bק����x+R��.�$	��hG�5�[T�]��6�e/ODb��!�K�toH4}6��VYn�΢���d�Ŋ2���d�1�'W�%�B��gʱ�!��{\��%�
�I�����r�{��/I".�_ ;tĲ�l$c��}��٧�i1�<�����ɍ�;�h�=9��Cn�E�e���m�i��m�&��T��qv�A&@�C�3%[�^�� �w��u�gݿ�����i���@J����x֪h�=J�,P(i3H;�"�͚%����vk��K�*,f\r��)vGlR��2�sd,巷m6��3�3Oq��.- b2�F(�S����!K�Yai��1S�;J��ٱ:��C$(��i �Ye���"�I-�|πB9�%gO#�he�K�4��
Z�v�@�y�����k��m�2I?��0�Z be����r'1lF�h�����_^1h�5˶ܥ�j�=h�t�Cޜ�0 wS���U����؉��)�@̡>�։�Ar��o�0��w0����aIA��L��k=F#�z�9�$znq�Y㤗^E���� ���u�D���&�˺"?ǯ$��,O�v��4��&�%i>�^�{�	��(x�KwsW���'޽���6cV�ˀ�5�ԯfO�2\Go"%?b��b/�\+�X`��)��}�غ<TԀș|4��~A�;ud�@�Z1b{�����!��ldl/�x� ��iQ;úX��o9���mn�²u1�54WŅ�S��.��P�wK���$##	�8�� ��b��c�� ֳԯ�2�N�S�x���#a�s4+ �&h�k&�2Ӭ��/��,���L��Zg%�f��t�y�1�j����S�ׂ��L��"�����liX�K��F2(��BgyeQ VwWb���)�M��G!�a�#�n �׫��p@�!S5�.2:d������?K�����E'�Wp9(����D�ؿ�̺[jLG9BZ"NĲls�̲�6��#jD�bJ� ���
�F!YPG YY�h�?)ӟ��g֤k4?8�����5V��d/�%���SВ�����】��ZM��@���*�s~�T䯦 ޲vp�Z��c)�������
�a�3�I �4�]&��m��r~ܰ�ԓe��A,<~��o��/�jnE2i�����Pu�qWC0mT�$��m� ��MSWbB����%7p��n% ����z�8��x�4����e�3���z�QIϠum�	Uz0$X�a�eߊ�Kʹ�4J�4�!T*��b�%$Q�=�P��O�I�0���z�6�a!��ܲ^�U't��Hb^0�Qb�M�:�E
�RE@la�12F�T�>�58^��-	2���'�wiz�cW��嵀�a�/ľ�6����K�{�P�4��f�����a��Z���f����}s �^6�ء)�yW7ga�c���*Ry�:�W�9��<T��7C�ʈ~,�#���Z:�[��,C��[�71]�+p��W.��F�
��
�U{D?��r�-�	��1G6~����q�nv���6���.� �g����@����]'}�v�^1��jQ*�~�:���K��h�¢�p��d���Ņ>8��Nzۏ^������G�	K��e" �՘N�y���q�yb|�N�����e&�5��5��˿:IuO��,Y:V8�f��R%& �V��`�m���D�ɇɧ
BD+7�x���J�ˍ�k��.�0��A���#�<��
� _����o1�&Y�b%y��b9������T�"%\�H>�ɽ>����%v�rNR�?k+\H��W��C��!�ً`�;�Fh����ZN��>��8{w��z��Ŷ2y�^"݆�	���wCF>x�ͷ���M
:ے�W7��zК�M�@Sxz*NH�~S_"��[��C�b9��>���9O�������q��w�&�8��`�<k�����=o��b
����U�E��Y<>�%y�JQ��j�
��e��F����.3G��R�Û�����5�ۍ!΢�bq��$_����cبM�ۣ@`?"|���RU'c���|B�}@v�tpL�Jw5�F+Z.�����h��Ey�CJ�m�
^!��������X	�����=����\X6ݜ�Tr\�ј���$�E�h�=Te
�>��;h��e
<�H���{�K�����b��?9�(��+�Ҫ���1Iw|MlU�7�H���h��F��f�|p414��ֱ��D�_0�)?0�u�=A��/XO%lL�{��dF�+��-6�j(�����y�TCP�Bm��<Nq�d᧰�՘�W^�ˍ]��1��6�3|d93��a�����و��f�"�.I�G4#y*c�����T��K9�U������[o_���1����v�	&)�n�������7��s�_�p�	5������m�]�}�MRm��P�9��${��|w��~��&��HE�L�|	S'_9�eMN�3�Xi�B�t=-/�o�e�����"��ANIM�`�����Z�@֩�@��r�������=#W��*���W��/����]�|f�4�b�H��uk�*�x��0n� _�)��K�s^º ��w.���exjx��i����燎@��_�x�o����ԞƱ��L��_�h	�{���l��'����N�����Q�(~���[7��;�mt����p��?)��Ղ�4������B��+�_m�p�K�[ɥ��\����g���k�Ou�N�NP���!+�����)B��i�7�C�K�7�~�X�O�>1��;��UF~�	���
�G�Ŗ@�mo_�*��V>R�~�ɓ�m�7@,.s�yG$�O�A�ǩZI��:�fc;k��:�
�P,l-	 1\%.��g�<hj��h־D&2 1�����,�>p�"�E�cs�ob�V1ю�i�[X�G�գ*�?>�� �R|9Q���0+o�Kl &����/��nW���J��{�D-��m����ۢ��)n:�o���diEk��(��H&������@,��O#��E'�,d����]��z?��,M�ߞ<m���U�&r�o{�Q��"���G6��g�̣׈�J*0at��1۷t+D�蓁��x+�z��M��awm�U��e�T�T7�9A��͹E%(���S�Н�_\�6��<�>~�u`1I��LC"�I�8^�v��R��m<�߻�F;,��8�+ZtX��j�C�\���У�e3I��c�@�L%��̲��(+�]\ςպ�A��_�H�+R�K�#��w��
�����"QQHfs:{���!���+�EF�e�t�hh�im��u��_��o@� �F�m�n�s���+*���}�Hl	M;G�2�&}��p��R��+qD���6�q}�X	)N�3���_b�Oٍ��e����W'_Y�a3)A�[~e�d�J,�7;�x�e`M�)W^��b�3Aӊ�pXY7����IŢ��S��\�ϵU�U�m7�4��IY���vv��t�~XD�`�/�t�L��)%G��n�o�����(�2ltW���!���Y:���9jd�P���9����\a-��6Y+�t�Me�۰���a4�ش�r�>1���a�X�t�t�rf8m�o�n:����
���zؖ�T���]{|��Ȟ��u�c̂'�b�̓u-���Q��&�n�q6��J���/��7����ß��nk���R1����M�HO��iǥ���5����eS�)Q+�cfQi�!���Ab����8MOH��������7�����0�l\�!�u�ۋ��"Z_;���XK��:��!Q3F'< �I��EӋ
+��Ҁ�D��<��b���SC�(@}��v2��Qχ��D)�(�f��YO�,bx��|a���3������0�#S�����y��i~b���q��	���&ԝ�-�4= ���˳ϥ.��L��_�����_������d$��[�<W?��sm;hjƠi턄�4����nE����-���jiA��c��r�k�Q��n��fY�)��̌i��^TG��e�˘����O')�~��掴��z4Q�ǁ�����F��]���%2���M�b=* H^{{8�����#R�X\/"-y|�
�}���S��#�yY�����k���8���j��M���k
�j0�?��E����B�f_h�	=iG�a6��[("!g�	^��o��xN'iRJ�z�`;�\�6) ��&LD���1j�'̿�*���{��ĵ�c짥K-D��'�v�����)��V�lI���f��n�Q��o+B`��l�a� 
.b	�ut�/�.���4	ȑ J�G�����b-3C���x�f�l��DʼY�bs������l�L5-J�fcWW���w��"��,�bD��b��8�sC�JOE5~7{1~-åK��na�g���Ao�����0�(n�p�z�ԛ؎�\��@̷�$:ጁWxe�%�d�.�XìzU���k���8��Q���9ww�����r��^]@u`ό���`�]�@�K(�l��T&��3j��s�1mФE�� �1M�ڐ#'�l���(�zL��2ؠ��q��Wu\�B��0��o%"���8��1�w�L��P:��_�1�DѨ�:Wn3��ϖ�;�{(���6�Z��&,���M�TM6�/׵�v��$��� ��[��I��㓱Jc<��!�װMGQw�a{��k?Ȟ��[Wk瓇Nǲ3�7�~N�8j/rٌ���~�8Qj�f �=�����!l�y�ж��mݟ�81�dc{E����*�+8THն�<��R�S�qv�%��B5�U��xʔ}�c�A�a��e5����VnO��y�;��?���&�2|���Vj}O��v�1C٣��̈́���G~���8�ï
4}�aw+��{�#d*a����ȡCv��zw��0W�5���af�a�M�瑃�fT�O�ق��� 1��� �~�#�}d��5�)a�_f��&��hb2'z���~ $Ee퐳u��>�FA�)Y*5���͵MU!�8�6�څ��`�B c[Y)��u�	�a��v'����)�.��\Z����Zci2��+��k@L�!1��ʌ9��9i �;����?6�@�ynL��y����ݧc͹5�Y$���0������aͼN��)�a��F%̑E�eV�c��T)J��WX��(�8�I�`x�ۯj��m�z��_���HW&�L�3,-����i���o;q����5�ۯ����$lq��ט?�W���KTfr�tk����@vz��fs��I�L_"�)���P�r���6�~t?�V�?T��Q��!A*|��ٍ����f��\-���7`VĠy=C�Ⓖv
C�0P
㒢�~Yq Fvdt$�V �H*i(s�Ӓ$��\TQoz=k0ν�Bd>ɩ2p�-^u�FZ�18?q$n<ͧ�MC���m�۳tE��ۙ�����|�<o�<�u�{�s���bնz�
����`S3��4>e�O����q�YK\㰀���r��>�W��~���]^��@O�>�됮3�p�1߼���)��)j��L��o��4HƟ���b	7&td8X+�?,�'�.:��#��U��x��y����2�������7a�i-�hʜ��@�<�Gr7�Eq�fr���J��q������ۗ^L��]4>�ud2f��¼Sj�ɏ���p��k<@�j���FL��G�Ӎ>�X=��Ő�?��yk�Xi��$����~x���*[��QO5�tc>e}`����o��C�'�@5��c�����A�b�~	��8��f�[�E-�c�����i�7|P�k]$j���c�^��U��2O�R��|��ƴ�H���;D>�%��[L4bM����0HNc���O�����b�R�EG�}��u{�
�뚶��˭�q�nB�J~Y�("�셵A�fJ9��k�Ħ��p*c>z�|�.����Uf$��\�����O& �æ:pܽu)��ܒ����e{���Č�-��W��H����x�~��e����Azgr#Wuc#Lx��XZ}����O�{��?b`�I��/��Ew�����z>�B�'^0��]�w�7�O�M��	�~l�+��/�[��������F�#n�c'!R
d�m fb��������&O�X$��7"��*�9d�i2��;չynQ��j�2h���eXf��a��C�KZJJ:��C������ �% ! ҍ���t7HH���8'�|����lg��Kէ]���5�ƽ{ka�'�`�%jis�0���LluH�s	 �v�܌�C��afR�b%'kRg,�e4EY�����)��+]��>���:ex�d4|��q�pܚ6@LZ�-��"�����"��,�ė�&i�F��^�GD�{�&
�Xр�kN���Lo��١��̽c;�F�M6a�vQ�0ʗ����E# +��Jef��ܚ!լ��A���U��Ҙ]��R �Z�@̺����G�ei�h&��K����⹺,�}?��S?\0��	b���/NM��7���Vo}DP�1���	R�5��X� �t��C3K�CC���-���).�Ke�ak�C#wC��xM�H\�mY��bg��&�*15�?����+�Qbo$�K��L:��n��PN�����>�#�~�,�iS��k ��E�ؕ1�׾L�¹Fͮ1�x���~����k�Ri�Q����Lh����~X�9_���)�c2�2�v<1'��sW�z�%�L�?a畫���?���� bݜ��
���Pr����|c:QCAl��3�G�#�{����ˈ����H��L49Yv7�~��|b6јO��G��ۤ�*��璞�k5���^�;y�zt���N1>���-k�PN��L9#�c�oM{�@̷��Y���U���;�_��͒�H�����\U`tك�A����:Җ,{����c\�H2�����B���TK/��T�3���+�F��:��I��{}�' �%�2i@I#���ȹv�Ĵ�/i��p0Ȏxs���s�&A�z]��\y�fv�ĩ�%/C55��u�%��d�0�p3�^�&V������y��w:�y>�[�-�8$�H�h��J��B(�jQfK�as��
6���=���k�8Q�YYb�����jMTD�4��w�o�,d�Xx�J��m3]�}T:{���q ���i�.)$0�� ���˿�C�=�ՙW��P�,�8c3kzDy�ح������		#��M�\�� 6X�t��Ù����(�7���ɵÅ�I�4�7qd��)
8-����FbW!
��G_�\�b%AL��q`���ufj�|���=k6�v��8^����.���ډUL��<G�8B�q'$�P�V�&�}��z���l���N,^r�qo� �!V�&6q�9q`�9�Q1�׊�K+�������5@��|�zC������~8fi���?�-*a�ʙ�j����q�X_X�<3���I砫��&��� v	.9�͞�`��fE�Ah����]�H�֟���=)R߇��=g-1�dF�P��#�X�����E�@�'Y��\c*��\�<�Q��[C�~��~T٘՚ȉ�� f�!%�&UzB|P�ҩ�?xn#��E]k���I����k��"Z�<�/kc�tA��jI��"�^IIB�{=���Q�	�¶
��F�qE�kYd!w��	�q�����lA���9�&���{_w�")�M632du�NX�L.�>#��(�Z�mLx&�|����}�*�0�M��I�O 6ʹ���%fF���h�g#X0?b�y��T�q�)�r����e�Ħ�
�M��||�U���1�AL�O�Uo����I����k�O�N�ÉmY�Z�p8\�����`��'����R����� f/f)=�A�c/6ط'Dfi �:ѕ﯑���T�u����X���G(N��h1�ˆ�I��s�C*�&aM�-ViUk�q�j���8��S��F3�D��#uX�b�{��&WONĆ��p�b��>��d�v����S���+C{-&g=�镖�#7��bˤQb�è:�؜۩a$�2,�?�~� 1��5"2�AU�v����� �0ʿ��U�R�cdo�́PK�lڳ���?"�d��L~4_��1-�Y�[��p�9S���+�?� ��`���#����VH��@�����wW�B�'.�97+m�;OF�m�^ޏ��p耆�������\���~�k�n��B!�
^>AP�;ZH��pz�j�����W�94IŇѪF�/�دVM b��c�=3^4����u�D��y�e1������4��m�.�M
_�����Gt��V��yU>"�;+#B�7��QCe�t{(x����uͫ�9���t~��&͖����&����=��wS�B���ӊ5V�p���9�zX���Ճ?X7�HI��֚�h�~���fm���ն���H�u�f;=o���'���Um�ֿ�Jzzt�Е�63^o���$CD&$���.��>���|��i��n2�յpEx]㭨�j����O��Oa���� 4�#��_���zhc%W�Ƥ���%���3K���B##z�>���NQR�S+����_��	��n�'<��h��_7k�a��n��gP���U�ϔ�Oc��;9� ^B�N�~�䷴�pG�	s�yi��+�(�$��>UC����=Xט�{�a�������ѓ��p̣�+f����H�6>'*�H���T��5� ��z户����a��j���χ�yQ���W��#kqo���/Ɨ�ڙL���j��
NX[�W���Ê�w�do����|�X���qsD:��=��X�/���;_m��.F���Ӵ14:Rԑ�o*�e�vu7����[w��=?2�C�8���_���u�5����5s�Kd���n����O�	j�4'��p�E��Z�K$�k�	�֌�:
�Rm���SY�T�U�J�Z&��M�q�+�({�wӚ�h�s?���S�)�r�I-� ���aS��oPt+�s2O)� ��d���}_�Ыl������W�
�F�X��������lJ��{���U<����G���Ӽ��"?�^���C��u��^�V�7'6ywE���%z����w3#4��9�ʿ����K��s��8D�z<70���g�����������<6��d�q���˵�(wO1�w��w?\�g�@��2�����%O'��������;n׹�i ����r����z�wȵK����6�ӻ��}�|M|~&ܡ�pa��Vؤ7@���K���V�k��?��r�t
���T�em<�o�>=�����,� �j��X��K[|����dJ�&��0���Ή���?����Ւ���������G~/���w?|�E�Aʶ\MbT����{vݡ�	vs�)�͜��|K���_�2������k)C廮����޲I�]P�[�!g�?�K$�Y����d���Hb���T�q^>[���Z/{J"�~���@�������x�[���KD�(V���o{,Q�X髡پ�7w�dÏk�5�jD-#D�mZ��������'�?l��n�-Ⱥ�'^TZ�x�\�$�(�a��XE�E�wQ��]Qov���W3�ܱ����]��T3:�i�y>"HU��ؔ��<&�p[�򧝄չ�.��F�J�0�m�~��4X�O�0�b3bk����Z�!�X���O+����ӗ�P��� 6���d+R�J�z�_�Q#�B$��-��f��vZu�cM��s�����w]��z�Y�̂�9G_)R$��;�b. ���55����L���ԣm���f�����5)꠹n����+�m-�ç��ɓ�ؓ~1}t&u2��>��ѽz�Ѿ"��N�2���j�Z_�ӧ�8�1�6���ȯZŬr�O�;�oσ���s�R�8�����c�4����=x}%"F�a$�Q�i2I��8�&��e�g&5,�j.M᫕�µ��g����"	& 嗵/�LR��}r�u8����hN��&4�s���t|���7t��u�i%�g�/��LS6b�{�AL{�9���]��p�H
_	���^G�W���������� �F�#�:�ơ�?j���I���7��94o5?D�ꮍ^-x���7�Wmn�K���`MQl6~�]U�� <T�`�n2_�a{e�'�p}ު_��]����������"( ��DDI��3s�%ˀ��e#t��.;���}�-D���{�B@>���36����������NT~���_6����rf;Ƌ"����\����L7������R7�_���wvQ.�nk|o?*��7z*�>�!	�?�P`�S\r� h��o�ɳ���D���~�w��'Ƶ�H��S���l�:>iR �V����E��1��u	�>�
��7���������u��Sf8ʒ�n���,ֿ��{��kv�?�A{�����T��w�}>7�5�m�=4k��_41��߲r�{b��žq���}�sN�Q糱#�z�]���K��Qlp��n��� /��"q�;�rlEs�+��dC|�P�˞�m���ֱ�ȃ�f��'V�ӊU{ 1"�esһ7]@'���x<t�ۮ�]�Sq��@H�o&�������s�=;L��p(�xE�ĳx���f��kf�y�~,"�l���j�� L˗��Wxm�PR<�m�C�kU{���	�C���U,=7X�smK޼�1���8]�|u���۲�i�8gensu ���w�?B*B豢������j��.b�P�c��c翚_���S����j��/�Ò��6(�z����͠u�0��^����=T�P�Mn1%�(�&N	���=։J�o&�ܼk��9���M��P��v�q�g*:���D��.@l(���m���7����ꉉd*>��F^���4C1�}��1�a�V��f��n��lw(�b�U���w���.���~��|�v�VՑp�0cB\a�lF������9%Ӂ�қ����7����'���b��W�6�h>�l�wny�c��yb\����XKӒ�+'i�B���6q����ӘW\ң�7t�Q�*oZ��W3rt/$� i�zA�°�&�4�w�y^�"�S�Ԗg&�-���Z��������-@S��}z�u�C^��@�}A�W-H��7�����N��=z$n��>�;�"��VNMﴚ~��M^!�%��uW�[Ï���i��d�)~f��5|���_-K���d�j�/�A�,o�r�>�rӮ+�]��.݃<�7V�f˼��m��C��n��	2h�^>zS�z�!��%L�� b4�f���f���HrQ�,0�̿��'�Ͱ����q�w��$��,!�@��=<, b~��qn�����o���Vu�O@����!���5NM8��#�]�O��&^�5řM2]"�lb�T�K�,����:M:�ԴT�U �9ޙ:ĕ8ٶ>������ Ę`|.L�K�ЗT��e$�hR�ǟh}C;qs<m���7��)A���BhH$���m[��m��4R�v�׭9^]�i'1.n�~Igb���B��*�u��b��и 6h�o�~	�S��[��s�b�a>�Y�8;�Ml,fI�X���U�:�%h�F��!2�F��Fz^8=0Z���L���b�����a�q�#�M=v�u V�8#��g�%�x�l
1����b;)KfԿ�g��?�Q�l˲��Y�j���x����I\���|#% fG$�xC�U���p��cN��@�S��?�)��J���-R��t��b�7�eY������Ta��] v6���+<.P��ސ��j�4�)�ʜ�M���"c��a�~��pĔ�]k�q�	H��Dn-G����X顟���󶖥���wȦ��� vF��|���)��d�ۤfik��CC'6#hIWzd�ݙ�	b+�&#�k�w0=+b��={��]�A��q��Y���:���č�7��N�i�~5F�>MdUC-�������)�����IP��<4��[�����l��ȋ�^��Kҥ�]9����?���b���.�O:^N(
)���<�<4�'��Hy��hd�+]\k±���:�����0)e�6�75�?�@Ϝ�'���J}g7uR���>�0H�A9�|�!��Y2��&���l9<&;O�nm�����ߪʳ��;-�#N�;[�,*�w������M�������V�+�g�'���s鴋Y��r�1���7�w����B��j>棓B��	�}� |���ٸJBп;� �FK��'D���]|�(=m9k�o/�m�@�;x�i?�,9��c�膡UƧ����;��Q;�.�?2��+�|�OC�����}���d�콕0*N�y1Ok�g�����ECf�XZg���M�R�t ���&�"��!9n$Y�£Ny?�G��	5fU������%��5 A��n/m�� +F��!���A���(i��3^����ʿ����U��ê̤�P���#ao'=����#k����Bb� �R����uR�K8��if��� ��Y9�hIi~�0IG�����@���~��.a(\�>�%lݩ�S���.j>�p���I�׹���kXw,�"���Ytu��bA���#�ݦ}����K�����-+�z�
Jyz�T�3m��P�t�֢���&�"�����l�>��g��� ��aB���-)��x?@���3�1�}
 54�i�Pf|QK/WCM�&b��!��Qi����5�v�@̒d���i��^�s��X���<Ok���y�W �G�+�b�L����J��K�WؘB� �ܤ�S�߱��2w;
-�HĈ�|Q�|��pr�͊p���+j��uH^%�߫Ãv>�O��X�
�`Vv���j����Vr-���	@�'&=��y��*�q�h�e���ͧ��K���]��Z�����M��Μ����Q��[�]�^P,o5&��b�����5�k��n���"'���e���h���eX�i��a��;�AJJ���D�FZ�F���V�ABx%���C������{ƙϽ����ǵ���O��A�l�U"���QRi��0Ng��}���2��"W%�]A�."�my���ln��j>�d��0�Q=V$\\���	��U�$�fjN ��aox�[ �׹��L�G��(��^J=^����qzv�B�7��i�c�ް):A��K��R���b.��ّ&�<��:�ɞ�] �>��W`-�䶰(��և�w��t9�Gu�D1�ſ�{���b���^�dMl>�ַL�~b麆��w��|�{�FEEHgǠb���策Y:I�:�¯t�T���J��Y�Š�6Z�AL%��$�g�S���q��>4W8���{X0�jX"6#�]���Pv?S�9Jwz4Y��e)�����!����)�1���'�l�	C�>��Ȃ�~��5�a�A]�Ʉ�û�͋ ����1%\lB_'��w���Z�b2�g"��{}��DC��09�5Ay��HI�*%v#�T�}bt%Y�l�͆�
{vn�kz=ί� b'��B�'��Sܬ���(�ށ5}�@���=���uT��c� �c� ���<pN@~3>�����&�=���k7�ֶ�U��+��XÓ$:�:IjF2m�$����&O@���S3��ղ��1��2��^��l-���f�I$���AG�ˣzCқ�SM8Rx�b[�]��Q�j��~;���4�"��#�4W�Q( �E�`�J��}4��ܴv6��Y��lcjN1�ಪأ��&
bkmX��מ���KU秹z�r������h�ӂx���3c��R�v��mo9>��M�����%Db�r�iN��Bm�P�D�/A�<A]���AK��VO�c�t�DU�Xf�q'�8*�:�` F�R��s�,�w��������� ��%�`Cϯ<ˉr�|�.�	>j_AH*4E/UȢ��=+����T?Jgo�5�k�٭	$�cA,���e
��8���޾�QH09�9�:����vI;g�Si�����{Hm�m=6���O�F�k���؝{T,g�����Y�%�}^# ���U׉����nKV�R�*|��sM�*���s�g�o}��;Le�i�.�)��_S��j�3Lw�C^���tuKĎ��Bk����S�MR����V���I�������jye�Rp���,��p݄���A�_b��a�����h�Ѿ0����?>�ra�/���<��_�y��SU�A��[�M�����w��C=Q.�I�s��s���c�򤹟�C�BebCqv%iE
TZ�FG|��J�> �De�7������x��gp�=���ʄ}(o9�M4zk\2ӹ����TĢ���Ia	�=�x=�!r�Ě�U�6;�*%]K%j�g�J�@�;���]x9#�@6%�h\�X	�F��en!~Rp����o���b�G��L%m��ٝՒ�Rn�Ư�����b���Ք)�x�]a�(sed9��^�Q�ձ&�y����.m�I��a��������-� �f�zXb���}|�=�V��f]
���_��Y-���W��&bB��1��c�|�W.��6�מ�#2�S�B���7����n��G|�@L���o��~���l~�3G6�$O�3f���j�-'ϐ+��=1 1���}�k��%:!pr������ VŚh��*@H����raxMxXĊB�%�O:��u2I�8(lR]1&��8�S����� ��U8�yb^�fNR֨�4>�����t��g���E�L.����4�įM7�s2-JVE��>��~|֢b��Q6y�+���vUm� �͋+�.|�����U��j_�pZl1����kRW'�um;�@�"T>�D����X��5���K��v�9��/��k"U�5Q�	����j�~�a��m��C\e���7�����ףe)�xO��<���� ���F��s��u#��X�k�@�o�Ś�ΰ�0�pT�[0�Q)�=���Ŧ�V4�:k={b�V�#�ka��b�p;JG�qG;H����ڱ����}t�;F~J �x{��&WT�/�g0P}�9��R_j�a�PёyVOb�K�/�f���?�i=�}�H���:�}�� �������оL�B���>�u�b؉�'�W4X��@��)��4�1�����E�k97.99�_�1�q4��D�{�Ymn�EP������0C�̂�.AlB�]"�1��6��~�{pG���e�Z�H�1��~6PK�CM<qv-�S+�J�1��#��l\f�헝%S�� V�iƍX�ZT~e�Ҷ�J�m���UMO�,�h�S	^J��?~by�S��kS#�-	�c���4�� �Gl�J$IL;{�jIJc�ˀqĈ-�E�5��0sM���$�$L@l�{pK�Y�榟�)}?�4���d�,ս�z�*����&��	b"߇���Ѷ�l�腎���� �y ���s*�?��u�GQ���z#�I,$������5�y�<�E����!���a��1J8�瑉@�ϊ25MbJ�ү�����Y=6��N.a+l���BM߭q�5�Y`�b|���sC5&3VG;O5Z㿃X
�����e������5R�ȥ$ ���u�*����r�9*C�1��X����h�N����d�U���
b�N�����&a�k2	'�C���'~������i2�%ג�Y�wu,�M�����|(Ʃf�1������S�RA���U��`s vOuf�<����?������϶ &��B�ޞ��(zx*}8�w0�nb�D�=E�-�LudH7w�6
�4@�ª���Sq�[��w�W��Q��ۏ�I�P�f���*R�4/�1_�-�;|�%��וV깂�{@, ��8����I���.��b<{��ɑڍɗ�u���
U8e;�,W��>�Pg4�W֙�Fيr�1Fy$�*8����z�n>)M�.�٘$�'��sLd�a���
b9��(6	�}�;)�$�a�/�Ÿ@�g�7/�X��[v��_��8 �ڗq�-���B��� ��H��o ��n��,2��aj��.�:��:����P����m;�P������|_x���QOf��*�������]~\s�����)'��/1���>O�bw�ٔ�0%�Y�j{�k��']�����u�;c�q�t���CRn֯�4�������b�$l�%3���ϧ��A��<I�wԛ���Z�r�T��m|�1�'.e�����Ά����ALV���!�/�
�ç0���B�	��F�긙���Xf5��LvɀXtܓ�<}2w�Eª��h��� F��W���c���}H��(z	biu���{�ְ�w�K([ Fqi�2��)�鶊��}�Z�*����i��^�c����y~lṘ b^����5��G�[ZE�-�RK��A��7i53�d�c���M����e�,W��pH,LƠM��$�Eₘ���L���u�um���@}��W+~���.&�cW���H���b����O�s)V2*�e���71�����7n9\B���uljs 6ԁ����RYu�&-�l'��	�^U���z.�Fa_����a�s3�5�@R�+�`e�u����cK4t�rǊ=b�D�)��������`���g��[�D�o�=�<A��C+��ì?BQ6� ���?ĈV����WŬWRaX)��� �?�^�@b�AsO��Nu�F?�U���&�������-�HRVX��b7q�SQ��'B��[�3��G�@̔{\������L��M������!E�3�@Y=��Sb��>%o��]e�5�mX)��g��Qv��X��̀��9�	�RY:�ͤlck�E]��9�A�)���W���
be�K3U�׫�����龥�Al+��i����n�&%[�� ����9��G�����)�$�p@G�E�jl���Ջ�;�k�=��O�����n斱�Πp���l�`��<�)�oȯ� ֱ�
�ln��(�~xb�� \W�+U�iTſ1�6�y߉_{3��&�y�k�Ԏ��.MN ��Td琭B�����B!�49a���Ho��y�}ޝ�<�v�n�Y��l��hv���P❫Bw�Z�aԕ�p$�V�<DSW��@o���5#�'��<�깲��z����ir�T����E�1d8�n�8 ��i������:u��8�\Æ�T��_��h�XP������d�5ٯdEK���Av+�2�?lA��R��2d?:i�,�d��B���UͲ���S����|��TU�_�2d�f�j(�~1$Ƞm�M]�bƠ��ץP)xZ6?y"��Hؓ\��w�L�֙��[3��� ��(�v����E����2A�Y�_ݧ�.�|^c"�Ĩt��Gx����1A��M��k-�T���v��D����,	��W��/��}S�,��3Y�X��E_S�`<P�����љL���aQ�� ��D���H#Ma:3|��P�]��W����[٧��}o�4;���A6a���ـ�$_(��.�&�+f�?��������z�X��V�᫨�̾##:�2+2I���ռq�L�-�)I��a�W�T [��f9dD���u�ۻ���g�\ۣ̚ʹ����i�=�i���t=t���`�̭�4ct�1��٣v�?��������mc�ehc]�H�5sX��r;Բ[|2����9m�bP|2y��!K���>=�K�^{-�o��m=��{�z�!.��o.���Cd9\���\�r��]qw�Ɇ�~ڦ:۩�%O�����[�W=tE���9yʝ�:z,��<�k���� ���/v d�]�L"��U�yI� Q���
1ܥL�/����A��j�0ć�c]!y�C
)��?V��0Y�/��#���7rgo�X����X��z����]����b�NȢ ��~t� �n�Oghe��b֣����kߋ	<��w�y+1��]�dB�/+��q3�Bcά7w��-�w϶��_c��)۷Xgr}���lZ0jL|&�n0<����������2�a�/���Ci8�]�oY7�X:ZN�س9�F�in-9iT�"�0���?�&@5��?���ɨ^���F����Þt�߬�-,��"��f�PDG���A�N2�m�_2hp�Q�#����r�Q��	
b��ͮ���i/�b>w��n�u �/�V�T�\Ӿd����>d��v+F�e�肒������܈�+ƐU@���ѱ�������8cq�>yȎ�rd��:�,:a O%s?qRy����z��bB��Z��ĥ_��:�����4\��9F���28<4�?4�Pd�ݔ�+U�	����ד�&ND��L.@����J�:=�J�?1�eyR �u,n�!;����p�����pZ��F��pBf鐟��\�a   �  8�{���Xq#�Qj{�!��=��ݔ���b?<�[+�*pl~*��=Tݏ��9	��,z*�	S�g�^*|"]h!���R'ϯ���N���K����?  ֑��>�Y��K���[7}���ae��}���':�����9�ݺ�;R:Tjm����k�ɇ�e>Z�2].��`bR���ο�;p;D̔�E�ד?����*5|�p��������O���'�V��{�7o���?e?�����x���>��5K�W�+;�@��Y��;���x;ab����b�8�#�M�oaLΞ��L���f�]����)b�[��sv���S�"�z��ٶ����x�x{�vj��xU�T~_�:R���=���F�#�����ݑ������\��x�Q�9��4F����#El�}�e���vlxT�Y�׫]��"��EH�g�Sv�wr3����[m}��n����V�V�{{�
�Yqm{0)bi�r��[5��؊�9�l"ELd���Go�_t.�����'x�&����� �+��}��������B>,
V2L3�i	S��כ[s�L
LL)��!v���r���_��_�d��;���_}�����Lr^U�$6����#����2�m_�����'�=�q]��_�v���SCl��t1/���xE7��ά��(~�1m��F# w4t�4��J��Y���4X�   �  "%  h���eS��a$�E�n�V��$���A�[��ii	�nA@��A�,3�ewv�������G
�Z�d5W�*�3�(�����b��_~��N���"��Cl;x����d풯t�L�3���孯�n�F���- ư����O��BIO�e^f&�tH+y*t^@uY�"�.,c�b��i�{0��k<!uQKJ���hbu��6�l�'#A���e6����3�3֮�n\���I��'Ą�û���h�ad�m�nS������^���y�]L7\����L�G�k��Pj�K�[��7tdϡG�R�J�q�[��O����q�Z��pL1d���E]&њC~�7���`�qG��J�?x]�V�F����{-� {��I"J*�c��՗4�����<���'�#(�����+�2+� &O�Tj5�t�B��W}�b?J>gS�a{�B0z��] ��N���%����Я��ʄ4��l�igkN��.�׎eO6��᪔���'�R��q
�~�Z3���Bܹ?�9�4�Jr����8�I�9h ���zl��}�5lK�HA+�M:u���KM� N�7}� f�p�-~�Ĵ�!:J��Z���ĸ���zS�_����B�.��k�14mXq��Ʌ�X{o�k����!�쓘QV��D1os��R-�1Q����O��AN��Cm�*e� �=?�4-�22Hs��$�
oG�i�Җm����E��p���ļ�H���?�eܢW\Ah��A��{7̓���|Qi��Tct�b�~��s�Gx��IgO��a�E���� �ޑ���<�>��2��E�$�MLn-%,�/&i�����؆W����MHc��OG�eB��3�AlֱP�Ķ���*ڂ���4�r���A�yc��_�-0j@l)V�����#K9zU佡�n����P���-��R���(=1-V%ʕ�nc�F���C�v�p ��;�b���KGw��L��-���/��%�!�EKM ��$����J��6�����W�u��O��!χ��Vj�Sd،�ۤ-G�/l_��0�CYɤv���ٖ�
b��G��=�X���j�)��Q�9
�E1�%T�V�`Ϸ���?:���<m5���6�ex4qXO�z����WR��g�׽�� �q�c��+y,�<�[����[���#3YL�MH�ir\�^��h�s���9$�E�F���m^���I2��6�յ�PwtOo�MR�l�%�C3G-ԣm2�N��]���
��I
@{�8���s���"� ����䔁�C��1/�+Zv�"b9"�á�ހ��A��h��b;ҵ�2BU5I�Ws�mg�0*�4��	�[�b2x���.zo�Rn���}���mQ�oC�h�p�a���Km�M(�!����a@̷Ĵg�<¾ɸf��D����kb��8�{7Y�*�I+�M�h�z.��!c|=9���ܛ&�R���?ńV���$���t�~-�n6d��A�6<��L�D}�iџ]���_�O|�1ߣ����}e������0]
_��tk�F��&�
�9)���t`g��.yü�����L3�	�Ք�?�㿐�'�<%��s���p��+t�DK!��"��U���������zʆ=��)�*�}����m�BVǇT��fJ%V��J��������������T����G�{�:�_���1����}�r�V~�� �QY�4ĈH�c�'�H��>�4e\�=�y��٠'zN�
�vO,���bm�S'�7��K,��ե���_��C��uw�늯�|F�v)k$OЂ�6���y�gg����|#
9���<�Ŀ�{�!�Ī�u �f[� n����?���k2��\tƯ�Ewg>j?�X�І�&���mR��O�Qc,O�!ec�S,��]��)S��3��VЊ����,�@�������~�j��h�ʌ�u%_yHa�3�ď�1Uc��ؒӥc�!+}��Z��pNȧɭ��l;�m3r��0{����24�/*�/�0Ҙ���kHb�2�E �?��
�ϛ~��Pj!t�3�)�2�H�J3(EO���麧t�λ�j���a�(�T�p��s�΅o�`��s�_��
�~-ox�⒚�h�[���4�3d�qx�#.�6T� �23x���T:��{*�m~��A���PRx�H�?�*%��{>1��������K.��� ���6zՃ�T�S��s�"������Z��f������M�en��Rm���bu�|������~:�7X�������x�yv�m��q$ǍA�k{�}+�*'@��,�R�f�6&�z�������n��dS�S1��أ5r�"���@�y�0�)�۝e�U)�hJO���&��-�D�\�^����9S1X��x?��Z�S�$Vi%W�6�����Է��X���΁�(Qң���W�O&��Χ���7�G<�T+���[��ۂY�����kÕ./cO�[�2<'�%\1��U̪�}b�h�B�w�a.��1��xCn�
 �ը�w�d�bEdJcV��m^����5�X�Ub�)h�yt�u��د���
[<��
��k�dt� �~3��@c�`�)�4j`��E�
b>R�*�J�d�XH>-�V��1����1�A�4TD� 7��! ����ýB���l� �lVbDs����w�k�체�y4�A��+��xm�d^G�&��*��:�Qj}��nK��7b�~|gb�)�v�|�/O\�<kNKd:�Al��H���°,��hR�C
b��U�L��4B)��r��A�!��}5���*���F��L����aC2�$�9$d��h�,A,
�w��-<�e��o]x�YQk������G��\u��c��a �XKu]��U�?�ޢ���������`�0N�q�XɌ�o�9� K�J��ԾX�f�,|g��Q8	b�N\S���,G�&S	w�K��@��&�}��R	~��T�Բֆ9�����2E)R0�8�����耘tNe��&ұ��wM�ω@l9�`��ʵg9޷#�v9‐e��3��\^4�f��H��n�D�1��w	��_U֘���+�m��XL,�׎�\=�K�(<�["SL��q�+5���yx�b�%��oWwc,hloH��z�6axI�[�Q���2�e�$,�%����rKf�x�"�76�vCK�	ľ���,[m��)P/��_ă�{b��{w7H����bhf5�x�� v���?*,�jh]!������� ��7�deHq���F�9��CC31��$�g��ab�ġ��HEK�	��&oj�ָ�}u�;�YdX��*w~��r��cB�\3�'��>�:r�ߝ��Џ9Nk��D��>n��������~�P�Ğ��R���G���:�����Pf�����l[M����9�����H�K�|}!I�j�Z~;#F &1|/��k��{Wm�,r^O	b�����OƦ�x�'�O�@���b�E�i$�~,g:Nrb��,ŷE<{$ƻԶ�y(;� F(ZZ��չ�;1[�"��}� ��)���	���P�r4MB����j�*���Z���M�Hk��PF�5l��Z?��`��}ϵ�b<o��3U�3�����+8��@�ی͕�x��F*z�1���,��2�z)�o�7�.x�L�$">q}����Z!uI#�tg��	��G] V�_*������7�Nx`��3�!RÍ �=�zS�dm"�dӃ��n'u�����,�|����z�_8��c:.6�w3k�*u�1⅟k�)ϴpr��e�����y[�No8Z�cwjLYFv�uz1����X��/=;�������8ĺ��X}6EJ�6�5��������(*�٘q�PR6.iRkXv�"�	e�<Q~7d���Ҹn���%39�qȜ�����:O�O��+|#�0��qx�@+�rڗ��(6�I�5@LC!���/Zene���m��� �밠g���+��۴F.����4<k��e�-\>�	<|�?��	'�t�?�b䰓�N%�
��%Z�Ŀ�㥤r�b�]i�a�.�u%k�����@�@?�=
M�ԛv��73<-l-��B]���t���{
�8�Ӷv��A���$%)�@<�9P[�ӯ���ĸ ���{���0�]R���OA,{Q}�1-J'[�aq�0i�E�v���R�R-�e;%}r�
-��@�����e��kz~�+�N9�i�0���xń�th��*A�HC�&v�^Ԏ�2�'~��� 1��}�%�r,[r\T�)��J�_x)|h}���Y�)�S�xJds�`1�i2
�q�6x�i�<���jN�H��<䟊]r.��leZ��] ��X]��p.s�uLF�Il�7�p�vG�Mbz��`_br1+������V�� �q�u/��@b�]��7ݶ���m�k)\��k�C��`�����m:�WƖ�<�����W�Dl��{_}�;�A����I��Q��.�����A���&�U|Hb�x�a�Q�����y���D�����>~9��`�l����EIv��	(�8���5S���C`�#�f��|�f�q���f����'S]���%ќ�`,y���t�;e���kVNL0<����1�Xr"�<�$��� ������۝J���u13Y�o�L��8@lh8uT;�ޠ��v�X\�9��b�!�vǯ�	)e�M����I���C��t]ւ��Ȓ �\�������V�R[��Ӌ�� ���kL�q?��,�N��O��bG_�=�CWH�.S��{��S;@k�͗I��7������������bb� �aι��Д�m�XU���6e {��m+y�H^[y��o*���BP�r?R0Fq`~��&��󞠹�9�4�l���u� f<�u�$\���������P	�VܙB�1��81C�d��:,@��ӽK�/�i��v��� �Co+�¦LS�$�F���W�b܅)���8�j����E/�E@�Wm�O�w{��b;~���d�P�:Tx��N/��k�����`����]�iC�(k�߆�nU!b'�a������_-������?�����F&9����{i�鎻ch�7
O\�Z�Ē��?�8_�}o��|k<��b�~y_z*�X��Ό'���o?1j{��o��_�OVR�j&A,�kqh��AE�;������p	�h�u]��0��o�D����ALHb�����[�����rkL����Ҵ�ryS$�z�23�,�-�Xc�<���%E�����}�I�� �@�����fHk^��1�&�FĠ��/���������l$|��J���i��-��儕l�`�"v��k;�����nT��`�dC,!l��Ĥ��9R�8��7�,�mkAf�mḕo��n}}xZ�[:���]+�H-mZ��^��Eقb�R8�z�1>�7[����i�NFD�V��>�аӥAMcb�ϯ*~�Ֆ4I:�F\ǡ��q˂X���k��Ye	)Vy*��� f��V�M�:�a�^�&~��Ns^[,�)M'-�cN�Y���BD 1>�=���R'��P����/{E�@�Qy��A>|IE}e6�,]� FV�Gg�b��x�&�kb_gbj����'������{��v��� $m`hh�)O���$���X1#?�@�d�\̄��������N��脎�ڳ�a�Y�+J{��o1�,r%")���i9��7�c� ����w@_w�m��#�7�,Ĉŋ#3����9��]�w#@��p/�v�!�&R�M�1�G-.��$Q"���e��'�}b9����� v���z�+���vj�;,�����dQ�}�P_sۼ���e� bk�pU��*m�aP�.��;Yk vd�����_^�rFg��ݾ��(�7̽�>*b�c�7{Fk�ԁ�%�`b=����׋h�4��Z�E��_�Z�&�@���j�M1X���!��e�$�SO�Tn:㧂��-��d(��-��A
b��8SN��e۞p{i{�5$�z &K�n��ԫ�n9@��:`���jc<�G� ��F���ȩ' 1X=�]�IJa'��c��P^�GH &�M��j�RC0��#�,i*O~bo��I�/Tqn�}�~�m--����@�sQ��KY�ooNl\V]�@,Ϣ>A؁�Xi{��p��~#6�q*��&?��k"-�'�g#�����T�-	r��穉P�9
o�@�S���;��XWc��o�V��D�t �����
�4
�9�>�f���z���h����# `+ٜ-#{$�JVo��Ȋ���u���rdfd+��蔽
9�8{���2���{>>�yEd}h
ߥ��lǆ�Ԉ�����b6�D=�1:��L�PЂ������J�OR�n�U��gU�u�q��ykœz�M��~������p�4W62/&R9��s�c�bd:���N#�Pj�̥���i�f˕9��;�%�6Z�??�ϭ���V�[ōދ�fa��͟�JF�t*�!׎�j��l.��wsE=����0�a3uė�p���M*.��Y��w�d���f���G�T%���a،N`K�0��2���5:rU�_݈�2�n�u�ܻl�Fȕ�6U����u4��6+�L��9�`2/?K�w8��👱/� ��T�8���R���[�T�x��9���g����M�ޫ�G.�R9�[��>��%���T[��rg&����M�tz�=Y.��vU1�Og���r�ȟ�_���aR��ȣ� GԞ�O���XO��#d�Y�jB�/'@�u�t��܇{�����&ȅ]|���(,�8�G�fO'��+ ��4[���EL�������vVT:����<;gC�r#�|�=\���\�!$�(g��Ul$CZtr��b�e���t���b��Z_�C�y�q�}=�j�қ�2�f{ѻm�C
=���fF�۹�h�.o�f�!���N��#�B�#�N��}�]7���g!�=7�����v�O�y(�'�sn�uy���6>�hb�0��B/�'�O��r�\�b��I~&�"����^a�\�`��#Q��sѴjK��9��d���if,�*anǵ�S"�0�-bQ���-Z-��jK>�����ͫ�%�aCV��j��F�����4�J���j3ߺ��qe�7�?5��k'�.B�����>�w��;����2S}, ]?M�2"~b����Nf����r�"6��G���)*K�c��lW6!���GE!KT�Ӵ���V�B�8��*`�bR�s�h����~1�m���DP�Pχ���Z�c�\ C�PK��d����9�q��r�©xo߀U��}��~�2�e�� ���8��(�������^>���NB�3�Q҆QL/�:��J��_Z�[Z?�֓sx(��%����1���.���Ag��9���2�aMݛw#l�
�hH��_��X3�0
�i��x���9�[a-�����o��)��iC΃o��X)�x���ڣ�u%ܣ��>��s�5��!�˙��w�6A��-_j.]��Ѻ���kZ��J!w��a�����άRփ��u��ȡT��ZQ��A;�����"� '$<��i�^�˗ٿ��DQP9�xD���)-��fk�Z
)�bH�M��|y��:���E?��E/��%�96�L&�G(�����#���d��t�51%:�q	Y�(��9� �I	��k�A�����{s)MbӐC����t�n2Z2{s�q=�)���<P��>�h!��[5��v�E;�!�����|�2r�s_�3�`K�ES�R�֢ђv���e��軏�� �g7��7'T��2��զ�Z��]�ܤu��ZKO�G0��{����ѨCN|�կ��i�s�)]Q<}Q3䊔�WY�>��M
�٥e�{�I$sT��
�����Ё͹��r�lm�2	�v�ӌV��y��M!����K�nqS����i�����7�g8�V:��;�xn�o�Bnĵ �l5eȶ�$�>��ziߩ9/��gJm����W�LE{9��
��tڦ�+�����7�~������9ٚ��K�j��F�ޤ1K?�8!n~�acO�A{;�>�?�	��:�^�B�fG���~����(�-�!lߑ៺�#+�0Z��>��\G���eѡ̃�;y�R)�4�BO �^��S���1�[O�q��k-�%�vŜ��ڇޑ��s�R3��!w���`O���ӯ"�>�w7�rX���t"驦M	Ꜵu�*�rO�&'�YurZl�-m5�r��~�1E�l���繘n#���J�9l�i;G�J�A�;�d�5' r-�ϼ���ڐ�-�'f)(
�!�+e~o�yܩ8�rS��b���p��m��]Y;���o?����r���̓�a<�򃔶�ǘ��I{p�4b�,M��Y.s�!.��JB�g{M�+�S�۔�-�_�ŭc�W ���c]+�[��6�Fa��Q� �E8
�3��
������^<����a�8Gq��0�A,�0��C�i,ɪ��j2���(����d9������C��\��S�5��ʻ�ǌ�ά��	n�-�\�=N[µ�X[T��a��_<�t^ab��f�x;ޚ��1�n�[h��jk��Z�w6Y+|�O���>��>�ыy�Tu¿��L~rJv���D$�Nƽ�o׌O=���v	څH�Tg����p�r���+��0���k�g<��G�ۈDk����7�<�mڎU�������d���˧����Y��!wP�t����b_e׏����AN�(mq��W����)!Y��s'�r�"e��v�U�VA�h��\Ƚ�/�$������P'aL��n��� �b�}T������	���$8�O">eo�Z_��2�W���U!�@��S�-E:mž�C.�럷e���*��ڐ�D��O��܀�_&�����:��$�d��Q���܌�����z�8���r�~�����4uR�7_�dM�q�b��*�2&��zsp.����3"�nC�����[��7�O�~0={!�d�Sё��AZ�e<p����&>�Q��E3Қ��!TZ]��)'!W�n����<lv��1
9�z��~Z���Sr�����.�9�[?l`�;���s�^��V����Sw��0O%���&W�& g&�g���۸
FNšD���v��l�>#�:,��u�M�ړ���R���lM�*�&;�'�Y3���c��~�6]n���)g*��r]�d���! ��#��Z��-Ƚ3{�d&���[��|D=��ID�*�Ҩ�>ֲ���nѨ�i�B��~���WIɫ��f�*i+.0�]������mZ�A����J��<�T�E����������*x2�0V�B���,   �  B  ;g    ��  ��  ��  ��  S�  � h���g<��q��l�W!#2���^�3*!�����2B�*;�B�d?{e��-�%���N�u������}�]`R���ΐ�)����I�U8N�j�4�x���(.=�a�}áN2]ʚc�?-/�6K���t��e|�u���Nzo����Q[�ҍ�@� ce�S{������v�W�+���`̮y�KCf��o�u��	Mv��˭c�,�=�3Y�o,VP)�
c��6�������6�>�;jc�8��/�%�g���)Ĩ�%B�l�y�GID���M&]�v�P�*�X�,���	�4�gw�k�EaLBR��y��h��&�G�(��{������6c����������y��d��?g�[0�e�!�Fc��8
�c1�9oSp,�l��XE���A��ϥ;�{����~ܠ��3����/����V=ˈ�T��Ս�0f���6��q�C�NL��~���-m�G��h`�$��=~��cDg�ew�̭Ɩ�ʕ�H�F�a,�4o*����%�ѬZ��E\0��Ga:o+�g���'�+	�_�sl����HԔ{jץ�HeJ�*��j�{dw�Q�e�Nu~�!�'N���		dxщ�nzD��ӄ6��4�Hd�+]*S�|�+eF���3n7Rj8`��2���dMØS�]U��]̱���&��`�J/�i����B���6����U0�~�TOC�O����&	}k�>�i��
�
�w]vs8%͔��!�$cׄ^��9�,[4��ʄ'�������E�����>S�S=E��:����4��+�2�>7�A~99םz�I �n�ΚR��/i�;�Y���M5�s�Q�Y�w���<�Gϐ���y�X�*y�����}����N��m�ݼ䈲��������K+S0��+��ԫ� ��cZJ�Z�s�{Ƹ:Ξ�o�o4W�b1l 90	c).<�'��e\u�5�B7k� ��41F��}7l9͡��^gGs�$�ƚ�fF%��J��E�Z?eS�"��6����ݬ��B!A�d�@�c��:k��c�\�BjT?�k�5������u��M��=��i^�,0��T�0ʓ��+��̧h-��dØ�q�`ml��`��F���:�^\06�v�@W�dQ��O�i"�0���ğ-��x�����ji�� c����=�gi�����*�06��s���ܖʩx���0O���'��X"$��S3����{�������t�W��aZ0�U)��ݷ��~i�`*[��Q�s3��ą*������&!�C��S�6x`����y�h��ܔ�Z-�}��1{iZ���&F���-���*A0�a����Ե�{�Nr8Q����9�צLy��9������d�|!�1,��S(p�{�؈�)7��c�Xsj�#Wz�Px��,��.��b̚�=F�m�����8w�����v��X��;3��E����2���W�s̶4��U�����ކ1!�4A�}�	���џ_Y��1�������(��O*�F�r�a��ի�H�E�#eF0���4#�TF�F��u�QM����(l�TV{e�	��[����lp�`L+�+�e#�zҧ���׊�.��X�ꎯ��2�(��z�f�#�Z�m��f�G���Y%pcX%���������V�_8�9�{7m�&}0g�9��~�aC@� �u��K8S��_���C�Z�?$	cX�5�iq�X�N��3f�z�cÏ��/�(�j1�E��Ld��XV;�q24֩i��9��}������2�{���4޾�g7a,չRl�-u����P���5�a�N�d]�6���/����Ct��3�
d�ޭ±�ΣP��x
c�..�)�"�)��5Qį����\pM�_��ݽ��Ќa����r�FdלS7ٮ�2�N;��v����	Lct������0Ɵ���U2�{K5��=��x��4��
�UE���.:Е����ؚx���z?zH`R�~�iLޮp�e9�H⧋L��������Oc����n�8y���w�4�����ۍ�x�Fk��{���jH�+-0�>�9�.����%��W�]uM��X�2ҿ�_�ܱ���~�T��|�/h�ʸ\�1a��x�&~j������jg�ki�ha�LE�s�ן�F�㛙��`�7�wdVX��Rw�h�3��7��b�ؼ��U�39�4�u-kP��������y�lp����li�S�����+��ȧ&=�u�^\�CI�A����E�Y����Q#���0�oOw3��Uo�r���1�%�s_k���Uk1��ح��X���ǆ�%�o/��$�������
�=�df'z	4+X�ד��Nأģc���:MFڡ�6���0&$�U�%��|6��JDZ����t���0=�,�pVG�nʶ�h��(���
�X���b���\ȻLc���!	cW����%��p�a�5*['��8DwZ$inA��z��*	i�. qH��QNvO��$��־+"^���L��݂e��uȊalK�v ��D�}�$ْvaO��KcN��^�L�Ё���DE����bKCsy��&��y���ǻ}C�F�ac�Fn~�KG���[�D�'s���K׶X�\7���e��q�Ԇ�Ė3ۉ�ƺ���<��5��>�C6��ex3��]R3�VD�o���4���H\��j�>ú�Mΰc8�c�.��+��*���WFE���X�vê����N�W7��r�f�	:��&QY���s[���S��:aL�C������3��s����mh��`���֍3Jn{�-�h�l*�ɟ`�)�[���h��y�y�4��p!��YL���є�ܭ(>����	c^8�j�Ք�_J=�Z�ʦ��W��{w!~J�+�j�2������'LA0����@�r%�iJ{(�k��5C��O�kS���]��3��Ӣ�K��<�?_ar	S\OU�'��s�<	6���kWk;1�Q`���-j1��y���Y�m���(:H�'���P-ۍ���Vւ�Y�R_Ja�Z��~A�M��`*��Z�1��kw��L�#��%y=5u�d�KV0�`f�g��܊��H65�2:�j�_Lr�~���16�l��CFA��J��������d�e�1����#��3����'F`L.����ǎ����z�E�a8�0f�J�u��������R_���FS�r
I���Į��Ќ�֍o'J�������u�?~�۸#�6���Q\�Y����h3/��cٟ�/�x.4]�c�]yv����4�	l���s=���ʛx�B��آs�µ�Cy�RB���G�N\�R�#,�}gc�w��<�P�S��r�hc��}݆1�� :�l>�oI�Z��5r��0���]"&};i��fA���\9�!F?����*�����$�(,�1�u�[���a��zϞ�'�i�.A��`�	1[/�ek9K�O�H��[#5%���������6j�"���s�C�'m��-�)P�u�?Ș������S�[SNq�L�����]a,����6T�GM|(�&���0V<;��nf��IF�ى�B�[É ����G�����u�u;�|�9	c׋H��%6�³w�5���-��^��$m�k�A#���7썍�m0F<ʯ��G�|$�lv_��Oe�e�c����}
R�c7p_�.��%�q�;뵛&��-�������݆�M[n��C��r�oZ3~�N(��0���&��-���(��2G�����
��i2��H�B�{Tf���"w`L��dѵ��)٥͹�鍒:�d0V�Nt�B���QC6[��'��.�Ͽ1}�Î-��`�*�a^�c��tE��)�%�'
ϩu��N��1W!������_d\�u;�>z�1���#�5�Nf����D��v�ik�h��'����s�c����1��ϲ'���G}�!�s	�'�խ�!��)��cșcoXRM�;�X;�-�C!|w�������&����0�8�X6�Z<�1�l�K'*c��J!�vW��q��lٲ�)�c�W��9�Bp/��`��Q��X���|���6��������������Я��$"���|0��|aL���!G�V�H#�	��c�ϭ��*��/��l7sG8ga,
��8�M!��Ҳk|e�kH_���=
�������A|NS�CΟ���,q	-��J�&�.�s�3O�a�`Я��Nq�$��^eAt����O��������1�����a�Ϟ=g��A*&��վ>s
�d�zN�`\!gt��]��V^�1;�y[����y�,a��06<���];��YWB:᧨xf�����CI�u�X{�u՛�,5�b�`仑|���,,�0�@���x����V�\������Dl�T����10k`O�us�,�y��{���0��8�6
�*R�8��l�f`׀} X���ꀍI�oP��I�XӼk	�d����|��5`��Ɓ1#V��0��jY��g{��E��Y�q��v����X-�]`7��� 	l	~Y��xoI��O�%d��+�k`��ҁIsv�5�7��S f
̄���o5c>�fI���K���*"�� ��
� `;���� ��w�����JL�a�h9��T���I`��Z��3��,�e`���t�{�m9\��!����s�A��*�d`����� Ck���|[4���u�[s_�&�^4�b��VlX
�Y`{�� ����5�e���;'bȪ��6�>�@7��l�:0?`[��m���*�Ϊ���dH"���}�P\���L�q���0K`���I �f�닖�-���`@��[A|Ͱ��`�����V��<0`����6��g$^��3�5�0tR��������^K �,X03`�?�N�� F�XXm��ZL��w֢�7��'��ā����e�V�nh����L�=�{+|0ލj;r������x7�?�{��2�}&�7�����ɬ�;����΃=`��\��2O��m�]�9�N�������kE^t��Bp���ɱ�77`�G�����#\'�D1������l��"��ud��(��oD8��~�=Y|�{��v8�6�(&��O`�l�Ўw�db�b��k>z���@�$t�Z;�7V`����km�b'0�\W&E�%s��jMNY:	ߣL��n��:��3�;�aܽn���N���������X�̡���`S�v�~�B�{�u��Ӂ}ڃ5�n�/0;d�HC:"�xg���[��^4E���l�h�����sG�~dJ����A��Mk^-�ך�^2�"X�]:��4��?�`[�z0{?��ۧE��7����L�0`��rů�~��A7l����U��OC�5"����]�6ÎY�t��� ����Ȼ+R�1�~M���G��~hL�V�%�;�M�p�*�z��,�J�Q�A�C������+H)w�[��?sG�V�1�dO��)���o3h�?��;�ˈ����mM�$�~�0m��T��f��w1�2_�C�&@$y!æ�2�O]��jwv:/0��ʤ?�͡5��lGa�*')�I.9ޤ������Et����/��~����_�nlHՊ("��J���D/2I��s��¿4���|4A�	B&uc��� a`~�0�Y���i�����yƧ]��b�j��g?���G�n�}̦�Q;�bu�����6����2���W�#�O}E�Է]�S�&�u�n�6�`n�.��޻69n��lBxg���#�[��10�#��=4s`��L�1u�B*�[�f�uC�Ak�A*����V���~wĤۭU�}(3ĝ�k�]�eIH���P����P�q�A�Nq���1��]G��2���G��c{������Z8"�ꦦQu�w�n��)����X'�����Y��C���2T���A�F ��G�DK�`n�昱������6�Z��ͯ.����7���}Q:;z[6�Mc͜���?Qp�P�ao+B�"�)��}K4�CF��]�������g���LV?3H��h�-U�Q� �
����xw���|����B[F�38���
[�����X׺�����/{r�|�,�Ȣ#������
qO�H�{E��Y��C�,�����{r_f���m�j[���R��aQ,�V���1���t�_dtFJ�ŽB�w��"�m]�InclI�6\Ǻ��_f���ܚ��O������ăw�~( �
�X
��������Rw�-'�VZ�4�\�X�e�3(	Xӡ�?2��n��������K�6�<o�*R�f$���4�S`w�S*]��y����%�~'��Y��g��W'��\�H/�(�8f;Gv���
��0�j��c+��8D#�%��؏,����;�سc݁3���5]e�w���%�J����QC=f�;�0K*�e-��w���b��B\�������6%2���~��1;wdu�E�3�-a�\�9�6#�H`��z���젓:�ִC��v���ݬ�]�Nv�r�*�E{7���"?�k�n+v�-���.Т��HR�{5yuZ��:���﷡$M����q���� n�h�m�g8���񄈈�̊����2Kʊ2����MFDf��ٕ�2�W�JhIvC��]��~�빟����=_�#B��K�r�,$�:O�j�x��vlL,��_��`'�:Y�.��>b�S�j]O}5��oI��}[�FM3�O�j8�*���z���lWcu!���-�
Ƈ���l��Y�OXi�ڧ�;��b�w���Sr�´ �G�Z�`�,l ���I��K�bC��{C�͙�B���``��OB�X�A��XWno��?��䮭�S-7ۆ��g	�C�Z�3�:�y)���~GGK�69Z�M�u��t�I�@�!�3�s�A	�[ 
g�����y�n���?]C��a�X�*�00|W���[�Gq��zͿe�f	2�>1��l�[�� f�MmL�,�	j��?�^X8�zi��h���J��f���F~~���.�\=Mi�ٽ�L��X=�ʐ���R���J^W�������7�8�V�7`2`e`�X7�8�t4bG��Ǵ=���a�.���1���:���X� ۼ�O�L��fx}�ӷ�?/`-�L�+��+���Yk_���kM}/�?=��,�c@ʺ��]����O�<�ش�8{��u����^�$�*�ER8���b��0/�I0i�7�����q��`�f]�^�~��>bvݝ�.Պ=�"�ۡ�	�
�gz;x���w�
T�N?�#�6��`��$a�c͢i�	�nF����U�43��Po������1`O�d�����r��������0�M+�x��������`�P��I��&2d�{q���������9~.f[��n���)��]QH�c����`�\'=n�j@'`Rl��w����z��+�-$�n5�,
�F�20�L�>�e0��>�1U�rz��jJ*��a�燚/f!`_�����a���2�m�r/���fĥ���?�+D���z����,#����f7��_f���ua�_0s���_��K���e��vO��?�-^JE~Pސ���X,�n��`v`H��������W�ݽ4��*ǩN��A�1�����,�#D�=��:�XX�w3!5_�'C,�4��j�d0W�S�}H0��wf��OA����9<.u���'���!m���Ĥ������R��z��.����-�4���;�4����5�,�LM�.̺M���ę���A�RU�~�כ�(�28;p�F�t��,S&��7���HɺM�D�(�q�!������w`�'�q������� ��ٚh墥~�fe����r��o�0� f/�QĬ��-��J�yŔgz�Iqq>$ǡ��`��Q�%2B7mJk�=�zFk�T��zi��h=ڽ��BR�~�;`�t-$`K��8;��1��%`�\�Uc�MeS��x�l7X�q��`��f�&=&�:/J��ڝ�wJM��q�:�I��`J`
�Z����
���<��H=\���{����ko����l�x�E��skr�
�nv>�%��A�?�?D�>tj��9��}���aF
�Vf&v�	����Z�ݗO�.JIy�{�W���kԊ���V�pb��d��m��yʬ]���^��R��h6�����Ữ�{O�nsB,,�XR8�v_ҍ���k_����G�p���8;��_#p��=���8E�;	u��Mq�x_#�\�v��L��&�	b����c\U�~�_#ĚA����d�I"K[AmL��|)�((*���q�|���L�0���=_�+Ҏ�d�.������3�>��O��ia5�������8�!00F�q0���H�6��Mcrc�j�p8��U%r�2�>u�<1�-ٛv�Ȑm�q�����"�$��p-3fv�"�l�=XSD���)���+���K ���,F���/��$^�^���(b�YfHwL	�=X=�(X�
3�mu��Ƽ}a�)�lM���9.����)�Q���9�������+�4�=�')_B�0��W�ứ����Sz\�&��Dt��ȼg��ғG5�>O�l�R��̓`��p6�����e��_�.<�љ2T�������r0k5@�<�Yr�u�A�\��"�YfѵVM!&�0�Fd��E������1�p�RN�-���0��W�k���#6���zz��}���r�^��O�mM���[�/�go��.���Z����Ƀ�[%��x�Z�;dnT��h�^��w��.#X�N��0�EǢU�3�/�w��W�/"ᙉ�Z�������uG| �1&��7w��5i��ߔ��>��4�Y��$�Ӧ��L�^��`�``��oȒ9�<����ۦ��B�#��fLz�=3���:Yrѷ�1���S�8NN{dsP2�&�K``y8#tŉ[m[�I��kέ)=qҽ[�8QPQ��Hˎi��`H'�n�igq�`��<[�Y�齺^�Q5:<�{�� v�i`V[o�c|�'�Y���E,�doM��#F�Vd%{k�Ȯۡv	L������%�~��uK�K��I�`?�*K4�9��lmֆvԳ���ۙ�F���S�|\7|��'1��#*R�}���/�i�|�C`\`�Xw��w�F���Y��*�;��%�(�EM��<�\����;�ֈ��M�������֔Ķ���<vlg�n�ޱ�S��[���]K�#"����Gv�����ע�H�k�4	�=��X9X�֓&)]���?D��F�$���<X!�f��Q��,L۝�����@$w��N3��C�t���j�`=D����/-i���}�N��ii��5��у���y��ָN;�Lk��N���N�6KB�� u���K�>`�`�``��>�GW�m��Y��l�g�Dz9]a�hغ7j#`�`�B���������,ϯ�Y]�/��"����``��\�[��%l����	��N(`o�A����%<�Bk�E�e�`f	�6VVv��P�K�SCQq�5�9Kk���ȍ0��A�����Clb�S��y��1�+�~�6l��r��B��	�2��Z�;�'vt�)ٚ�[��N��m1�;��*�`�'XD�I������L3/����������&B�H,�>����� C����x��V���q�����	Yy���k�k�<?�@d��Q�K�̵qO[�Nܙ�ܱI�c[_�e��O�9L��1�����ő�:O�
��\�dg?k�y�+�+˹%1��`m`�`������:33^��M��2�v���S���vl�L�5����{�Sgu*%Z�7��t�]�3v!p̷g�`R`H��+m�@�N1�^�,h}/4���mc��3z��㨛����.o�7��1�[ �}�c��Mդu�N��ȴ���쿁ف}�j����"�b]u�;S�\k���>Q��l��lB��y�����.��ݞbe.&������N��-�|q-\�N3s���q;�~�`H'I���������z���]���:˩��,`�``�`�`�n3�2�}N����.�7����Ҡ���#�15�4�[��jћ&^K}���������r?�Ŭ���	c�'��SS�T���ng�,f��ަ}���_�y�e��F�3ǌ�lL,���R���_,s�d
}h�>��������`�`�`�D]�?�%m�Lup[y��0�>:(�ngJ��Id�N��s���ib��މ��{����-�.K%�+߮}A��޷�k_��*�kq���s�D0�C$��E����.��;����=��l�vԨ�|���Ļ�yޣW��§��.#�xUES��.�����3��[�[w�I�$ɕF�X>�Z"�$�k��
[;�o9����)��N_�^��Փm����Lve5�3�; 6��������������w�bC{v� �Պ�*X�-qK��D�l)�GT?��yK?���%��z��1k��~�-��%�l��k��]3t��K_{��n��<����ozr�>8���L�ll�,��d�<K=��,_��)�W�߂0sB�����C�N�8���M�op�Μc�t8ۂ��j�`a`wq����ל/s�_<)�L�i�9�G1��Up��`�9�'#�Ʃo��%f�{�'�sO4�mI�k�����I0m�E�&0%0���l��b��M%W�"(�,䌵�}��aV��:�Q���
"Q� S�����M�!�%܅�\έdջ�
�3W<C4F^��KIj��՟�N�["�d�6�/�� ��S��ԁ�q�H��`����n��u/K�H/��=w<�@Xձ��\��f0#00_j�^b�/�@X Ϊd���)3;L�߳NfQP+ÙX��k��x0;�B�����O�m)�.6I$�UZ�<�=�΁=��3̐���X�Ƽ��U��.��S������l�(j�`�``=X��������k�����I���j�`�`�8#t4����jn6��q�,�4��i$9�X"n����&ҽ`۴.��&�Nj�G�Xۻ��^�r�f.��#�2��{�Y�x"o�@f�c�҄�6���~Z*6`��u̾<~Z*Jd|٨فɐnS�퉚��#�JF���o=�ٯoN�d4l�������2K����[�U�QݳrրI�9�ށт-����=�ƺ'��7�c/֏9���s/���3���7`�`e`�D�Ǌ�Nd��A����ݵC���0[�+~�Kd�`�`�8�w�q|􆗞#��J�q+o����Ü�5�,_�B����b-�u��q��YX2��Z�=�:c��V���lEm4`b`�`j`٘�B�4X	ؼ�~�ѧ�o�kG�u��_�/�%��.�~�����,�wd˳� ��f��g�u��	v�lh�����N����Z�-� L���C�	g۳Mq>.�gY��D���������Gw,)Xf�"����%�B��4��Mā��&��%_�aI"C��g�}R�^:��L�7��2��+���;
F5y���/�I�ֲ]��n�<�@�wꛠ'�R<4���L\p�����]k �kQ/�:�1��H:ֱY��G�2f]��}[;������dy'A������F���nz�L�f��q����p,��ˬo�{��{�R�*ID��qv���2�S!I/���4�avA|J�Q�Yv��@�7ݼg�O� k�#+C�̎G���R��jk��ѽ[Ǵ��p�Z�E�[�5�"�M���,l�������+�I�?<�M��6M�uf�[|�R��tWd����q�N�;�g��fbo���1��b�`%`g�������V���aE�:���sK9���e)�/����q 5�;f�s}g���t�
�~�*���2�j*���~;β�Z���e��˚�k/	�ԫK7��{���������E�����&��o�!]
?�����r��i�zx���m��nZw�:���xP{���֝�Mq�$��U���^U;�⚌��!V
�K5�9"C��`�N�]W�c�]�7^�!�%N�z��zt�u߁��6���A��mVc3������R����;�GV�vЯ���w`d`�`����-f���ǝ�����F�E.d9��(R 
����,�P"KZ@-l�}t��l��Y�7A����:`~`�q���o���׵W6Gl����|�h�4�/x��p=ݺ�� ���f̞�Y��������)a��۬j��߲�P��b��FͿM�100w01\�V�D͏l�gz]��Ӷnc���t>�3&փ3|�i��b��ч�I�����|0�����Y�S
	[�~V�7�+�^�YfK`V`���{|y:)z�g���p���eCU�0>01�Ø��&
v����h3_ܵ�B��oo����/�!2�J���^�������ȩ��|2�~J��w�}x����P�������}�=��:��_��9���ז�ǲN�.�u�s�S%���R>���TkӤ5v>_���<
l6�	�
���7�s8�C����Ɋ�듋�^���#���] b�`�����4b9�7*�{s�U��{�U����YGcc{D8��\{��z���3�� k+ k��!��vq��������������Bm,����'sgͼ��O�}%�]��F*!�Y5�)�g8�wf#맼F�ϓOȦ�1��Lh���,0�Ə�]B���M���fb1_��z<�Sy)�{ẙ��Ir��`�`�����N�K&�{��+�'+����=��G���GE`#��L׈�9��``�6Z��� 9�E���o�	�ɝQ�o�&g{G0�(ֆ ���.���6��<����p:�(}��,b�`v`��t���΃�%�4T����u�����4�M}�$��,j�	�t����^佧��ȣ�x���U�����@�����!�{m��{*R�ED>}��?d_�j���OAb�i���!U+}��6�p������Հ����x�Cf�{-#���Y�P���`�`o1;���`#`~`�XwiOH�)���I�?׿�1�nr^&X�e�H�R���Ś'�}��恹���ʷ�Y��ƙ��wx( 8�O�ұ�x�}�WzI�wgn��n�3�=ߎ���q�]+� ��w���z�ߥ�k�k=Z��q�}���_Lk��@�/?�&��D��(��{������޲��(؞+篕"X�cuQ������뤀���*fɚ>�zsǎʰ���m������1��Ss; �u݊B
��	&��E�h�2b���sB-�,��=3M�6�l)�$�r�Ħ�h�1fN_�7�l�"2|g�3�7W�9-b<J�"B�|N;J:#�o��1�[U�ކ� �u���f=`�`�6�n����f(r��ޞ�	�
�
V&���7j�`"`F`����~,��}��������&Q^8��a��(�S�#ؾ��Ън��k�z��Z
�����d6��9{XK����tx7��ߪV��t��,K��g�O��bc ks������1/7٭���j֞֊���I��B�Z5fe�c^���>�)��Y����S5���������́�\5}��m�@��CV'2�L��&�R��B�b��f����mOxY��̐.�	,�1�"�����ȟMy�1?&qCKy'�y̶����L�!��W;_��"��>�E�^�����oP�+�����tDn�ؿ�)y��\�?�yU��F��!�_Ù�gmR����j��^-�Kɞ|�g��ަ��%I=5���u�̓!�G��	��
v��uZ�Qgx����Qo��T�w��;�:�����`9`�`���>O,��k���?f�:��Ь�P���}�0����ؒ��-�yr�8iEŎ�플Z�-�I�����Kԭ*���3���呤�_���x{Dc�,��	5��6�O�΀3���s��R8�l�d����%#��~�s`�`��\������C��F�b�U]���	�Շ���>t��Z�'f?�����.��,Ǌ�Pe�RS�	�J[�N�;�Y$j�`��(��c��c�?�J8�wҙܵ�,��� -�f��������T���>Hmi���{����.��$)η�Bۖl�`H��7F;��3yA�#9N��/u����o���DkF	V
�v�%b���q��"3��k'���ڜ���
��"������ADF��-�+�0�9��`���bs&�'�#���m��9i:g�J0�s֫AR_�O���u�^�
Yi��'�N�6�3��c�,	l��>�
��X���T�>%�a�9�'�,�B�|���¨1�Հe�u�:�l����mE��@eoͫ��?y���>�~�*��i�ỿF��d��3#f�V�j=+���Zw���FO8bW�2������w�3�cK
ޒ��(6�ok"aRg��]� �����8�����Zhl�\ߑ\S�5�k<�x�&��mQA�� X3���h�߳�p��I��C�A2�]��2/��F|5�`����̓	���Y$9����9p�V�@�k����``�`�`a`��i�Q�ے����T��<�AaO��$��4jS��Iے������ ��g���g/���Q�c��v�?C�@��?�_-��n\�*>��$|=.3��Zĵ�(�lM���c�t�`S`�`z`.`\��C��΅ �2�T{�X������]3�%��;O�lY&��=�8�E��>=;5E�� ��(O��4z�!���r���hߒ��}y�FOnO�7$�����l�*��0�'y��ݏ6��v�'lk�N�`��$�>�I�!�f}*�倹ڤ�They5�q.M��D���m���V��D��Z=X���{ߡ����8�/�d��"d�_^���!X�����͎�Eöwٺc��s�����߯�}�")b��ށ�;��f�.�"J׵#U3#�g��ȯ�����`0/�<�ɨ�bf��3)�3a���h����;v�;�(,����8;��X3��&����.,���YAٍ�)���7�S<�T�޴8;��� {f&ڪ�S�8��z[��<����������0sC����,����f��;�g	��T�-j��6Z�)XX��ڪKi��
�Ɵ3�V6�v�X��Z�P����b�Oc�mv�N��g<N�;t�Ӣmu�t�+��zZ8�
�v����c�K�sG��[2�5��Oצ�g��i�Ls��e،s�mD�;�Wn�7���]Nl=ܔ���1��9�����l��M�|�`��Gn0ov����N���x"why �n�I����l1KcS���:��b��a������I��]����`�&�뾂�h���l��r�e�e��?�V#�"�C�Ê�C�`�8�wL���>�!���X�qw�K;��h�2�폿z#v�8����ܦ��3�>0{jsu� }��~�Q� y���`:`�``�03wC��,l(�#]]@��"Q_����jDfz��"3Hz�vU�v@1����=��.�T�v$�{C����h��);�bd�<�0�@��[w��ԧ�k#��%�5���+���5�M�K���_N��ҹ�ͽ��| l�Y��9Xn�K�."C�F�i�W]~ߨ�{_u��goI��\���2?���ig&�}U�������%uFqR_w�8��~^|����A��`6  f	v
������xq��.���/�a�|l�1s�B���_0U����V����Ƿ����ˏ�"aCm��g�.���=��i�5��7KX~7xVUY�ה�_��f��Ui%�6-g��ڻ�R�||��`Q@����1�N`-`M`�`T`H��� �x��8��p�;)SkwB���#���x��Bj�`��ݑ��鐓��}Rhf(9��P=��ق�r>�Z�u���NFZ׹��Jh�i�_�M�Mʼu�'�݉�؅�X	���A��`_��#I
�>t�Սs�Դ�����0��y���5G�����
R���c'�}�쫉G�bO����7$�#�}�|��V�$l6��=)�a����Qϕ�#�G�׹wo�#-�/f�`���������s����~U���M����`�81[rE��l��2����
'�Q���kI{�g�-�yP��;�3B'w1�O���8-'��y�.�=�bMًm~�l��9LC�vvK�\&��ѐW��t��q>����7��� ��3�0|��Y�������
��\���*:�\�*���VN9���"j�`j�4M�����ה��EQ�tl�Ō3�ձ��c��k�˿dk݉��������e�s���ئ[Z�[[Č�L����ֱ^��Y��UDhf�E��*�粯 'j�`{�
��qb��.�"[����"���=�����(�b� V�g�����!V{��˾Nh���g<���qd&��&doe$�de��d�*QY!�"I-3!{�*2"�]�W"#��st|����������z�y��>p��Ю��`ǻ���$��y`R�v�z���1�
1T����!�ٹ��|���|���jN�1������3�.�����QUhz�ZW�,�H�t��ʯ�&����6q������L���r����:n���[������1���dj�0��30
�5��wp���u�cx�'%\ϊ�{��L�
ll�?tc`Q6�_8���$�����>�;�!5�������0�0Ԗ(W��UR��M��#��Os�U�)���k�<Ǫ4�;�e<��V�M9��H�Ŧ��J	H7���2�OU0)İ[����`O�ހł��h6���?��6�P^i��3T[���ھ�]Sc��P�D�-�X<>9}�����ڪz��������1��=.S��ք���a� ������W�,Vk��[6�<���� �T>�ay�y��w�֜��<����U����1�%�X��F��ڮ�)/�oQ�g��Bq��ُ��Q�u�����VA[�0Y�ق���_�pV
�E�i/s�جZ��&?���w��o��Z-T�n�n��f�P�E��?���=�F1ʮ��]��K 3���8\��t�~K�|}eX��^i�a?��`%`�Ih���%���S[n?�ke>*�41Cw�ʑl �΂a!�;�y?*;u�D�^�߽<�&�yb/m��^K�H��I	n�`
{51�!bZ`�`g���:*�5�;-�@3,��~czL�0J�"��������'�kiS��r�������7P�
Fsmx`�;ձ�IH��$��qv
}�`#i�~���W�n�ps%p���G�:E��`��o1�*W>J���#ۻ���l|3��\��+��V�����k����;�Er�}9�O�zΡ,1���'7vX[�Z��-y����(b��O���/�#:��AiG��e<�:7^BG{�1E�o��4��,NMR�V	�.�*��$bT`m``F``�`�H�yX6�O�M��Wjw=N4S�B[�8�j�x��0:�Sf(���4m�FBt�����T��<x"b L��0;&eN�؃'DQv]�^���P�%�W�r���e��E���2�)�sL���JCu]`7EDB霩3��c%,qI�Ro'�Y���9��"�ǃ6{0�0-�}�rO<��/y�2n,N^���ab��vLL ��:}�bf�:/��H�at�shf9b��OG>;�1�!:��=�D�����Nb��?if�Z����xyQ�f�C����p�|&Ǿ����y��\��Q֏�����G��;���Ι�+����0� �2پ���y*����>|XLz�6��|;�lg��Z�#9���/��ߒN�]�{X2~q��2N�+����p���/םF]�S�$�?a+\������G���J��F��3��|�\�v�����缝�rO�?�M�M.�
zz�[/b��Yf�&h"5�9���mI���k���s����l�`tt��B[+bq`&�h{rT��9gR�x����	�K�&���)�a�`X`x`}��eӡ{�'��S�;��f,c#���	�Ö����p	$�)R����ΈD5xKM��F&F�XX&�/��;Չ�<���ngṁ��lQ�t�Gd4���
��B��7�)�:>�4���(�q�+a'�)ڜ���u��nwo���>0���S���f]7(>�7<-T İA��`��gF��P����Zd�ؗ���F���j"6Ɔ�"X�2�;���y��@�5:���k��
Q���i۶
vL�՘d����	�Z����vI�*;w�޼fP>J��b�`��5��~����1G�j�lw�꺨��|]Qig��7m��1`��.�p���0���G762�-۬	k���v�ػ��G7���6j�B�.�̓���o����L)�V�=��#N��҅IY���JUI�S�)��aM;:���D�M�v2VR��Rzl�j=PN��,��m͈Q���6�Zo)o5�p���'�](���*l��`�%�=�`>
1#z|B4���b'��
����bFt�.��N���9�k��g@��Z�L�>�!���U!O�/�.��6āY �	�v��Ow���ӏwY���惜,'&q����wFb��1��"�\	�tĵ����o��(��?+��r�N�Y�łubt�gP�s��T�(��p��=�C���RI)槈q�Ub�'�Zb�|�o#0=�ZT���S��t���_ݒKh�3� [�����������.E3f�3ă�ANb`70�L�ou���_����L��~Bc�ؒ�A�>��S���i#v�k�郕�Q�1�<<GyK�EX+ڷ� �r��[�����)�%�)����]YӠߡ�W:�[�l��6/�5 �
��P���%t�F&��ew�9Urۿ��s�XX��%9|��b`�`u��] F��hO)�A���Wg�<�>���m8��)e��9+(6�f��j��]�������q�6��IM�.�8�z��u�ǰ�e�`�K�<����pk4������d�(9�	� ����muo�^��o��H��zՆ?Zi(��-��a��2��2z0��f�s��<ߝX��N���wXG⑘��� �@������J�i��z�f�������S��$�ӵ��ik`O�����8���D�9ԙ���3�Z��J@�"X0�#�mRƷÆ��7l:Rj�޹�~�oY��ٍa�J��KF��wW�ݣ��+�;B��݁���ZWJ���t���0=0sĂEOTi(V�="�����伕���#��v�bE��#� X[��ښ:��=\Nr��Ҳ�T~]�=p�)��@����ݶ�55�Hj*�Ӟ��}��zfٓ{iM�`��m ֌t�``�P[����gL:e?�o^>u��z`�5��!f�7��N����u/�'���ǜ��X��������Ə�W��`l``��݋�s�#=!�t��;���1�ܮU��<0	�h~���i�]��Z�s�ޟdE#��6cf���q��Z�{�;6	ffqn�P7n��oy�{Ymy���!Em!��š�>`1``�`u��#]1�)���-�1��S��ۈh�7��;A�_�,� �.b[��kb����k�T}ΦE�j}ͣ]dh��ow)`�`o�����$*�hD��X�>�j}�p���3 k\ٶ��ð%*,hH,�6}�/��Eih�$�63�V�h�F���Z�t���ߩ����Uy;(�yk��|~���N�Y��ݝ�ݙ0���:F���_b:N�_k�4g��&�XX��X)�1.�09��WKбp�\���6�Y��ﯾv,����0�}'Q]�����<e/��ri.�a���n�A���E���q"���������]��r�D3��2�kQlܐd��� �b?�����ѷաl	���-K��#>Ί��G	*`3ꃕ��@L,�݅�E�i�]*!�|�/o2*�y���A]�e{y��c {�)熲r�(����:�q����7�KO��)�9�� FICޣVF	�v:e0C�[�EO	���m���^��@�0���`z���t.�M��x22X�tW�iV�(	\D��22����1�łq@G�F��5�*�@�����^������=����x[�,�e��"��1�������:�+�&[X�����.�fv,�m
���6��/c�Gm�^��]�M[.Ᏹv��f�����v(��4����w��O>>h}�yG"z}o��$�\ާ`Y`�o�-��v��Q[�K�wb��췴��]Vl�:x\ mu?��L��u0w�S�e�)��hg}{�2�u�D]vcI=�$�{v�D0q�*�rj2��}E%_OZ�8���s��DY%bB`�`�`�����|�8~��\{�y�T��d1C������ �	vL�������P���%!iO�*,E��a�ԙ��Fv�	���vǵ���s���n���t1K�\�f�o��~���#�6&�ͭ��o�W+-���0U���gn�W� �f��2�N	�s ���(������]������^y�ah�6v�(����N,�w7}�����L*�i�ٯ쿈joN�e@�
lu���1%�.�/�1l����-�y�M��2����6_V��q�e2?�].��_����L�CC�:��&�#IFJ�c�ŵ���z��s�R�F�l�f�і���W�f����|G6�4%�R��8ٴ[�����]ؒX�R�1��6ڜ2�r�b�R5�1J�`�`r`�`�ih�A���}���\5���s���zV��G�Ο,����|����N l�,�S����Ǟ�u�oD=��������G�!���c�Am3S.�zkn�R2�j<J�y�Y��m�/�p�L��#X4b�z�E۞T�%��W�I���{���XT�m����� f�&=FR-ta^��N���ڙ�9��g'�n��m00&0&�P]�����<r�Zk\r���u�Jg���h�~���M!��FVC��e�G���ԈN=�c�w�+�\՚� �X X �k�P��1�k\Cm��ϗ���IM���Ct?�W�a�8b�`/����'�mY�o��l�����!�T.u�r'�룉��`�`҈���6�;Q0_0^��ֽd]#���=�Ğe��u�g�@��[�=`���(�ư��;l�R���\�.���]�YrNaö(A��kv�9�����3h+1"��8H��n��Dh�(��ʚq�.�80���'�����:��H� 9%aG�&�y���xib��O`Ѫ�`�`2`E`��f�Xwd��l��xq6N��D�5�DY����-�ClfG	�S?��2K��;G�*����RW�&��̯`�b����C[/b�`��-���7����X��=c'�B�uNmX b��(��~�}���%0��ď0�$J�y���gt�� ��0i0l�y#v� b>��m��L������מ7��M��+ɡ�k��
����i����R�i����]��5����'O��1[:��C���F00:��&����uj�%4����Wxx��L�	l�4b��a��b��"���}*��ٞGċ�Xb<`_����������{��_�������ό�%U�[y����]SE�]�����|��Ӯ�_<�t�Z�!��ׂT����W��#���8;����?�;���������Y�����/��NZ�ŀ� �ȋ�l�������fgr�_0Q��_�x̀kq$�G.��.�q��L墌����]�w8�?��m�������f>K^�AL,�ぽ�`�`D`:`^h�	��qbk:# �|'������8�`�`5�bQ� v1쿺�ŝ���G^W+����z^ָG�y�4�Ru��X&��p���h{�،�c̨���ͱA�l��`�O�1$���(�FldG'��>�T�ۅ���o/%����ީ96��X��I�&�|[����^�b���[?l�ɣ�BԳ� ��X�D�ʶ�|�00�X�9�yv���S�i�Ӿ�=G:w�o|۬���Q`�uG�|c��M����@�{rc�Jh{���k��e�A�60�?����iGSua�}�s�O��|*�I�[X�����W��<t��H2�%<�@/�C.%^�8���vL,�3c@u\�/�r#�O���YIu�&j\�6M�7�LL��#�e$m�$,��.D���y��P��O	m�`�`�`�J�]M�vw�UlI�lL��#K��\���է^����İ�����#(��c�K����4d���`Y�:P��R]:&	�1f�V���LL�S��qV�eKq�y�Xx�7���Y�����L��ư�ߝ�)���2Ն�F�޲�"y,p���`*�\��;i0?�W�����띗�b��B�W��2�O�4x{����n{�a�u$%����'���C�G��9�AKR�Ɓߠ�6��6��m�`JZe�z�q��r�Iڴ�GF]S�*�G�'��1LwG�fߪy��cUȇ�K������@ˡy� X;�M�%�/������IX�ʩ~3?ڭ��r߱��
���=N��Q%����f����O�_%�-)�b�m��r��D/�i���`�`��&V��a���������=����=-�1?�~mEZQ�1"�~0Y��?݇�6+Oi]cʶ/�_�b$�����o�ǰM�c`��C�F�bY���ԇKI�H?���ˏKE��,,�k�Eu��	�?Ш�/���(�\\۶;`1�,�Ӧ�0=�a�x��7��6b#�LB����̠�,�Lzf���ݣ9k�_v)�٦g��+ފ���^Agl��1��l�zĲ&��+1廮�2��΍^�%����ݣ�%����������D����_��XZ�l��&�Y���n*�����m�=|����Bwϧ�h�Ȗ��\{��Ѭ�[�C��i}�Z�������])X�R˖�+T,׌��~��]A��qjG�;�t;��ö;�� ���S���ֿ��.���d{�DGG�glj�ܞP�Ǡ�L����!���r�$�fh�D ��}a���-��מ����yr:�7ʄ�ǧ>ˢ"]>���4S���o���FeWc�C�T�q>@|�-|��M|^��U��1�%���J�Y��R̋ˊl�拝u7����I��@�Vp���p<��9%�s˛�f"ſ�f����@�?(//s�i�e%��Q�S`��~��|�{k�ٴ������<������B���9gcH�{b���������yjOVR��cJ��0*;���~��	�$X�
b�`c`S��[���ʵ��5�yMW�3�B<%j��������UY�1�Ҭ�qƏ#B��߲�o67-����?X�қ|���M]��;	�^'o�$	?��6&��;`�;,�)���{9�G5�j�x�j�vc���J���oɮ]g�\�;֊i�=h��� �5�ڨ��~���Ѭ�faQ8��2����CƉX��S��w�T�٠�v�e��Y�g*�#Wz5�2�|��1g��Y�dIT��#]�*�U���I�q�]��=�;��-�v�o\���������,��_&)]s��ύL<�:���{�:��,�\� م��f׷���C��W�H�=x� Y�.�����eŇ��b(�=Qv���b�c�&��� ��w�z]q�]�fӾ���S��xY��`\�����<c�Y咣�(�N#����ɠw����Y'&MÕ��=e�]�@���~�����y�P�_Uw����a�/�-��e�?F����L�?t�`��f�ڇS���:g���[ ݍͱg�:�:|1~���qeAs��l����$���H�E���I9��y���<F3X�l�IT�F�������Hl�"٥����B#s���O_�Qȁ�鑵O�8B���I���N���+8U|^qh�tu�c�L%��B���?����W�a�U����8���}UY��I˟���U����:��`�%�d}J�Ă�^�����W?���4�j�t����^ֽ��ӘǺe�?��mu��~�8�2Q;'`���,3)�޽��WU&:���Y��!V�l�cb�iM��!��:-DɡR$}��קWS����z_���R���X.�U�UA��^z�k�t�)���S�,��{�ƞd�����d->���fqqh����a�Q��L`k`]������}-�
o��)XYwcd�8��ʐ�t�W8U����l��F���Ւ�����`J`��7DUhj�J];����v�}��1�:�}`��/��ɒE���꽞�dC��g�9;��n�:谌��%�qI�����e$�d�� �Z�Q�G,"��#k��M�^��5"aa0�g�L��`!G�U�&=��6<u��mk b#`Q�����+�o�g����rY��Jc���g;}���f)����gF@�q*�@oeĲ�R�<b_�=qUF,�Y��at�`n����t�d^
?]��V���&V�ר���SU�ԖU ]!ҽ�)�^�/�װ�Y���}]�n~�c�M�XĲgs/����\�Z��@c���NYF���Y~���BJ��O3�2El�I�X,����X�.��Bh²+Q?]'��Y�'^�jLs#�/��?��.��L�k��>J���f::b��j0쟼���iA�}�z�mF#����-z`�`4`ռ��B���(X;b�D��Y�ot�Wĕ>a��חǴ�����n-ܤЫֳ��r����ڞ�|ٛ�8��b֯40k�w�ߌH��۰RQV/L�l
���/��M9M�i?	�������c��wc������x
�M�����ҳ��o޲�T��vv/X�R�:�"�V�뇅���U�1�<"�3�C3!DBJ��Kf�1��)N�3xZ���r%sRVvcv#�?:}�U�f�o�H2=%����&r��5(�ޯU�'�|M3�n��饡/�*OK��zx��޻����a'
�����Y��	վl��j�؍���3�j���}O�+꫓D"�����sY��7%�+�S6!e��܍�![_2�����/��kCx=e`7�N�����M5�sO�<Q�M�n,�HP�^����}��	vcqW*�d'd0�W=}1w�8S-�n��aA܏j�?7&?��t���Y4V��I�{�#+�����J~��n��B�bR��
�Q���8sn����11O��{2x(7]��*���8��2���+�K�5Y,�؍�\~�9l��$-%����.�q7�=�"�"[��~�)^������wcÍ��.��?p1���7=��_Qk7��ݯb���8s�ŏ�2��wcd�C{�+_�������|E����n��ZVRΆ;������|b=}#���iz²\�i��L��@���C���;��m��6���^*f;Bu)�Iz7�(��x�8݊+q��jX�<�n�X����Z��O�.�.����5���X�{<S9u��<�i.I����o��&�HNuIJ�$ͺ5v����q7�Ae_��f{��a�iӦi��X��1� z�b_��j�[R칵�c�� Üᕔc����ͽ��vc�:m�̛s����	���b�;��j����6&̦'����7܍񟨸�Z��B���cQ���⻱u���X��:��W����Lν��2�bX���gS���~���Xy��¬����lZQ����ؽ��<ϵ�-q�+7�]��ݍ�?�
��h���e[�a$�%���[A��yh���CBR�;�iiA�Si�P���3�����_��Z?`yۯ�?׆"K�#$���H�!�`>K5���vb�E,�1L�@,^d���"}lƾ�ho�y b=L8>;��k�I���UǂXt�<?������;;�{�1g�r"廨���A�QR]�3X����r/��)x��IXu,-E]+~�C�fS5$��̵x��'�rĴ�=Պ'�O�{飛"���NY�a�_h�R�~��D�Ǖ=�޳{�����b�N���_䖪(�(�z���K&=�
N���~��a�4ƶ���[L-�d�t�! �����`��<i��W��?����m��e�������?{ՒXq��2c��$,+�֨	�7ҧ5��T�S�y뚹�ˈ�Ϥ�β �lP��o��FR�|ߒ�d^1埦����g�b�s�pv��ȳ69]s��H"CS?Z�{ۅ��7��7���'bF0��M_J��>Щ:>8�!�iO	b�,��÷�%��y׽��/@l�F�p#[�E���%}k=�y֖hj��d~�v��"�Ć�+��	���ί˘�g���ء&z�!Jע�~56�V��Ѹ�+����/v6
�SͦY��{vƅ�eZ���T�'A��t�K��A�0`��vR|1��f��y����*��Q�[�б��w���%��Z�XtS�tjV�Ġ�Q��(*��*��17��=�a��������X�5��/�<�����L	=�Ht�@�Zl���n�o����p�p]@,S���|��|�Cz"c��'�����Pi���١��Fu�Ӻ1��g�D��]l������jSTۜ�Q�����8U�S&���
�������1u��5M=�b���O�L[���l��n���V�W<Fm�j?0x��`��p�)��L�I����m/k�:���}�<��iԛP�aBeY��h�C�@�FO��و�Rv�ü�����QI���2���VZ��thT�_��#�a�+����2?e(C���Q �>�^f�lM���7vB$��!����WK�B���؆₋�'fӪ��D�(3���q�y�ݬӫ���ڜ"�C�϶�Y��2�\���6%���2��&���]�ާ"T�c��¦���W����Ԑ�;�7_S~��|�>(�h=�{H$��{n��VS�}�.��Ƽ����F�"S�z>R�%S��	�ѧ3�a��0���aLgt�ߊ� ���}��!z�o�O���A$��u�LxD2	�LQ�v^Ϩ�}�#J���7�N����W��n�IF?#=���'�ۢ�zPI��+m,JR�����v�`������:g�߷w��p�;���5ߞw���;E����pHg=qZ��+�܇HK&F�%��d7���J��<)V�ݙ�#U��g��	�m����(������q���!�2�f�'5�T��h��A��5�����J{B�N}���@���e�0O���x7&�����li9��mL��*��?:��O�r4t�DȾn�`vwS�uU��ƫ�B��.��2�;�*����L[����+�؍%�!����YV��v �J=�Fz��� �8|uV����2���.^��@uXڴ�� �ܢ�]9�|��}E7w�al"���w�-�Ґwv��j�Q��`l�|69oD��ʮ��0���,s�,i4Q�ec��=c�N�(��Ok?Q��_;'��[Ȁ�&���Q���!ɐ�C8:O�6{t�e����`nX�&�Oxv8ķ�ߢSa=�>K8\�̓�`S��貮0��Ox]��u�٥W���d����!M�o��_C��"�%�o�A���ӣ?��Z*�'3���5�uYQ��������S���&|̍�h$��2����A짶���+�]m5P3уͼ1iG���<v��2Yf��� B&s�m��^�6n�v���R�͙���c]�:�E�/���_�^C�5/)�2:�ĻF����x�χvі�������+��(��ٶOIX�ŗ̷���} �B���q���I�1W�L�,n��u�?쏎ۙb�ׅ|��6���S���0�q�i��R�U�L������Kn��"��%j����a�����3e�M�ޣ��	��=��%@�:ۘ��H_X�64Y__���6�*_ylA�|3,��hi���D�r�&;]�؆�uOchl�dP2�1�ۈ�%����s%\�Y���g7�������}���K�C�U��f�n�'c���2��z,�)q�$�T]��zBi��3y}��oF��u�[%���.If6�}�CW�4��N�gZ�i�#��wB=l�v���t_�Ј�N���hg&6_neFᝁ�C�Ĺ*���o8Oo�<�Bz���]�+45wڴ2��_���?:l��l��^�˸�o��8��5�,�!�)&��I͟�?�T����q��j&2�:.5$�5���N[H�w(�0�s�.F2|l�3�u��վ&6���VȽ�� �76r�8XZp�Ӭ� 6\�kE����C�+��P�P/K���pd�3�Z1å!��Љ.�<�:�:$�0T��*��1/���Xg[��p�J���_�gS��Џws?��o��.KԒçb�g�u{�q�`�5A�j	��H�`��:�qs�P�>�-�xL�Y�M#K�a�Z}hF[���M���kG^�O��"��7ZJA*�û/��B~g�s�a���N�ݑ���'-!�SwM�#G�#�lX�ث0~o����FBA#l��H�W�T��Ѧ��v,������"�b҅Ժq�������"t��卟r��4H�2���C�_���s�����b(��K�o�Ϩ�`ߺ$��Z���~�<ү�yᾓ�OS�}�H[��e4U�f�o}3N��:m2.n�ǟ]aj�xVr�X5��^ V(��`�!������Hg���X�۩�������/�h�?K���^�Rz�*�ɉƘ���u�����ru[�ݵ�9��y�̋M�;)��*�g�����|lh��;�kLt��"�O�u�|�#��(K�+�SϠ���\'o�AwM�8 t��i�f�o�$G�E
�{ϓ�&D�4g�͕���L���B�eQЇ�'�#��Dw�2�j���,���0]�x�\�ĉ��2
T� 񊧥�<���؛���,PM����갹dL5�kͳ��fn���R$vv9;�1�V�/�W��
� ���vKy��א�d�}D/'j��ȭ�(�OUYv=7�����?�$Ǩ��������;_��p,��*��j�5�ԁL��_�������`D��ܷryQ>��"���r6/�d.��a(���}N���*Yp�}�\HZ'���E�PBNu-:E��h���˜u�-G�/�n�_[9Ȏ������b<�/X�,p&���u0���Fi�L�P�px0X~{>.�{���V�-�:�ps���bd�e�o6��34sv(U�����ܶ]R�j75���vZS�V�-�D��X�z�����zK~b�|wf�£��x�'���:K��Mzi_�z,A�������4��g��bf���6K3(����x V�K78�1�A��Nw�F�Sv�C��[An��?P����'jIH��0�"ė�j7N���|���0۴1�	}M
��%U�F�Oa�=4�� 6�ƨ�]��}e���?7���F19��I���oz��Ӟ����y"�@�Ĉ��T44_���>�o|I�b|:�J~H�3���E*VH' ���I`�����:�M���M.T�}�_z:?'P������DܥX{7��lK�SI"���^&�x�b����?S������-ĕ ΁���nҖ��Jb�N�#�������9Hվ��c�.@��D*b��wNr��[���U�|��' 1DE���*��ȕ�)�Bz5� V~:���U��ށ���N�a��u:��3�l��b����̜>��m3eaW�������B�9�B,�\ �J��V1.�J>-�X��h��m�n�Ë��;{�
� F�'����J��n{o}2{~�5¡C�s&��¨�GK3v���A���˷�Z���G���# �B��j��U#=��g��̭s=��Gٯ��G;�x��ի �j��w�Z��Z'�~�d�r~S�v���1U�,�夌�����I1�fѩ�H���nL��byQA/��(P�^S��u�v:M��
�/ɸ��B\�����5Nu��;� ��q\L��ʣ�������oA̵<el�J���I�q�"U�i��eG����>�Y���r��������ok[j$K����X��-{%�rOj<Ok��K�`���,���3v�������8P�V��:1�R���C�K��:���1���[�/^	lx��`:�z	��1=7��y/��
W��m�9\ f�m�&��y��݋Xc�n�+b�%B�3W��Md�\?=�];�������W�,\ԤO�Ë��t���-9]��CMQ_����AՀ2[�$\D���N�T�"J��)�b�o�2�IM]R�}��u@�,|_�d��ܕEu�5�i�����K�5�H
u��i+��/�ؗ�p�z!���U��E�ҽ+@l��Xb$���y�4��D}�4�F�I�ۤU��7�x�J&�XV��B�dF>K��g��p��� 6Q�ej�n����/��X��U�5b�o�#4R�]�z��12�6�ALyʔ�a���"O��n���Ĵ�W?�W
'"p��վ��y}�h>��ݣ��l�C��]�(���0"�g�)]}�#��?s��H�<���6���G�C7;)(��k@���Ԟvnx��� t3�bY*Į�5�\�q�pz�G!~&ss� ��~e|�B�踝1w)Վ�(Ī�,���1�zu��|��z���n�>��O�/=�#ޱQ݃���b&��c���cOF��Lw�e�X�KD���бO�GR6-���N�I 6%\���·T^�,�o7�Dbp���7_X�xI9���ޥ1��w����>�s#UD7���X.�������	�vϿ$w��� ���!���*8ÚF������0 �4����ڴ�R���k4�D���8tn`<��J&lo��4��q?b1��އV�C����F�x׮� �{~aD_� "�s'%�H�H��NMV7&��JG������_��o�����{W3(��{��! �����@���pc�K��2 i'�ts�e��^hs��'#���1)��;=�d]f�r�:�W&�@�o-�|���؊�I��'�%X V���p��HN����d�R�Bb�X^�<�2�S�����_���XU���ѳ7�w�^{��r$���1���<��&�EL�&"2�'�=�� �ؼhzC��Q��З*^���V'�P�J��O���O��&��Uh��J8����MӢ����"�y ֺ>���(n�=o�rXh���ĄT�!j�K�l3�< �k* F���!ZǾer�ը�vnu��rB ��\������]��l� �/�=�(�L�t!����*�b�3��SP+0֓�m���>A�A��i;�F���H�+.�%�9��1��w��=�J=R1������;�i@l����P���87�}t@&�G�͔b?�Ƃ2��՝u�Acw'6��I�A{v/�$�0ɏ*���m�����c;:~�[ olfNaC4��io�zF�6_�!_�w�Q^霍��σXs07�LN��� {��??�t���fW��dC���؛���k1QJ�A�d���;H͝���� ��J +.�Â�O�̝+���b���p~.�+���O3U���AL��5�0[��C�|Z��c�.�}�t#]$ ��jj��W��� bh%!�;�,<��Fq��O��LhA��e�21ӗ&f��]���1T>��s|uJ��w�J�ԴAL�G��̢^�2̅i��a%���o-���|�/㲰7�Jb�^��ĔX�r��8.�\����2W�X$
a^�l�uܜ�a΍��d��"�����Ș��^n>��yu<�DW%�<v 3m�d2ew��A�a�C��PJ��&)�0:�=3=F�U�<���,��z�ĺ�[֖�Β�Fw>5�܀��ff��|�*LL�iS/b/��KU\A�啋B���� 'Q��Uc}��`-��aؖ�Y��i��3U�e��ASU�%��V�6×@�bc���!�k�Ɔ�ݬ��j�ALk���¨d�����KOw+��Bqo��7�����3wzflb�wl�t�Z�n���V��陃�փ/ۨSV�}{��a���== �WxY'f���<��b���9T�rFw�;n���o��4��נ91%�س�
Զ�Yh)U�tz�M���M�5�v�z4����{�^���H�>�ߥof`�j$�o�1MQ	6{۹���B)Za��W�@��M���>օ�N�����mbO�[�rS���5�����$u1܀\�JB�N�67r�b�ʄ0+m�IDe�(ʹ�X�T�3��Ys��?�XF��?��Ng\cu��H�5&�㥕,l>a�0�M���:�Z��]��zL�j�f�5�������
��K��aך
b5����v�O������r1C�k¿�:�7��?�eܯZ�:�����a����e��B��]�g �E���h���UP�� PRB�%�iPZIQ��FQ�C@��Ii��RBi�.���3����^�����<Ba�B���G{;
 {�#r�%w�i:�N�eٝ�� 1��׾+>��C���xZ�e^B��,��l����k����1Ŭ.�N���$+b�~r�Y*�aa>�@���X�?����!5��&�Ŵ�Kk��R�s2��"�I˖z�z�Ěno���J5�Bf�5��z�!&�"�G�\���o�wԏb�U�1u���/�(�?�Go��[#@�.r���{���o$�z�W��M��;�L�Q����`��Ԕok�B,#��#��,߫�Ӫf���3Scb�zs|
��]q	����F���Al	_Y�bL��e"Bl��i�"b�Tƌ"K#=6
I���b�u@,�����)J�U����ӻ"VgUb���5�1���;DNc��bn�vU΃dS�BF��Y�?!&����wƣ;o�vrz���ާ5�B��W��u
"��� b��#���o�iH�d�%%n�K�b|Z�#��b$�׎,��O����(������B�9��l�WO�qf@���27A�b�z�xx�X���uo���6G}-����Ѫ*��r���Y��Q��
�B�*���$1�w����g0��0���� ����M����&;��(U�cKz�#k�BET)��b���T{w��m�E]��>v�>����˒Vq������159��H��?pn�қ�o�w�9�C���>�<9��C�tL�^�����1���<t������0%~�b���~�2L��'ۻ��)[��F������Q��^&��g,,�z�O��o��qR�&�͢A��TF��"�x�	V���g5��$��\���@�s��K�$�׺b� �g�g��6����*�w�jÑ���>�������_V�(�n��g��˲ob~b�\��aɨ�X.�F����7/bK5G�>�_��������6��C,�w�����i�ЛNmS!����!1�����֝�~c{�:O�e�jǶ��6���}�Q{1K��������nP=Y�q��[�05�a���W�>�
7|�����,�
M��
�?"'�~EEC-c@3p)����+U������?����*�A;&�n�W����6Ė�c���%(�cb�\�t@��Q��u�j��J���n�Z!&m����m3#��ͫ�?zc�ޥOCl�M��b2�޳
F��B_Տ# +��Զڵ�v���u\�71�XKb���\y���J�5%ξ�m���H�G�~vǳ�����6����	bA�/)�[����^LJ�dQ�A���T�a�v�A�S�J�]���w!&���a��;�t섒W�yY>3bKm\�ތ��lc��煵�j�S<���֌5r�)�����q�O�1�w��z��3�}����Уf!��4}3&H@3U���g�2��|Q7���\/�P{���bE�}H1�����E^	ͺDe��~��S
7�V��
g'��wA�6%l��1�3fJ���U�h.�ź�z��B��������C˥�>ɶh��6�<ļ�f*����_W�� T�@�<p)@t�(}� �)��}bt/I�\Ww�`�L�vӍ&"C�m⁯Y�P� s!��5w'cb�1�v���\��1<*�����A������k�U���\� [�9�*��}Gy!���&�%~p�MY���	䞗qK��qa˙fR��D6͏��#;Ԭ�Q	��n��{�L��)^����������AL�vj�r�����V�Y��)�by9
�j����I^u�TYّCl7a�e�i�s�eJ���	H3�̸���k���1A8��v���m���"?�Fcj�䛧e�J�"=�*jܛ`ݶ��V�M������S���f!������@l�K�#7�z�.!�9�]Q��/�}�u�|����K��u6w}���j��boq;X�T�~��[���E��̶��h5k�ϰU�h4��kx)�� �(�������A�"Պ�
�����zs���u5Z��W8r�XG�P���>�$j��ݧ�	�(z�]o!����Ҙm�کw��b��4f�.�K���eZ/�Y�h!&/q�p�r*�@�_'��g�$��b�$��)I�sMo�U��H�|�Xv��};��`���%���������_a����#!Ɏ���V���n	V7FK�Y{z!�Q�m���w�5�'������;&i��U��@�]oܐ��pNj�!��|�m�bm)"M&p?"�v��O��WB��<Y���UⶤΈ�{\mļVZtn��s̰�,ND��Y�XV"~�ן�I��q��ݭ~@L$�a�p!ˢ�%�:�B�b���H�6�پI�do���@�m|��m�VM�D�._+����D��d�x��{=��}>��0�ض�u����_�u�S�-�ꈫ[���8�QWe:7�d����:�#ꀘ��偧F���{�)]�*N�&�k���3�{;��q�s폋4�1���-��wL�kU��n��q�?& �0�G|�ٵ����L �}|�����sf-�D��{*%w�b��^RC���A�uo��	WU���]�e�p�&i�%!S�ݼ}�}�w��Zχ��p2�4IS�8�B��.�/�af3�ʏ�ug5����۷桷�˙��EF<\}Mm-~�7���p������*=��Y��Lٛ����Y��a�t*DN�!&�\�������jtp��`Y�b��d��oG�	�����u떆X��
C!B�pL��s\.5�����L�f��b���:��A<�b$B'���Yt��O����Mhh� �L�F@0B?��T��=�:Mjb�LM�Z�H
����V'xl�C,�KA2ڴ=G	-����_3nb�X�/�VO������J֩G@���Lʇϸ0�c�8�	
��]_����d�l��־<=�u6P5��B��"{i�n�5e߸"�A	�ܽgg�b:�r�o3��9�b ��.w��l6������ی!b(ǁ��u|W�9Z]�����?��b?�6~�6�Jڔ����3x �b>�G�D"3,������Cl
I{���g�dL:�Me3�p�-�����ԯ�pk�PU[�����1�_E����¼��'y��S#�)�
��t����ސ{���,Ii]\��5���Q�W�h�[��Y_F_�Pߵ������`���&�)9���{t�4�p��pK1w�ߡ/)7�ڭs���{% �j.Ji�'�7�|�:#�����\�@Τ�?�n5�aE}�1y�^f�	���$Vl_&UB1���;���o��n�Z��Ĉc��j�X��e�QN�6�G���d('�C')�J����O����֫`{���C�MV��Z�V�t�SU!�WK+a�>Ĝ��b��[ElF�����s����C�+��N��
���k���/��my)�R��~��7��K1���UY���2_L6L��E���������#Җuj��	��o�������mRX\��h����V����ػ�3�'���S���A�eѰ�U<���7��c�Y=9Og!bE�#�R�qs��~�"yl��^1z�"��g�^+�d/�O�)�m�!��3�[��8�����w� �3�4���VT]
\~�O,��71b� b��	b��1ş�����j�ؘ��n��~�=�O�d�Av�Z� �2 �!͇��Y>?��8
U��bAV�hTe��W����E��JC� ^��]�eN�4���K���zf��ο��KYf?*�cv��>��12N-�'�qT��h�ܩ-~C$���f��U���ܖt�r������\=�������.�F�b���gn/6�y4�i�g�,V�AL�N��Nx����c����Ά}���k0۽�n"�������b�:8(-�{���V�����sN�dsy��2H���ꗯn�*�n�>Ť�����I��ܵ�x�O�ǃ�Q��:�B?����'Z� ���sQ̃YS.'�ʑQ����
b��l��m�^�E>���f�``b#�"]�Gf�Q���($Lw* �jd���`V�5�9!$'<\KibJI����E�6*�WV�.@-r�ϟ3��ְ��C�Qb�ECvIY6�r��n�,S+���T��Y���l����Z�2��e�����h#�5'5��7������I��wL"��dr�?����8Y���9�&E��r�x�����׺g8
ʄ/j���	�{0 F������}!7�\Z5t�^�h*�R�ƦP~>j����5O�1˘ﲥ�~MW(��L�,G?��!V������2���r��s2��uc�YTwU�n�&�R��{⮵� ���ݗ6C8�϶��N�Cd=���#�L��k�����1�W��5u�t�̚�d�oq��OgD�T1{��*D�H����?�iM�l��ݧ�V�ø\�-� 1�j9��_<��<b
A��O� &��j���U�W"w��f%n�\�A�
������F�����!�J�Ծ�c�ҳݿOel��@�)���vw6�e��=���]������71)ĦfO�D���.p��!���=�7|$���j��Ӽc	�OA�gwi�}Q�)�h1b��d1�g9�a_���+��.	W1o�Cl�i	�Ȁ��jꒀTTz���M FI���o����҇�\�a�Ʀ�� 6�7�G�Ƣ�͸��u�4��J b���S�s���֚*�E>���CL1�fi�)�*�e��HN�(��|��~N��SP/6f�a���z}�v/:��Fn�,{>�Z|�"�'M�s0�)Y��U�w� v�D�֓8C�����$�Zb���M��Ak��SȺ�g�G��&���G���@\�8˵U
;��j+�5�0�)n?0�|��v�1�<\U�#F���?����]��5���15!�n��Q��3��2��{tTѨ�*%'��ө��!C��J˭�1.�;=�x���X��QCi� F��z����k�����GՊ3з3a�(%[}ɛ����`�7k�CW�%9=a�eo�%I����!V`�}�/�' b����/v{GZ�b�)2#�Îc=�	�V蓝�lS���9CW���O��8Ng£�?,��5���߄c�v��I{��}t>�$���g��lF�|���Iq��J#.M�
բ�ǤV3�Rrt��%P~{���qZ�P�@�,��w<�����+f쉩6[�f��q��*��˱p�qϻ�� &�����`M{(69(E}.��
��g��~و5&> �Lj�g`����;mV�=s����]�~�����0���iP;yf�oc�rbIt�bS������).���D*�o�<��̤{�@Ĳ�N���ҔTq��;Z�UB,HW�[Y��*}U�2�.�
�=��I��h�h�U,��`8y?1O��!���h��s�kv�eO�Z�[��f� �M�.�Y֧s��L��1���C�3|�A�zԈ!C1��#_�/��u>	�;7C����E��ؿ �X�h���w8|� `��:dd�H����g"{'{D�8�&����ޅ��1�Wddk_�u=�{��������;a����x�����fB�[��Z M�㶥�����(rrR
W��5����i�7�xR�����X�ɭ���Ʉ�w,RKݻM��`9ۃ��kݸ��{:�~���=��X�?��5�Ԯ�x5-�jI�uA�T��}��ݙ�s�6�e�U��߶�o�l�����z���!C�g���b��.�&L7l�%�	-E��v�DW�溍�DSg.�s�<'$y���E�X�깖�2��t���C��Fy�~�����2]��78�\�!?������f̌H-944%�5���q ���뻊���M�M�Sb�#�tU�'�!���cSN��$�v[w|��Q#�h�fנ����,��M�7x�F��^\s�"K�rH��� .�о\�ĈT�aĀ��n�����p
�H|R0_W?L���4�� b��"?X�Th��j�����
'$��2/{�!1;,$�m�r����",���/X��O�5�4c�q��%Mk�g�������@Nw��q+hĪ����\�����8R_Գ3|>���i j^%[�>+�S~$-�^v��_��_������K=����>����bCZ3���D.�G�k!5���� &t���{���ਚE�� b�Fd9ÂU�r:���k=VD] �����ᶾ��ɇ��8F_��&Xg����?�`{�|u���ĎЃ�D�I�0��'
==�A��1��-z�&l����G�|��m�YA�g�"BbZ����=,�S����[�p����]���ƊN�[?-���!vLe�C=��6!��	1s�>E�\�SԘ?g�ͮ�~�bkJK�����Yo}����y/A��[/,���6G"��d��(��\b�=6Q��Փ�^
iDd.�e���54�Ha�	�I�1԰"��o����&���i}�4喟�0(xG��ǋ�=Q�o{�����/�����Nn�ö���GnU��9�07���)G��b�c?��t��Ǚͧ�+��_k�0Ո2S�4K����M̍���x���:�WQ{$%� V[eEN��4|��Ee����7/�_��o���;G}���栎ի�.���a�`1�N�G��N#�=���
�Շ �,��"r}|'Y-���(��D��L�Z�_�E�ș
�g�F�L&�Xy�������v��X�e��������P��%�����\0�K��GW������Q������a\�1բ�3#q���ic���-�l��ﻝ�<U-���@T��ur�=�����-nu�R��]�}�1�N b��}sϞ���l����e��A@L3�8�h*��8Ev\��� bd�~\�'�!g+rC>7g.X�%����Q�M�|��zg$@T��J�~��0�$,��P�Rk�մ��ȁ�������+�}��0;o
�0�QB�J�d�Ą�3?O����g|@���VH���Ȋ`��U�4�mC�������p�,p�h���b�g11>��G��̧����G�Ux�@L+_��\ް�0�{��w3h��z �:�U>��0Mr��+��,R�o[�`Ǘ=
�U�nu��Ů��ebΰ�~�}�o+v��=�N�/1�x���1��B	��2��Z��A�9�)M *ee�8"k���˭6���V�1 f��pR+�0]e!�\/�X�����	����~��a黢�4*Do����M�{ph//�������aZ�'syG�o{s����$�D/�� �dŦ}-W�W%��Où`T�3!����FB��,E:����7$N y�Z�%? ��e�I���8Zߍ>^V2�h^e�Z�b��*�����-M{a�}��Z VwB��`� �監I�([o5�1������H+�}�R��'(I ��\�.�?�{�s[<4��nO,��u�5¶�������-�#s1�Z,΢��!�o�|˯U�pA�ld��Aj�X���G�-�l��fd�\����8��.�eG�,O�v�F~�����S�b-�2g�����A� ���qÇ�-���֑OQ��$⑚K)�&�#C9��d&�A�=�s��q:]nU9t�0!�S����G��"�#o�E��<F�{�C�v?oad�2-Y��T~��۲�?����f����ɱH�ص�i��3Ψ@��E��g���m����}�zj���;%�Pѳ��H���aR��˾h�FU�^�x[.-�|M#*��4��U�n�������(�`�pt�X�'�R���7�{�B��Ǭ�����~S�F/�Ĕ�6�;�������̝������֢�g�!4�o>�1��<L�e���{���0�u{T��֔�j�B�q�s�z�/V�f����Fy!�4��wm[jO2b--���WS�f�:iZ<�FɣY@�%��ݨ�Rϩ��'��[�Fb�8+�D��)un"���(Ks�z|ϢZ�BV������ř�����N�Ԉ���g�5�ꯖRee�؃@��*Q��75�6`|KIi� f��D�ߊS4��)>��I��ɋĖ��BDK�°E��i�o�ށ���������h-�Ū��+�s� 6�{��=�~%'�J�乷$AH2����kd�S��a8���NAL�����i��=z�<�bQL�(v�RP��s,��B�r�TEZy�N����W����2����Yi
M�q���*܏E֏�.1��}�2�gcE���V����� F����=h��c䝦P�n��MV#*����l)N�������*�_����'�އ	y��Gnl\�߿$��n}�z����Me�y���ѻG/ �8�B�� 6s���@GËZ�����֬~�_��_v�Uaf�Ǫ*UR�3AZ���9r;���6;No���j��]mS��1�zT�������$����@�M��z�Qq(�>4��b(nz�3UH�T���4^�-w��q8C�d&�S������Wk�� �n�Q����o�BJ�7<�geb��?�N?�>9��l����ݣ��P�`[vChԓ��!��f�* f��H$t�׸s�Y��-w'P1~�*�\�x��_/�ۃ�� v �}��
N1n�##[�Zs$�]b�{f�W��D�l�l`W���&��X�ES��A(�(5]��@S�fcd�]�j�{t:��(Әb�X��v_7��[�C���	'��� �+��.w��W���Tk���q�%��=���*��l�Ϯ�[i������3����AS��,�8��i�^0ӟ��wO�@��j:��I�CT�<ZD*㪇��ǀN�Ekh�W�pcŁ'����xKT�Z1���	N[���f��.>\9�z�&-�Ģ��� �r���"�ux��ӥ���XqJh���cv�d�R���r�*�/R��1e�c��#�;N}bXL4�E��n���j(�/Y�А�Al6n=�\���S��"��QiU
�l�?�uX�vh�a�c��� 1G]FU�ڵ@��7h�ɜ?]tA1d�[���9D"�wHHWAL� _��]�M�����L�E3���'��P�b��d�_���s����LL���Y��p�w
��*�?�(��1澧�Z�{zbH[�D�<�Kqv2}�fy׍��X@P�z�S)����s��M��AL"���+[*��a�C*�;�b���w�}J$�r̗��Hhl�#_0�?�԰�ܞ����wc�Y�b\�/ v+@���k�9�.�N�����qϬ-o>��6�_N��'��Ĕ���&z3�;��oUjU��%u&�s�t�d	�Sk�z�}+:�,JH-v�A쀦��PE�-b�Fr����T��}��>F;�2��I�	�l\�k� 1�Q�WسC
��=����8H �7 v�OAL^��۬m��	>�'���J�����%�^q}i�ii��o9`�Ÿ���Q\I�OC���~J��\���I#Y5:d-�Mo<�������KA��e�����G=|{�3�����E����%���W}��3]<���N��"�A����S�˘�c��Z n��=#�������ꓻ:YF��p��\�`��d�����cp�-2Ϭ�@��BS��M���@Ni*��J�U�U5�K[�5r����'�u�:�J� �N�P�+?h?��%��-����0�no-�!ex?ū2���y9ӈ���O$E����N_��I���:�6`��=���+
�u~1�K��n��s�����x�����%v�wFڰ��+��"�߶)��&'�8{�?b�Pe]��;��Wg.�b��K|iQ�ЛQYB�R4@�����j~��_T�P������~9���4&�1f,F�n3V�L�Ɂ�_���{����xA*T&�M��o����x�a����͵6��S?��
b�v�%��~=nD����U�R�7@%���vzڂ�`�W�]�&U/@��U�f�q�#�`�c���s�o��G]%g=-H�Uʖ2r���ؕ0 �"K�i�֕�f��x��"W�X���W���mm��&��
6�6��g�>��e�d�(11�z ��?���͒�2�o�̟��ѳ�Q}1�������p� wS(�Ua�Ik��>�我N��u`JǄ��Ȭ��ux S��:鞝�KWKeALP�h�T�z����""������LK�/�l�w�]ѻS����*I��<�'7^�D��*Cw��%�Al- ���-E;<RU6��x��6� ST�T?<DG�x����y��Z�Nx�$�|X����ϯ�قX�v7�i�.����)˳��� 61��Ds���&�&�����2��\ӕ4�y���}r!�hY�������	�Lg��[�����%g@�b�Mz{-]�g�=V�mŝϾ�!@l�,��m��i��`ޏw��s�@l���)2���i7�t��LP��m.�i�f J2��+��Նt<�"69@�PU}��dʹB��g"���9� �bÞGA���~r� �Nǐ$s�#����3�z��d�I�=0����i���eO�O+Z`�NѸ����~��Nq�7�Bυl��\�<�����+����b�?2��ELR��%��]��fQ�@���v��U��G�WO9@̰L����-hb[�~�O�4OĨ�<���(����G��� l�Al_9��Ŝ����A���<כ F=7�S��8��k��(����b-�{qC���q�ܮ啵���; �E?�t ����g��/��U�����AHy��	A�f��R��M�A,�;�%_�Pz����T+ �їB��9��4o.�D�h���[����6��2�f4ԝY�O�d�y�2� b��R���,;�A�1f�c�s ��B���D���,{7��@�c�_`6?_�g􈲾3�B&������w�B���e��c3ALdT�?%7�9jt��G�
GWG[�P-c�ITQ�˿e?t�\ 'b<yX�mS�-Q���1�!3F9I���?�Q����(�ٸcL�`ק8#*�6�@��06D���.Wd��Jrý�︼�e5e�ŧ�:O�1n���
�]~SsީlS�KL*����˩�o[;�`���OY�N2nz�{<���޹����f �I�}��vU�3wR�g;c�� vD}���j�>��/��f;S �W7����\i�gVE4-3�e�Q�EX���*=��HYK��Gn5�ؚ3�hx�O�@u�L,�>f�4��P�Ih����S���q���.)��FA�[�^RJA�y�Ii$A@������ݙ�;�����g���$n:#�Vͭ�����q�S���1ʹ�Ͼ�	�f���wC}�U�����܄����^���ɗͪ�Y��.��º����ˀ*%����t��y�V�Ul�q�͈�y�2�X���r��"�!t�c����A���*,�����W��F�3��d1�0�
łT����8Wq,���@L!�,�m����_; �M�:Ī�K�	�n�Ů��܃d��}@LJ�����b0����a\�����%�=�������:7��$�E�b���1�(�p̹�)\b�`������E__��e��W0bő��9˿1-�Ϋ�=��{xӚv�{?;S3w�~�
�ᶁ��B�/J�r���ݑ¢@��_ުYC.��vL%���<k�?�U��M����X�aQb�'v���VY�,���`q]����i��]沩�|o�!$�&���AE����Mw7�&���+2��z�vʇG���,M;��{+bC���[F������B�ܫ�1'	�	�áKa��sdv#k}��V}k��J�s(��	���N�����S���ƭ	�̼�7rC)'�I%����dW�_`�X�������V��ѥ�L��Ӕ F� ���	���+^�e�ˆ-1;��)�\��qw���.囦�s�t��K?��ڌ������wURu�~�ꍟ��F��`
/����}?��R�����\��� �����,�r�����yǲK��ا?uJ��Ӣ���,�ũ�cpgF@��d���b!�"ʪ�6I���R�b}��8�����8�3�g!f�ذԝ��y[����ވ]���'[��w��?��$9�LyI�4ޘ��q�ä��O�vEM��8�A����c�c}�DDK#����9��_V������W�%y�}�s��}�"}��G.W#]>��e���5u(������!c
b��?��sG_R^�M����7���{�gzM�~g�\9NVRA� ��V�v��y?��=�Q�Kم�3�	�-����Ɵ]^���P��0��>�X�X''���k�61a�d�� 5�
/��	�(�Em�VY$	+0�Rz�h��1lU�*!�Yc�@l5�
�>�YР5L�b����7��4�,�MKb��{i�eR<�;h#��NU�����J|� n�$&nO�`�Mܐ�x=���]�u�U�������
U��1T?��h93�\a��0��9�F���k/�X~o��,�����W8vĕo���Ǔ܉�Z�<c@L'�����d�a�-re~�L�Q}}������+!�W�rSbO���Lʗ�G�"*��>(@F>�»��G�Ϡ@WQ��T�	b�9j��u{���X�~��H@S�AlBH���k���Ok0[���GI� �����v5��x}���3�|-��j��ӥ=3�+����R���1�⽱��r�c�	U=�@~&��]��d]Xm|�PlG!�L����8�;;[<�{�4���k#�9]�l�d�뉿���}� 6b�f!Xv���a��+�3D] f��	��շ,5��2�sIkNi1��W�s��U������������ي|f�T9�	�(C����W�d5O�z�]y1)��+:1ƃX����f�y���O�{1�7 6����@n┒"rz�1���Ldb"�
���¸glXhȾ)* �{#�[/:#�9����it���n�ڹ_���ܝ:`�����X4c�7!��|s׳#�����A��oκ���g���O�V(� �=o�Db脽]6���Ra�}
b���bgK�I���6-��)F� F���Z�U���"�@� ���I�6N���^��K�-�{���1d+���/|8eM�HpGr88�T V12"��0@��_d:ܒ�W!?�Qu;��<�-0(i���'�c��G�I��$�s:2�CQ�"�B�� �:u�Xu�Q���)�b��&�8��9���0˹v�f��$[��z?W�G��wv�$d���"�S9���[\��ļXj˫��ŵ��7;�O}b�7F�6�Q�Toe�b���r8�rȟK��W���AL#ښ5Ǻ�3�@!�|���]� ���;|Ox�5��%1�f����Y�J,��zW�9�C~[�K�[���Tϧ���4B�@,V�壘��������[��ۜ[![5�m�9\c�M���Q���oİ�_��h�l+3��k��#~.���/���=b�3��IHp���T&@l����L�v��I�s|9����26��8�o���1ԌOGb�50#Z(d�sp����|�5Q ���=+�����:��[�X����l�?�@�PQ�e�����Ǹ��2 6�j��Y������]��H|^~|��ݐr&����q+�p��؂ؽ��K6h��ia�a��;,wS#ܾW�>�{�h�ʖg5�ed�n b�-�4�6�0���	��H'�!� FS˝5%���=c)��:-�\�>�_6�O�ҵF�u�v����G�l��V���g��$*��򒈥4S��h��Xu'+c����8b_P�9���@Lױ�3���S�� �_N�� ��8���_��,���d�E�{���X\63�.�ᗳ��Q1,�0�EA���ؚ��k��@Pn1����1-�0"g��s�š����xB�A�*9���)�r��r����"�Z��R��i��R���������~�6s�E���[�m7�����!fĉ�<�
'��g)j.��1	��]��D���8�u��t�}=���
���y�C�M��Nq`��dϮevQ��!�������yJq���L&f�n�E9�m�,��"a芺DEO�^�,�'�X�5+3��S�C��<<K�e�8���S	�r�◶O���}��H��)����	T9�(U����_-r�tg���Rm���X���"׼\�=�Hh���M6k�L���q$BD©�m[��b�����f1���3��A��|i�I F��1\�O4��{��}��n�����R9?m٫�̦�,���"����N<fy)z0G���@�����s*2�S����.��D� c�n�am��~^*��A�Pb��J=�>��4nD����Xb
� �e?��F�,~�X��x�>���}�<��G��e�����X����M����u�1@j���j��Ӿ`~ؓp	 ���7�r��1I�� ~m����>{V�s��B�7[OI&�W�D��8��X��d5�F֊��e���~��3K��D�qS��UR{��k́�j}�,b�``=�-L�JW��l����DW���\�칢�+�0��C���t{�N-��S�}����~*�e3���?�샄�U-R�r����a^7�3#��d��V}�b�=��2�8F���>���GS�Xb	��$8��}K��<A�
.L(��
&��gaϪ%����y��ӹbH^�3�1G�+�Wl!���P�0�?C\J��+鵘}��*ӒLh�ǡ|��&=��V�	]G:��a*G���߷���I$�!�1��!ˁ<���a�:}��̰��A��r`z£��a����Y�>�)����vy�ջt���[�g=� �����Z^3x�΍�S�یX[���+@R���ʦ���Z�L�����|��x�o����Z�f@�:��,"�Ru��`%�g�B��YA�{�?ՇV�5�1:="\��h�7����`\h-ϋ������μ&��^�<��n�0v�po���FS����֩�q��!�义��̚���g��LwƊ����)7����@@̄��[��g�N������Њ(use[�/�zp5�.���0�	��,�O�_�X��]�C��ϓ�%�@����=/����c>�R۵K<�&��}�5�|B�F���\ߣ��4ͥ?��5�u)���氱��V��z�b�8���Ok��F�Mu�����܀��U�
��	�x�SVfѥ�6�M$��X�l1�W��K�ۄB@Lz�FɎ����}v��8	��f=�1`��M�I����9�q��#�X�A�q�E�P�?�/t=i.P��h��	 ْt��~o�۾�~�bx�⍃��ʺ:Э�������hi�m�i��������cH1o�L���8�;�Z�~��ڃ7���n���\��6zS�CY�r�8b8�2��~�a������,��}��bKq�sI�~#��L?J�[<h@�mY�N�υ���� �'w�k�u�?�r�{P�*�]4�My�X�㧑;��A�MjU�߄��� 6gf��Q�'�������+0��w)W�ն�@�Y�N?#6��XfK����l�n�^��c���
��{�P/�j�ޗH�j��������i�u�T��n$y���O�8S뭁X��R�;���+����oT�zY@l���*�Ѫ*c��U���`v�ĠҭC�F�	�Tuخ����� fS #H�����J�a��?�n�^�Sq�Q�uv�]t�C3Al��CY�5�7�79�Ż���2@L�>�oe�AO!�ˋ�7Ĩ�:��\jZ�d*�����CE#@,+�Ҕy��$0��;(��m���Hu^��dY=���x�Eb�3��]�g��x��Cw�pA�ھf�F�(|b��D�ȣ���J�S�Wd���y�\��BXaA�.��^0AM���M���ɀC���}��2�ɮĹ~q����hQ��=��y�j�|4�;�F=
b;C��l�	s��'i�׼A���Xj�t@y�J����E&��a6K&���<���eU֕=�H�EH����B38H�Kw�i�$����X釳>��$���Kڞ�L�b���<xS�V�9Ʀɉ8�q �B�$pY1��T0�N���t�ĔK[n�Jn��괸�+g��X�a	U�ɘ�����,��k��я ��e����rl�>��+�/�G�Xq��j�
��\}c��B<,z�7�=	�{�-����S��c*k@7�����W?󾒓�r�f �T1_���C�W6�
վo�6�@�.W:Lϙ3,]�^h�B%2ݡ���h5��Vv����k�Br�zkA�ۜ$s�v�7��)V�O���|u�C��V$�k�Z����� �����[e��mΉ�#�]���9�-I%*W��������u���61<}�� ���'s;�i�zx+ f�R�/��0.��4��"P57�Į42��MR\)z�3�\�' &O�O���+�]�źfM�Ƅ��4:��9;�9�w<���M֑�ih$Z7�ѯ�Ƚ#ӁZ���Se!��8Ǝ,� 1|_�����y.�*��{�"8�(ɿ'?���#�I;�uK������p�m��T���@3b����G�<�E����$�%C���s��5�����W�2b�:m�%�#L?�����zq�4��U��6�	�o>F'�/��1�@l��!�f�rae�1aH�G Ħic'�#5��V/���+D���@̀�J�Ŋ�5�`�E�I�0���/�F�Gh���w<z� pٲ�M�B�t�-{d��q�Yd��MD���"[���d+3{���t�}�۹������-� +&�$h,u��������" k���z�Hc����HJ�u���TKM_J���iԼ�m �E�~b��g;2{��nf�)cļ���d �jK������k?�y�(�����ʰ�ҩt�Nn4�%�|+��1�.�����ʆ���`ߺsAL53�ꟍ��YD��(�an����{<+?��J-MG��G�Ҁi5��;�qI}�MoRFؖ"�;�ɗ�G���Rg��D]�}$�Q�1^�Ζ��RfZD2�kwqH�A�+LH��)�����p$�R�\�	���{�Q�?H�y\�:0g���C�w���Ӻ�zs�F�u�0=9���D�Mz�4ύ]9դO��2��zݒ�YzQ�����&��N�C��AߴK��s���-�Mi�h���W˷�1��Q�.?��T�1q���3J���m����:ȓZ�����[w~�����m��Z���Vk��p����A���b� f�H'��ٚ�ᘽ��;k�� 
�\�j�|�>,��d�UG���b�1�(C��lӗd)\�-F8/@,[̉Z'/	�".���1����b��v�m�̱�8����u�>��$�j9��o9���ݵ�F�\m �PI�tc�*����`��8�G%��>7Ì��P<P7����Uhaw�@l�����9k&�KaӖ��6}b�.�,�&C�h�2����&N� y�_F�]����>� $���Ć�^�V�a'�JO�'N<��3K 1N����{G��Lb���A�%ڏ�6�[�U��Ҏ+E֯@Lf���_5�\�+�Ll�+���
b��q�#�(OЊ�l�q��ѱo�����6	��!�����uӔ &��i5Î;Ϭ�d�!��q^�b� ���K�K��3,�G�: F6�@���1H�������yĬx��#��团z8�Y�q'A��K�k�U��'�
���U�� �����ֱ�>PXL�!;6�Ĩ#�� Mϫ��.�Mx�*�X�ѝ4f��n����_�I���F@��]w�� V��ĸ�җ3ő�zFoq5쮣RV���#�7� ����WEN�:L�=���bS9*�'�����Z�P��|��b�Y���	��g�� �ꆸ��M�.����Z؁ F�K�g�۟�r��3�E����1�y��Ht��_0IW���X5�wX��=�l{֎�z��U��$G��X_",`��j>\W��ILe�1��\rl�M�m�y#r���̟��6W�?���\!n0F1����><7w+�9r�.I4S{��%��+ka�3qϱ�������]~�ʷq��n_a疠L|d!b�Y������v�	��v32�e���9u/�%�f�);=iI	��=A�v�;�VqbS_��萄}��#�?�Ipz��W���~���#b^����/�'�!���]'H� ����z"��l�T�?S%�>��gMݫ}�|�*or�6s�� ��J���9���v��U����b���KV_rvT���Q�W��kAlْ}HE�[iE����S&�T�.Rc�,�tC����R���8� ߒʘZR���H���3�����t�vrWi��u�+��ٺ6�љ?hC����=Ê,p��M���t��k-�^����WLA�eȁ䦐�m����~:�#]W��P������$�x�����(MĢ�f�aR[m�-W_�j>���b�l�,��9ݭðJdysz�V�Fb�.��Ұ�ދ�0�ȭEVQ�����V�����L��=����U(RO�i�J�*7m6���{�˶�K�م�Z��rtU�@l� Op"*��R2��-7U�l�P(���mv��9{���$��h�D�E�^�Y�{�,�r��d�J &B?�1*�;��?H⦫p����ަ��[5%d��E���JZ�W�'*0����!�N!;C9��{2��"�BvG���V�6�u㫫�E�/�2XR�l)��T 1�.Y[��AEb��gR����y� &F )�>{=����D��Ya](�Y>E��8-^����/���yĐ9��K,��5e>dh����?T�}U����W�k��s�f ���\� [U2����7�!Y���B�Q��)�>���ٷ�s���!�bb���Jӻ�?�2s���]FU������ߖs$���=�]|�z bS��`�a��Yy��͈�������!a�f�K!D�����m}�� vu3i��b-=��Z�3��}�%k��:l6�cys�Q�j'�X~���~���V����m�Psw$�v��.���y&�m�N��Ǝ��4f��q_V�9���1�f����)T���PB����tA�����;o��SM�av�[I�0��GQ� �������ַ�Z��A@,3XS���ĬG�e��`1�ϵ��xD�4����ۖڰ=�7;(d��[���)�#/}ݓK%����@�y�{,,l?�BҤ*=���A
K�25��6H@��ے�HaC�b������<I�b.�$��A,�L�V5o_�S���"�[� ���J�a��m��͉��FU�_|�1�/���K܆�1��J�qZ3A��X��$���s��JaS�
C) v��>����*?о%ٔr�1��
*��-�q��ݦg5IV����F�Q�*/+a�A/�@�?Aߏ9����n�g��� &6���U�Tx�j~�,��b�:����ɧ颛=��~���M�An�~�^}l=��d��.�6{��}z��پ�x�U��4��]:�S>٪qܼA��	b{���WX}�G���&Ѝ���@,9�4o�h5�ַ��tt/��M�ai7���@�G��T��n�����i�쇡a�ˠ칃\��&S�7� F�v��
��a�W���<n%��� �w�,_YRy�P���{q�pa�|�朞��C�G ��:���� �d�}��T�jo�<��8b\��^�*-����\��~K�+�Ć=�{��L��(0��1����ybJ}քt��'��EKi����p+�4�g!��1��\W��Зk*XF��nA[Yh��4]���m������X�q�>wJ��%�y	�v�1g5�4Y<��®cr��<ԣI�$=8٠��.����Z��'�S���d��f��j�{7[�L6R5���Iñ�~^(��Z�&�1C�*�k��G V��*7�<�0��0���6�w��,u���Z�Eʘ��;S�ղ� v�`oC�Xz��e��Gg���i�y��/��gA�,��A��ua���3V�@���^�y�a	���ˡ$3��O��~<�e�ӑx��F33��5����MK����v9�ۣQ^}݉
��ߌ3��E�|�U�����q� &�`B�jd��:{�>_x?%0u�P5�b`(�_v:N�[��z��>����ak��gS�*�%u�N�s��f���F� ��VC~�SG@\	����xC�����%��2R	3�FWI}��T�E��P�v
�_Z=���Z��2c�I�����s�1~�X5�����ɡ���)I�/�ù����d"o8��!�Z�>�U���.�7/�� ���:�e����x��l��`L��	ށ�T�i�M���A�a�k����K���>�~��g�������Q�Q��1�H-�h8���Ä6B���)bm�`[U�l���~�$�\�nӌ?|13�i~�y�''I�����aۦ�ߨM����7]}��R�1"
�����<U��H���/�I
b*�k��4�58Y���u�U��l�h�߭��w� ���dh5G��&�*�� ��Kc[Oy�ae.�T�G	ӥxFV v-]���z�N?��>��9�cc�u��	R�3Xܿ>�<|u^�"�_?ǌ�C$?3Y��#
��*���|��M�N�u�`i�8xmqрW�g����5�,��5�s˝_��?�A|�].	jS���u.F9�	[�tإD�q,�=��m��D�cM����=����<[rk�x�@?�1}1^Y�>����|�������jY���݈دPe��~�K�'0sŎ��rtX��q��&�=\�
��/��7K��\	��Mj�1Vtr�ˣ��r�?�����v�[^�1�:~���}�nm��m��xA���;; ��/ه���0G]��������t4�LcU"Am��^p�n#�A�m@3���ǸX)��ߞB�:+9��b^��U�|yx�Ὶ�_&�c�-��zj�n�J���̽���T-�'�F���iU�?F@��G�QޫP��<��2�����u�-�D�P��܍�X$+e��Ê��.#`�|%9p��<H�?g�wK��?���N>%vi/;	��2����Pv��$�1x�9��!��m$0�-h��M�c0������1T����V`1�r�}b��Nӊ9�8��2���Z����-�gC��d�S�I�1�����*�qW�qg����I�L�C��<	D˯%�j��Yc���r�PM���w�1�	:k�����|����+a�錝ɉ����#�$�[ &`��y4����v�9��6w�n�o6��|:�]9��d��hO������	@�-#����Ew-�[�}J���N�����;O�2/�X��zj*ٿ������/%� Q=�\�,�4t1Kn�&�Ħ�}�'j�"i��2B���d�5��EC�nI�N�&��Ï�e�%�����A��k�R�׵(�cM�J�..R ���1'Iy����pO�j�<���bj�cy���*.�L\
��λ�f�p����~Nm�L�ʳOc)B`�&�ĸ�Sո�e��EOg�*�X�.fy����W����|�`�cC�6��o�4�L�mK]y����^N+2��$�2��;ُW٬�����X.ùB�!Zs]V�k2�A��)�l`Eh�3m�!����QiId����?VH��0A�Z�G޷`$o���b�0�����N.�9���Z��A�yX_rǅ'UI�c����i�Zw��f@N�A)7�ع�PU8�b
bC�!C)N���xI�\t����5[���X��<% Z����T7��Q�㍅<v{�8�M��|V���7�c��t�� �!E,ҭtL̩���:S���Ҵڌ����j7H/���L1S�=g���n�.�����$GH<��@�6̱c���b~�8	o���^·bZ���=�fX%�̫#�n�o�8�?_k>�C>W[�f�>��b���沕݌���������ۿ3����u�[���=�nG��rP�1ѫ56҂O�fٛ�0Ky:@�x���KTR9�f�-�K"�*�{C5�W?A��ܕ���ϖb���n���Z�BC�����@l�p��[���{�D�-�U۷' v��,`�U�_���������?�
��l�zYr8#DB��ӭ�X��b}w.��4%�#���f����.��a{p��o�>���e�����V�e�8�<����6N(}x�;����攖��ƺP��n���z2�۟��baT��L3_�o�6Y��b�-*��Kf�'����"G���c������/{��wlV4�_�S���=�$�-��%��3c8���I ����K���g���~78�}�$��������G�L���X-��!��u>����:��AȓA|�	������Gc����d�����x��xj��V�	��F��|���pfa�h;�ዲ=E���Q�h���UX�چa��� �F�A@��Q�P����NA�C��FJB�E�C�w�g\�f�5���q=��c-��W�˟l=kA{��������(d�-�Y�L������xxf@��:RNk��+Y�!?�%���=Q�j����)f�!59�W"��e�j�9���������u�噩���s�slo�����i�Q$����ݢ�nT;Yy��G	qO���bAL�*z� �u� +�v���x$�Y"y8�ŕ�4g��ę���'�)�;Ƨ3�N;�4mdz6 F�S�sG^����$i�z��	�9�Q\�y`c���v������@�T<�	�mdؠ�=AL�o#Am���?�:���<>q]��#����0:,�o�Z���U9L�:<�QqZ��f�A^�Q��'bf��@i�Å�~<|�U��N4�|���8����b��s�|E�vQR�cź��/7��O��������`ExA�HA��ԝlS�I���=�����r���R�`�Ѭ���t�OǮ�?�X�2Uҳ��"��﹍��=1�
D&��#����(����A%N�PQ���WV;�gMK�֬ ��|,vk�����ԕEy��b�y6d���J��b(�O|�6·139��#��7��.[e�̢x@��\����~�M�	=2���2+��ok�^��ɑ:uݑ|��@bFcI�8�C�\82M╬<}p4 6W&U.վ�;��� ��BY�|��C�G�Z�v�Ft�+���$گ�@�(�K�D��u�\�Y~	��Ī
c��s/��SQ�c���b+�^��[	_ᛔd�i�YC럀�\�����h��[ɺ��Z V��P����g��%��5%�k���G�|4�<fS�$�L?�>$�Z�>mL%n�7�!7oy�p�u>�T��kG�:�w�S���<� f!���ܣA#c1��4�Y�� �dvR�5U�5\�'�1H��'+aĆ�/鱶��y��W v�t�n���4g���~�5�
�uc�8{�=PN�\�hY�U�.,1�"��;��,������JA��D�Kk:��F����=��vs,uv����l��{��ڼbYΛ����3ݚ}����V@,���`��`7����@*�Pq�.3�ܚ����熼cM�ҩ@b�)�uY;O=^=�T--pl� �F��t8br��ĭy�0�z�Z�ng��J�@�#$SC�� 1"H�M�F(v�|϶�h��L6�	�� rz���g|%�=:���!��j���M2ڦ��o3h�@̇�*��b7��0��V��YgVc�	rdN����%=pjh�S'ͿbEΎ"���zw��]d~A�h�}l�\~�߽�6*�Ȭ���`Ď�d�"�!�иW��8��cD�A,��iͳ��WŰE�a����P����ZϿ<@&�W�a�?��L�$��!IT}软��g�^H��Xe�gM�(|H�]H�ۡgC�'�����A�?�'�x��i\��<����79Q�E+g�ʋ�*�@leQ�|�u���1[�y]�%g� �����<���O�_'J�����bP_���;e�!V
b v���\*�ʈ�bAKE��X���:�{f��Kӟ�r_ߔ�Y%1��[C���2ˢ���!���� v����al"��?Ia���<?W�bb���"�i��v-s��'ALvx�l�D2'9W�"�lc:	�xs����ף�i�p��3�o?�b�9�պ5Ι:Y������ �jĉ.7Ϲ��A^(Du��˄�b�i=��s�s���2&���9WsgL
jP���i����P{ǧ�b�>�T)��7�T��/��$K�@,ص����������,��Ķ��a�,nu���V��yW���Q_�.���j��|^I�d������_�g
���E�-�9m��T��Z����+b�x���� g{�#�|VG-��~0f]��2�\�	�:�ޤq��XPCP~;\�Q������m���˳ޡÎ���A���~9�l|��uZ���<ܥ�T�� �|mJ����\V��<�ke��	��&�^���"��0���]3��@�de'4�#	��ee�K?��Ռ^�VDe��.�t��++����1�cO��աdi���>bL!�UC��s�٫�=��L3.����f FUNC}�a��l�H��W���F͒��R���N(A���(�M-s��(���`u$Q�b�q�22����ũ]�v��ج�؅�mⶥY�-2N>l2B�$Cy`Zt��L�ZA^��2x�3Į�Up�l�`�
���J��#A,7<,}ɶ�L��ODF5���x;Hf0>B��D�����ƲR�L�Ma�zHaz�C;d�Y&�̡��B�O�'	�K��/<d��K;8���V�\�r��$�	�����8�YV����_�>�Iؔ�&�Y$
b�ٍvB=�}?o�b�+�mFI1{��g<CF��(^iLj�TzPKs4�.��F*?t��~�E�/�b�,~��w�W�4� yўE �j�T�b9��a��_�eŔ
b�^�Hɬ�!�%ϕ�u�MA��ڕ��������sZd�1����YZEYM��/�j���M뀘BPk�QgTU��=�1{azK��2;c!��
�`Zd��<�N#ʻ�~�F���|�j�$����݋vfvk�]6l|�6��.���l��}%�\"}ʤ�VbL��R$ @���_�̾�!W�gI�}��{Gr����Co=[�Vi�]J���4|����RºO�����we�u�iZx�A����3ʑ�����ϻ���w�0c�U���Л���YC;��e�Ϳ��U)nϴ�v:֣b��7�rNT�k	���N
�a�׊�W{?��T�GŔյ�M�\���(�Pb�i�u��!�˯�M&�M�K�l�V���� �2q%�
z�*�^�L�5�SEy?�
q�*V�J�!��&��N�4*��Y��}8H���X�t��g�\�ӥU98��s�>O�h�A�82�EH.��3/OڷKw��m�6��询-<����.ÿv����g��v���{d��KO໾�6w�ڗ�(&�ƺ��fw)����;��_��t%�+T����P�ߠ∢����^P��]����*�ܽe�����y�PM��}?-n)$T��@G����;!9$a8�֠�^t;ÿ�H�C"�CJ����P�iۖ�_0�)���ӃJx�ϵ�x� ��+�
P�������^�ݓ��̸��0y�=�p��Q9�w[�A����_�[{/wu�T�،�N�ĆP��$�r���t-4e�z͝Z������>gn����,z(�� 5�Ɋ=lO�+%��S���ѓ~�K�Ô�c�1�)(��8�uw��뷾�25���r�b99}����HD*��A���!.~�)�2�e/Ì}C�]�2p|u������q�1���Y�����L�����Sk�'!TM��y6��y4�����+/X+ӆ~��e��7����ӿ����Vr���V�G��ZYXn�`گ0�j��WR���̍�fS�I�#��
�,�S����Ϥ~~%�.C*-�S�R��I�*�����.��CHl�K	���S6�� ��5���%�v�K�m7�6�t�&4E�i�&2l�Lp��b���5�I�|�e�o�b�'K"7b3#y�f����3�8��&�zʢ�ֈ��A\\�;��,*B�����1���y��~{Ҹ!��G���h��yRz L;�>�E���p�����/X��U�m�(�R�PD�-V��覩<g�8��7�{�p.ݱݎ}���{����]ct��è,�`[W>o8�W�D��f���[�n���5N!�5��Ti"
WlO4泛P'4"6�cA
:{ƍ��З�Nw{}�"S�Ɉ�հ��4(����e)pv�K����c�8#G�*4$gV��̅���&��C��^�n�r�����0|��]e�h�j\�/o��{w��:*���a�B�%�N*�E:\���H�����W'���^��o�ђ���Њ���_�ov��N�=g��c�V���t����]�X������^�x��{
��a��9~�J؊1	��0�P?S������}�2Z��Ĕ-O:��v�!��Tľ�<��
��Ln��!fn!FD�Q�����&��'���M\bJ3�����������s轝�8���q;��!�_��4x��ca�E<P��ٷi=��0�l&�a�f�]T�7O�2w�[b�\6��3���L��NZ$���:ܻvT?�_��꓆�ɟ�����I¥�R!��1T�7�o�B7ѶϷGp���ROGO�=t��^�.|!;eY�U�p�kf��y��H�a��_�"S��}��_�`����� �Sj��Q�rfJש|�ڽe8k��� �|�;�a��l�����w��b������@o)��Y�=d+�v-aZ!�����vd}�	b�nrP��D��F~j�|G��P�TX�o��K�������&�@��sۘ2L6�P@��s�_6E�^�7SHk��$�KYIl�n����kf*Q6��	Vr���}��o�Ӆ������z6*>�a4�K�r��x�Fi4��u+Vf	�E���Ѱ`- ��m�1�w!������l�}7�b�����V�C���ޙPx������	e�|���L��5�5��i�d/�w�w�Z_�R@[�C����1�a��6~�}�
��6�ٳ�A�(�O7PV��Al�.����]n����v:u�7K�s�_ɯ�����˓� �H��R��V��S-*����N��}��M����m�q��d創Z%��A ���J��I�Z�k<�R������/��������_���T�Z�3��ؤ�<`RԺ 
b��ℙ����i�B$��2Rd���N�d?�~3���"�br"����%��k! vKIP�j{
=�
���8�f�7��wۙA���n�7��B�
z���:*�������7�i��c@�k^:��h��8�u�J������ &��*m�� ��󆬳�b�'�`��۷;���S/z�mzR��ɨS}��@6����0���J�6�	���ĪްRJ�'s��k��v��?T�#��z��[?HVS0��X�]C�VG�7$Ԃ������*S
���e�6��ӑu�
-C�,;����f1�qt~��msn��Eb��zX7��
9ҕ�N}>]	��P���Vd2���a'�"q" &��z竒8��M,i�<?|��ek�v�@���
$��4t����+B+�N��Y��>n}��g ����z"ԙo�#獘��ab�o��]r�G|	��M�w�EJ��}��7_�4�B��^t]��G��G=��&rW�jj����n2nkӞe���x�?���]Nh�U��6K�M�f��(NC��0R7o�1������pOg�Q�#LyA!A�U��C�9�^�Ǣ���f_���D�OO������宀XS@&�A����սִe$u�W ��o�ee=_�I�;�'��Х!�bA�,�9j�i��f�=2H�_�X��pCTױ��Q5[nC�L��6�5U ��e.��hi*G�FEI�� �72�/4�LGx�E�_�b�����X��MO��x'�Oh�Q������w�>��N�ok�9̔�@,V��9���ʭT}-jmheY������I�iQKk��2�S1�X��s��p��>�Ћ\��Rv�m��BFs}�e������	�JL������D8��/�Y��31ɝ�~^bd*g���� Vy�>V,h���v5�iw�N�'ϊ1b��q�5���T�c�C��U�B�3<6�Y.����a F�2��ip���J.��F�nz
ĊW��m����y���U�D�]������>yi;�#�]�êK>󂘀>g�_��["}2��\@� ���G=%H�"��
�q��_����ɜ	��o�(��Dp7c?��!�4C�]��I;^�K-��g�Tg� 6�h�۹��7$Fj�@iVy�pw��#ԏ#_:��F�pܓ~�{�f��nox:�}M�Pu��O�X�k1Į�6�-b�BmB/2�=j�F��,��?�XDx���p��W��b�%k���#��4v����o},���M��b�٭/h��l�v�S@/�G�TC��d}�`��S
U��9h�l����Q��=h�č�d2�=��ꂳK���3����?���!w��gx<|�z>%����\�S,C:yj�=Z�!$y>��o��b�HfxI�����査��d�,��Xl������6�:��lq�ڈ� &�����Sʮ�F�]���=*a4�U(�`�Q�xΌ(�I�@R@�$���Kg���cғ�`yl�h���"��j��m�486a����=@�	fyeG�0���[�Z�*�b���|*�(��j��M��ޢ�1��<�\8d�HsJ!���x ���a�6���\������=���K�8h���w<�� `{ee��-#�d��l�MV�:eoJYe���-{{�c��2����v��������<:I΁b�VZ�E�'g�D��EC: Ǝؓ/"W�Jd��JNg�a�bxM�'m���j�ʺ��atQ fK�g�ݐ}؅�(:�I� =�j��R\�ס�*\~��w^R�Q��*u���ºe��N���3�<��?���Z��H8���JR��Ĩ�O0�G�<Fr4�-�-16&!�Ԃ�k�g�����GAL�F.(P�NR_6W$"�>l�bn��ژ�:j�V+Ҵ=��1�S�X,���!B�S&>�U���� bYn�${>�E̫�[W��X�����-�k���|v_�C@l�V+�27ԝ+���y\��_:`����3��Tn��\�_���U�$�'s%e�Nc���Å���2{�?�R&�uRW���W��~����˂����fJ@��>Lq$��@���K�F-i:� �z+d% Y-���q�a[F2�,V[L�U���7���y�H���A�@9o�)S�P2�%m���OC~GR'�͹4��%E^\�`1-ѷ��/lؤ�>��:���{S�ǃ�"$-��a��2ِ�jL���.!&�@R��k�A/�E� 1W�؋��*�6R�a�m��y��'���|'|�ù�Z�b$.h���&ؤ�CԸBcx>7�Q{��5��JA9
���,��6S�=�q8��sA��1{S8u�e	b�,���m��/]:���2Y��+x�A�~���5Cn��J59kA���W�P9�S�v[@�vށX�O]��6�KcHk[S�rruP�iF�jג�7I�}���L�u�Tb���8�Ư��TpHi5�A��s�ui�t�j�������(f�'LT:{��F�����^���*À;	��(oe�]��j�:
���q֥Wo��g3�>����͡S��)������]�'��k�/�`����9<2G��l��J��]<D#�1s�C�;�P�Ki������ �|L/��G�[05Đ��8=��8�Z7H�=<Ã&����Ԫ�eA�3w�u&H����`�;5��k ��蔎&Ӕ��23�A���@-bJHK��,r��h��ʯ��q�����!{k��km��GԘM��X#9;>��5�3��v7�_KĞ���C<��n�U���ǧy�Xhu"uS�`B�|���P�w�=;Kg`��� (���Y�]N��51�k�,C"���0u���\]➃��§��y�M��K�X�A����+[��J������(mK�Î�F�p�nV�x�������&����q�v�z�^1h�$�nb���(�����{ ���w%&����m����m~+[���'f7l[�J��(mђb�K�y��j2%ބ�F�Ə
jR@����^���VV_�����\�b �c~CU`�v���3ݩ�MJ��������������=��f��ܛ"Rko��?�}ɉ;I����W�3�a�&�������՗��b���1�O�}�-/�U���-㿘6ᑦפU��2L#�>��j������IS
���F��n�Oh��g�cY��n���$I��l-��o_�4�d۵�`9|�f���B�����_������x�o�y�g���s���.K���-��x�߶�]��驙�{J��!�lT ��C���x��pj�`����b�lX���;n�d�̎f"�F�Z�0���&�j�%��"UU.�s�3Z���i�k]��P��#�c�)�t��M �)�[x~�0_(~R"�1�"��-Ó�G����tX	»<�.��B��7�]��)\UB���?p8�+�~E5�m����u2�d"%ݲ8�<2���5���9˰v ��c��Ѳ���4	��I�L���2�O�!˒t>�.���F�������<��,�_K��%E���
}�����VXP���2��=[�TYm
�N���rKfGs�3�dZ���+�xa{Y�*4~1���Z�іlUG�L��$�~{o*��������ڻ�Z�ۛ9�Q�E�tEXc߾�1���8,�����B���m��؇��/��Dl�W�����`�9�n{o7��I�8�x�]�[�J'��ǟ��4꒶�D����=�l5���<d���ܪ �v8i ;ps��n.co_��8�V�G��ݬr��_O烺T�yM��y .ֆ���I��`g�2>�z_!UN���î�' KF��/"��;���~[K�G���_��'2�@4�.<��AQ�	�g�_�K����fiD�����!����ލ@�PG|U 6�Abf��өh1��;I���CZ��Q�[7��p���<�ﬖ��ЅӸ~�u}�3��� ����o����b��1}�z�h>d�2���$\���=��{���cD_�4;S+Lj��t�P�����]�Y�Ï/��ٌ���0�G�6��Ո���b�}�F�����}�eB�k�����|��4B�����n\�n�IL\��ɥs�5jrw0NQ0��]�L����<L �3k��7�|�uW��iF|���	�W3�N�m�s�{C��Z�ᡇѯ4��t�,D4(A�[��Ƕ����_O�U ����$p�A�g��ub���.h���ҽ��MX:��Xt��p���-u<�w��'��WHlw����x��۵�Ȥb���-�t�Vi��dHNEc�I�n�����1HL���L:�!ط��Н��}�y="����	�A��o��G&���ed�{�_Q��B~[����9rXIK!3�E�86�;�p����⛦L:d��Y��^E�v�!R������wf��A,0�
�aM}�gXœ���眶�߬��x�4�U4��~�ߟ�W�.��Ķ���Rd�S\o&�a+��]tll�\z*�Mb�EP<Z� �EԹ������|��*w{����ʭ�9�9��)-��2ϔ��Y��^�%�#e��^{���!X�%}#H5@�[3�����FJ���R����:|>�4L�V��b��^�F�y�MR%�1b����N�e� &���k�l�б|��`����?Y��A����`B��}:���)��?qo��h���� 13wL��+�3�B��f\1wSf'8�T�����v�﫵)$�#�,xKP��A�~�LK�b(�#o�R���6�įO�p�~�
Ƌx��2�[��٤�ļvZ���z������I忘���0��ýR�<<1�]��U��0�˻W*o�
�)���(	VK��bZ�bChZ�pLw~���C��rr���}���<(>�t*1#�t�Uc^)+ �y��^kbc�X�q����\�u쁜Ueng�����aT��4��j:-��D �erB^ �q��h���v����~��'4�!_l��q�����T�z�dR�Q1B����@�*��r_�ބ�r����T���}{P�B����R�᚟�J���[_��R8�g���jN���:�bap�sx����sj}	�aL�Kb��~��%����~��b>#�%�A��&�O�~$�a[9�$��	�����!��W�b`%ʮ����@Lc��,���<* /Zw�3�΀
b.��dˊF�3��I^�|�0����Ya�\hM�Xz m̐��(���ƭDmn`�8z�Bg�l�hQ�Ex?�|Ż9d;�D�.����R�Q���:/�c]��Hc��=�(y���*��3�XwE~������_$&=�A��bV//�{�Z�}�"�2�61��<����>��f���� F�G�����M��kO��Uu�)!�t�+�㹀BfIR������.����SǏ�kI�U12�P�f����)�ZO��m^��]e��ʄ�z�)�bf�cq�;m���]>2����� ��Iy��fhe�� �cS�<MeF>`ˇ�e&W��Θb0$�����7��^o]Be}����}�@L�hǾ
��P��L�TL���R�l^�[�x�2ɢ�"�ܾɮ?��b/<S���j�	�5���?ƽ�b��p�MH��
����ov���u�ڍ4M��hK�#a�4�DP�x���Kb�-��䮈��3 �7RI�6��l�4�BE��v}�@LZ��CR�>Ů���rs
�2�{��O�\�����L��zC�@L3[� o!��<�~{pu�Lk�-.���}�E��w�)��wÔ � �<;�e�F���}��:h�̝� �2��s	gVj�W�f�x!D����$�
TtDa(jn*��]kb�̓�I�5|4׎�:Q(b�,A�xӖ�&�y���dZTq V�2����
�/���q/��jr�־N�rO���I�m�u��%Sx�m���z�M�Ε��T����m�V���I�@)@��GT-*�RI�b]�gTcI:-Ė΋y�m��|'L���uQ
@N�oO�͕N��Π��AaSN���Zra��2�y�R�CH�EA����HW��3���"	�
�p_1�ħ���G��g��|2 ��f%��pr|�Z�lC�z�E>�X|����x�&ý{�O�r0��a va�+B|X�]�rC;à����"�*�q٢�[G�/8U,�F����A���h�}o�K��@ѻP��X���%�3����u�D����WJ&��b�h��u�y���i�kV�����=T� ��7�BT����ˮ
��&��9A�B�`��'����c~�L�]n�5���Q��X�����	b�|����;�r5]&'F~H� V|!�`N@�E���ٻ_C(�	bt>�I��'p�e�����B����Ĉ$O��+n8�?��=X�BX�v�������W6�� ��~���\Z1�%`��!��1���Jzh���nIô���+t:�@z���r<R���,z�/6��A1��-�)�ԟ-���z��5������1ڎ=���FS"�+U�?yR���,�>�5�E	U*�/�j�0%�����=M� ]���xƉ`�?�U����-�?��5�v&|�e�������O����[D-�����)w�Ӑ��C��h߇���k�H�o_jp��n�������4�,U���?�Z!�P�?OֹKSw��FQ������� �r��QT�Yr��V�Hۗ��@�w1�P���wd���<?���c��U^��5�l� ʹ[�J�|��ˠ�P�S��Ƈ"�nE�.�59�]�w/��~�qϹ�o�7N���&��K���/V�5�'�K�F�/��+����G_f��v;���U�!�k����_.j�'��3�X#�o>hh��p�1D2�����.�8f����g1�ؤ�V�����
�v��M-�
�k+���3F�k������t�[4X]務�����֡�S���U2��Im�_�.�
ӄ�k�
�1�oor����~xn]%�y��.V|�5>��������\/�F�w�����!q&oM�����hs1S�BR�8�o���ds�\�`{�K�Ý��Qk~�_��\�:Z�;�{������XkA���fs�{�	~A���Ey��� �a¯ϣ)����&�:D���17�8����ա1��A�{�Δ���Fie�YO��|��Howg��x�~�7&�5�|	��;fs���f^�"�q�8��2A�Z�R���J'��additionalMissiles
game
hero
perml00
perml01
W?MzUx�G�I�@����Ka``�����ݧ����Y�x���\���)l���{�8�)e<�v��1�{��V߬��K2��m�9�z��E�|g�(�����b��*�冕�
'}��nD\�_����j�E���"Z���}�B+���<��+��)�� =�<���ܫ����Ȧ�xHET   -   ��<�'�g0��`M<��|`��8a�h�y�^j:;�K��dL����0�����8�?�H���BET   �   =gH=0�� �5���5h���2R�6xexd6�oG�����3�\��)+W�U����<̚W������J��W-W�F��[���ZvBVt���U�aq�m\�E_��lS }P���Z�4�Ѐ1n�𯺾��c��	�����N�=/���#���U_Fݷ��Q���ձ��_E��U��µ&) :���H,�O8��:̓Ė`dEn|�-�d�M�O�;@7������#�j� �ѿ�Jl:��gH_Dނ3�Q��?�`�l�Q�ͣ�<����(�ry�ysy!͹�FaQ�6Kݵ�R�H�R3-�[gH=`����5�g6�X��7G$����#,IW�6כ�{�����A�a��d!}�&9��6۷�Q��L� �8�(u�!�_�i\���B��ۂ	�7�\�����\a"ڃ�Ƣb�