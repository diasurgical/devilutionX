MPQ�   ��   �� s�                   ��     !�     ��     �       p               9       �        @  <�^A���"y9c梽A/��)�z�:b=����Dss                �UL� �h�-���Q�0�����8�?�H��ވ�*Em��11:P�u&�   1   �{���Xq����ʫ
���.O�X�.CW �< ����V�R����2�@     �?  fh  d�  ��  ��  ��  ��  �  �3 �N �j ׃ � h���w8��� `{�-{���J�����;�l"��"�RY�3�R�^���~�Q�I�����}ݕք��&��o�ky0b���{�ĢbC�Ә��Na� [fq�j����ŋD�Hh赉Ra
x�x��^���Ǽ-/�)�٥�q3u��֊�8#��H�
s�қj��TR���y�����5��fߦA�-��Y5��+���6�C��k=�}���p��Lv� ��[�X���(�[3�Ch��L3���G��d�]��jl`OL�/^yo����y{~���{�p�S`W����	X[T��Z[�ȭ0��x����M �V
���C�;4K`��f�͗89]*צ����!P��2.�;0ř��n`��^�*H���Vba��y�v�q�5h�Гߡ�����L_�S>��D�Y�5��&�^c�W/ڟX,h��W�`������d$��n��
�0�h���[��j���S�6��	`��b�-����7k��L��oߋǚQ䕪.sV�!*^�p/^nS-І�?�[/4oG-���t
S����1����'�8�#G��#04��6�7}:Ns�>�Rw�:��e��?l��=(�!���rz��?f��O��
�!zH�c��m�LSZ픺��<�����8���_2_uf��	E�fLP[j��?����?A� d�03�w�}�O~�H���0�G��Ԣ�w{dnB�����U�|�v(.�|��R#X��YUYm���������:�l���d<h݂G�,�YC�#3lH�|ܡ�b6a[B��W'n*{F.1���o�A1�A�e����qBԩ��؞��bu/��nS�����q}I[�2�1m]����R�FEU��u��k�uk0��d5Zh&��PU�� dז��)`��ԎcUd32���O��b�5n���f(�.`Q5G�ʹ۠le�9/�]�2�b���#���w�V�s���vǑkA1���O���O���0�\�����j!xC�,&E�M�.9�W7\�P��� v�~<3`w��2��g�N<,��=��k�ӏ#g�A�̀w،+��e��&Ъ�zB1��S��*%����I����P��jS=����+��KŘw�+��A ��K3��]�TLFhh�~�_/����%wڗV��oH'z��	���0'`��쏇�-Ğ cl%N�W��u�_Kǝ�U^����6�U�ɨb�B1��g��ܚ;�����W��>�b��;H��-�B���� �/�z4�P�40(4Rp�L��� �������p���O�bcs�],V�UA���m�ӧk�!b'`�U�{��I�=`��~�s�D�"I��&��)7[�B7���M��c�%����A�o��)��d/a�W���[UeO�y����m`�r�a {��nE?;�UQA�tL;�r��\������ȶd'q�����%��l��4�;�ڹI����N�b?ШV�{@k����k�O�3;�~�	0G�RG�N��5�B,��D
�F�����KӖ�M��Î>1�)Ώ�w:ɼ{^�w03����"_��ѧ�zK.�a2��%�D&|D׳'����)AX0
�G�6�Ȑ^�04��-5��c l�Ň�9`�����=���OJs�zw�f~.�?,�+�W�[�\�S�F��ጪ�Õ^ٷ�5{�R��>�6?y�P���yh�I������Q��>�����sk>gO�;����z���u���"���
�d���#j��i�&�4��xh�ޞي���J'CwILe���Sg�]�CKc�&l�:4�� �!�rG������6j��E��Þ�1�ގJ��1栮g��g�D��:J�gL�A]:x�g5���{ލCC/�{�F�,h%�$^�,���kMp���v�`�����*͹���O�i��~p[��i�Ś��Z��Jg��*�P[����f��Wq��Ʉ�Z�7U���mF�*�����;_8�U�8�_)�.N���71.�n�6^�bw���\�6xM-n���j�&y* gr��]�p6a��� ��# �2o�=r�I�͞���G�����:MX!0���"�����^S�s�@`[3\����٪L��Js��[��jOMȧ:�W׾�� �\�JY!��.J��|�ٜ(�YM10'`ο,�Ek1�7'9ݣ�@�#K�4�� {��Y�[Nԇd��kƮ��:�
�1�o���TY�@ex�x�:[�T�8�
��C���l��4��_�ͯc!�հ�Ķ�pʥ�f1���r&��+��S.�ҶxW;$�x6�F\S�>��W��5 9������j%d^�j9���N���4\�m��4�>���u�R�I9Y&b������6���2�V`r���*`'c����R>����5�}#i�
�4���� �v�ez����b���D���~A��=���<��{}�]����n;����ҩ07�y���~hӓ�.�IL��D�"�?�V�ۡ��J�f�#�ۨ��Aa���fNE���'h�J�#�m��Q��	UT�-���q`V�to����?x�^;יnvNScc,-�9�T���_6�������X'F�L��i�l�//�3H^K:�Ůq���hJL�.5���S��D>4φ�-��?�;�a%���V�0J�,��)���gӼYѡ-"aSq���8�Y`�Z~��u��81��/G��e|�8t��~�q�#��K(=^�Ë2k����]BF����1k�i��x��<V\���rM�����~�"��� �uh����XD�:��W�wBWY�zܣ����H̡X���}n|��D�ÛlW4��(&�-`-p�� u9����4�x�s�%՜�`�D���k���Lع#�5��=bjytvA�n޸�a����0�_�Lha�P�+���:�Ŕ�Ok����qv�f.��:GH�
���e���p%4%#���7��;�� Gf�W��e�O�*��O��h��2�K������uBn�|�3�QN���b�60���{�S��6��k���w/��K�C1�s�βκ�}ϼ��8�uI�֠����b����\6'gj�+�e(��2�6l�5����z����FO�?�;���b�,���f�$Fk�-�=b`����G��cfl��1��$�9�<�D0��k���㎠5x.�:�9;NN��]A˄bb�s�X��˜�V~EO�D�_�bF��l��G;D�J䓫	��Xʽ�(L�C�CB-hS���-��o���k&3h�����zx����v����9��g<<��rX�&_NHҾ��R�&�ѵpx�Z�x����6��ٗ�XQh���Ț����;^m��y(6I8���vf;���tr3e�2��i�aWg��G�M\��V����/��h>��疃��*�/^��.��4se���R�n��g������f��uW���"�ٶ7R+�<�V ���r�'c�F.�<_�P���b����z3�=DYҲ�:PL0�,��l��;l�ŝ��Ǵ�`����L��|�@3���%�������!z��'#��˳b�ٱ	�e�����?����*��+p72��p��fm��[x�}#cY�O.��!n� ��ɦܠ5��HJ�6��ŵn��b��bOˋ�rxlK��t"Y��z��]HW�4�^���24��ur0���MJ%�Q���Uk�e�׻b�.=6o�^Pq�R6�~�����\sSV���Ř|�k��	�ֵ��"mK�u�qER�ҡ�k�f�H~#�7��9��4X+TϠX�l�+y�؝��A�������I�f�����n�J����>X�<{���#��ݠCC",�p�
�>�������M��/�G1��Qu�A�3{���/�g���Rb�p9��l��;D��+EmQ&�Х��P�ih�5`K��A|��f�%t;(v��)7��"�J/��/���I8�\Dl�44?�k��0=�[��~�^K����%��W`�G�o;��c��!aR�<i���iV6(ƕ�6�Ly���v�zV={	���b�6�#`GO�oEUw�&�]
Ŵ�%(��6�ֲ�2;S�����%c��O��}�Ը~W�^v�r��%�o� zh�[e��$Uw��$ĥ_Rj{��q���p����v�� gn..ꫝ�PL�M|2��'4�vZ� ��ʁ,��Q���ݴ�B�u%Y&a��<�פ+*Iz�UZ��DoV6,������+�.�#�cbTR~�`�@]�X�F��}�~<`o���2����3�25�}��pX���H���"��0�"��'oc�';��蠘N�C��4����l�.�V�w^Q|�b�N
JX�U�Χ�TmyHbP8��b�\�_҅��z���ӎb��Z[�����/?#����s�嚕�����殘C��yd	,�?���,��3o�����ґ���VՁbI��K�.�>/m�(��O�b��xO��H>��+rV9q�1-wr �-�.�%��R��me�J����Z�6�w5Ec{P[�����V�	�kk�4u�:�W�>����c�X(�ׁ9��`(G�oS����jT��O��l|�d�J�X.?h��ǩ�߁پ���B�ۆbq���&��7�I�hb���^��b��v�E%k#��90����(�� �2�
�eG𱖬=<�L �@`������;{���\B��;	)����G��p+I��b_XNO�`sn��E�2,&��ν0��(�0T�p���Y�aSA�V��v)�G�}��$-��D(��{�Yq�SD���ċ�2q5ͩؽ�ޒ}�.�
�ך)���'t)ϰ;@�'<j?0Y`8�l ��s��QGcz������ (fs�����Pi��My��g�>;@�jr��ZA3s*%����AK(6�g���)x�ggfD��<����Sf��IȜ�Z�(u*|_���zػC�S���z������۩[�O�y��yuh1O�'��ˁ�?g��Y�L�Z�����H-8���+?1,�2b�K7�	��a�{�ٵDH&$[JN��o$َ�b�V0�#�\��`���7�1PL��Jc����/�L��L��8��FlᔖH?��k�;75�B��������r�|������,j�·�/
[l��GP��VB�����Z�j��-,/CfUr�ҡS�n�V��J?[9���l�SqP��)�(�<S#�H}���x�4MV`�F��	!%�Ww���F�"0[��%D�}�K,�m�:�q��Mï���x��]Fv������{ѯ�%|�R��a=�r��j�
�m��8[a�<���B�{�Dϖ�F[�BM��,
�$r-Kt�ʱO��-�w��ᥐ0�Ô#x��;�G6���ub��������w���x�M�����Σ�Z��S�XN[W�]�?Z9[f�w@��SQ�t� (&MUwes���8}�6�}E1�{^%�TC��-%g�L}�;5]�S/{�K�Ɨ��0R�'!�2��?t���$X����u��7CT�$����	:9j�I��eQ�LX���dU�r�G��UZT�HYKb�b����[s�/j^HWJה��-އb��̈��f>cbW51KpR
��b.��$x��l����H��@1��M:!���8!� �>r�}�68�x���>!?�i$2a���ۍ�g:�U*lx��K��u`3G�o{o���I�0&�YQ1��\�!(6B�V�ͥ�(M�W��RϠ����=��m�\M�ի:�uK���*hl�	����B��$��f}L��6f���<3-���sAgb�ңy���1eD"z���k<5���Ӓ�Ό��,�8���)�3�<���~���EEa�6(�e���;����*�s�-[�������Λ��y{Q��|D���>+Ƣ��}�R���O'��7E�H��?,@
��ؕ�H�	�*��+�N�>��1��Q��f�)��eYUh�3�	W�O���Pay��{@��"w�Ҏ�>6|�9�lw��.(�Vs����r��k�5q�|�uPLm\�۩V����g��܃dRˠ�5Z�Ɂ�Oc�|�ֻo��'Se��������s�3I*{z�X.�{^%�C��ܤ�,X���ގ졙���J'ɋ�咬vS�A��ը���]Ѽ@�a�m[(��q����F�ݭ���!-K](V��d�+lE����rF���ϒvPlth}�T��7n��h�tѬ	�<��6#65��������9W�D�+�K�:��s>_fg�D���tM`l��*������=(��M�	�L�'�PMy�ڜ= meV��߈͈t9�L\B�9hOױ�\e���r�z�}�D[��M��P�cZr(��4�R�g����(�PVґ�h!�'Vl��^_�O�gS�n]g��n%�R�h����P�,�֌]k0YQgL/�}�w��b�҅N#���&��ԗ����sC�wQ�ۏ$aON��>�_����ҽ���?�����(�SU�m�����ĸ\w�l�����K�$H�^�E�;j?�M`>�PY�,�}UA)Ef��g���m���C1�9�+�/�/�Hf�e���
�C�w��C��ň�:s�����t�	�5���Q.����xS�O8��AŊ뿷h��G��hTR���·�'�C����ä���#ŰO}���=phL�[�)�����?^�
��ǯ�hm�-���l�I��2���Y��#���Oj�6���C��;��F�E����^��z��Y�}�碊U�S8����*��j8��b�/R�mz�j��|�\��E�,���D�����E]�v���l�Ѹqrz__X=���8�~�cd�'f"S�P��IiU��[����JW��+u]i�����4(�w9y�3�l����d��]��P�� �̓$�v˫|��ޣ;���cZ�(0m��S>L�!���M�"n�K#�J��o�ޗ��Uk�9i�1���a�*$_���L�8�������J$G'%n��}uFX��Be<h���Np53����YP�� nU�-h���w<֋���dJ�� �%Y��ٔ�U�J�.##{o2B6�GFȎ�.�R2��o������}��������1�-�����%]·�JJ�+ַn܁9�%�"�`h�Nlb�"I 0���z����H[��K���ճR�;�(�d��t⤶�S�������C������?�4i�fF����9�����L25��N��#��e'�"���݋��"[��W�ބ[���L�f��2O�ܙ1d�<`ZJ�){'�W���3��J���٫���S�����S�>m`@U����}�問D(n�b��_��{�e���r����|��\UX��e�c�-��vƌR��>��������e;��'�9/6
�6դ���p����;��cT�'^ȑ�7g��9w�qۉ��+���_1��� ���L��� �[noɯ_l���|���BJ�|�2��C��`����wK��N&�r^���2jK=eV�J�]�3hv	��<x%�L?�X��w�;1�W�,ֲ|��5��%f�z|�S؉u�3��W���}��JF?������`�͒��LOUp|�z9_xԴmc\f�K�����Xf�>{o#�����C�<_Ll����W����U�3�g�>��{admO�+|L-mtZY��8�N�uC4�W���:�Y�إy�wbNir���K,M}�u=~��\�fٵM窢m��m��1�uW�A�yON����x�����n��ǘ�&�a]ش�%�?*=��7�vb-��]2q�����a/�=ط[oɿ|�cܯ��e/ݱ ���t;�J�'��<R������w(�����|�Q"�A"�Ĥ����t�$�������)g��E�+�,�߿oD,S�c����Ø�K��u�
��,�t!��~41g����l��BH�`Dz�nI�t���T�;�[O���۵^�~2^��|,e�0q;�n�{RZ>�|1���CO`ҽ�ٷ�|��f��ғ"f�ĸ��8�Y�~_�X"vw�gT��&�N� �i�����hb���*�-��Qԝ6�;�u6�V�A��`	|����_�ʛF�{�X�bʥ�8�#�><(���ҡ,,��3����h������%�
	鷉`QרBV�P���c>^�f�]��|��+�F�O9D�;IE(i� e=o�TU����xIV��?���n���&��-=5T}:��e/%Ln�Y��Vǁ��5%Q-\Ǚ؅<F_Bj���;��p{>�}8/
�O����~4�c��ݾ� pU��I���ע���G&=C��0�0&�x�PW}���`�`T`��=K9���;�����{��׷:�z�|J�ur>s!s*'S�j�Y�3��ja��ژ8:2�pz�w��������2�\�*��X\�9�ş�0�V���1%�m�a~m����n�w5�M�޴�`M�X;ʎ\#����5�y|��V�I}�C�N�����<㽻��s4�s�����m��	��kxGb�[$2��x~�|����$=���*�њײK��*b`�`�n�{�$v��ֆ'K��7�8�&�����i��grˮ�KrVa�Ƕ��c�����*<����i����ep68M�O�Γ7�e�����Э+/��mo��vq`��	��sN��R`�
�p����i���=&Ma� gN"xx���J����vb.\wbOk���\cӊ���O�&�*b1v��4��S�!�i{�-��4��ձo���͛�M�(|��k�s��%b�`�``���R&߆�Ig�B:��*��:��Sb���=yϿQ<j\��겝�i+q��~�NtU��&@��!�Jcg�Xʗ'/{���:����w�� ���D���і�Φ�~8apAqQ��7b`�����
5��׫�*�������?X�k�(/LԦ��k�w��{Iޖ���&���'�-t`e�Tꡳ��:�����TWR����Wki��;�}'����W8Ŧ�qGwb_�7��?�/��Z<|�\�l'�3�iy�>�l�A���]���8��N,�t�d�;"9����U�:�2+��ml����*G>� �Z���D�}�w�S,�f{D��W���<�����\e�ϊΐڢ�Z�&��k��N̠���L4:uU�|��$����;1������x|����o��-j؉1�ܭDMGT�R�>R����ҝX�aS�l��4ũ|wqh>ły;�۶�nG�I�6�{`z�����Ꮇ��`re�O����ȱ�_]�&m<~oS%��U�cU"��C>;�g�����<�v���f��GN{'�!���Ou���{��#��܆�e;�w���e)]�x��+��3a*ۉY�g8�Xpeǲ��~E�ה�����ڭ�(-�uYX"���>�:��5:�O���Htce�˜� �fFl�Woϛ�e�.���)��3o�<�5B�j�ng����	HU�l�6���$����J!���|����v����L��X�[a�d蔸x��������K!_����o��:O-S�أV\W�i���I������v�b)�zSMp[~�V�.�G�Sx#F��uK�1a���
���.���{�ܐ��_�V��'��诽~Vd�Q���3���{s#�o���%T��]M뽗uf�R����*���l�C���U[:���	�O8k%a)�ŵ���@K���э|�u��12.��?V�����3�e��?D{3��(����������x�i���P����-�&��7��"�����O�&���ح�?��1��}Aw���8vs�Q7�/�j'9��M���ǚx{�G��Q�r�}�xრ�y���B#�z������x`��f.�\Q#Ϛ��0���pi�l�JC,�a��پ3a�W)׶�p}�.K&΢c��T�}�x�]��ǐe�q2�S#���DϷ���!����
�u�H���%�z��1N�w�\Շ�);	��C	;h���J q\ٴ`��v�t(S.X/�4*>�D�|��'��.
*�K!O�o��i��N���!��Y��(YϨV��8+��S���٥�6�b���~g=�V���wtwzK��q�߷�0�|�`����,��/�t�� Sò�2t�����WZ�+��'I�IU�a�3�`�H��o�����]��,R����p�|��ǫS�;���K�F���>M�gs���w�y��VI�՛�070��7k�l���S�b�)f��ajA"0�=��,#��xBl\}�15��	��I�J�o'���W�յ�o�r�+֔��vbUmt<������$���.�Y�����i���E���o���g�s'�vb��»1���W)Z��3�tޑ��[�8Qv���c]~��g!��Y����� fo<Ťӗ�N,N+t�e]f�Uc#`�I�LL,L�"�"�2X(�۾;}�O������z_���)�8�;}�`.``�p�<�D�
�*���NUD��~�4��W���r�(�H5Q	X!�
�4X2X&��X)XBDs�j�q�Sץ�[��ĵi��E��p���D��������i��qCL�D.��r�����Q(�g��`�����������U���yߠ�.q��!�?� �5#�{��VW���� X2XX>�>�{�����a����;넫�-��^:�
� Vv,�l����%�ݷ������֩u_���v�F0=��`#`�`�����e����I��j��H��@���/��'Q�V��Y���	�[ �c���<"{�"5��|hv��A���#```�`����=��s=Bi�z̶�>@�<��H�[��q���� �&�M0s�K`�`j`����'�^�wD�ea����Y8�4X>X$X�<��I05�<0U��]l	:�}�r��þ�3拓�kc�`k�%n�Q�&I<��H$ϿD!g)DK!]sm�q�Mn�()��P&���wFBg��}�l�ɨ�������DY,چ�:��Q>�f���@Ya�F�ҕ'�����j�"PV��W�`Cuu(^ H9����~� /�{��\0B���c�]�̡�p�_�ώ2��~:bNF��������e�H��Z<�b��,?M��he��� ?�&���y���auw��҈�Q&��ǥK�`y7C���'��j���@�,c�nӤ���-�L�-Ү�z�+�U�;�ڪ�u�;�Ş@w>Y4���ȁ�{�s��������:�/�u�2�n�8{�dѳ+Fu�ǡK�ѫ�R|�Ƙ&����򞒊��`3{�Xvo�o���u�Wp_S��O�Zra��m1C��-ݫ�ݜ��o��;P!�w�F6s�	�d����,���+�=����q�����*���a����7�X�i0<�Z,�A��)~d������
�nvI�����;v��Gٗ��E2s
5b��e�\��_���9��),m�R�^��Ns��(���.�{E���u�Q\Uߟ�?����PF&t4B�ҨtѫÈ�C���R�W�<���������8�l�o���)�e�i������&�����IE�sr���:�]� #�؇�0<��O�9	�-�o,�gCR2&�vWxΏs��X6���f>��'C�1�z�9qa��OwEmY��H\�g�wഄহ`+b�[�ߘ�燆���'��.�U'1���"����&��1]ka���5[��u����{*�ޥ"Vƃ�"�F��X��k��0v8Ʋ�-�e@��c*��&[�N�Ox�{ 	1T�HeӲ�L�����7�r��f�cOj��f�G� �����ԥ<n�Q��Fd<�)�g����C�c��N������&m�Y�~Ig��v˗�z������f��_��#�-90��LL���0tv/�1]������ے�Zh��`d����X
�0!�ݘnhT{�H�J����
��(��{��0U0<0R�N�����e�$�U���2�"��?g�dT�'�ȩ�����-cu��f8��%�6��Tܷ��)�s`_���C{m�
�n�.ƃU=N�2�P�4�S�i~����zoc�y�v%Z������Q� sG�*ڨ������>1.<�k-0V+k�!�;�@��-�ǋ'�s����X֙�t���9c��o��f��=�1���t����3�BՃյ>^���F�]��O"��>Ʀ�������
�6ֱM��9���*��;9��z�0 i�_D[#bZ���[,��;d3W���Sgnv콗��D����j<�x�'Z{�&�Y����cL�z�����U�I���i�鍉�� k�q�>�S,@��	ll�.�0�$�]�2��Z���cX �}D�b��xڸ����bu`2c�/���x^�r$NС�0���&<.~�/�Pc��aw̷v�V<�"/a�lF�Aq\� ���h9OEX&Ǝ*�&�jL�=Ϥ��f��m�qJ��FI���q�<��1X�Q��N�hĈ����\��T���
6l���2��<�d��ۣ�V�j��^G��a��3����|`�D}�S/z׷R���k���}1�|�@�L˿�I�VW���� +�]I�B��a���*��D�:�V�V��vl-)�w_~;n�&�Ɯ9�
6	����a�c�9��m��|��P�i�_��R?w~W!i+�͂كՁ	�9�R#�c��u|4�`5��
]`�k��P�Q:D�i�Xv1T7��v���W%��:};/�ޢ|A�f�X 3�ށف=��t��ē����rzM��ON�	��#f�����f�yI,�tF8�Z8�+g�qM��&Ykt�wwi�V����޳����e���p��5IOKp�s|��m�U(~rU�'�3X0�(��b��b�_��͎���~�!˲+�����#�O������i�ql��h�3�V~7�������!��2��`3`#F��:�06��Ww_g�s�t�G�[�z-黤�Ї��Һ= f��,�/�1�Lg*՜t&,��[���#|G[S�FYж�v
��C�\u�Y3�B��3�x��M�n���;���j~�%ϳ�L,��2�Jz}�iW��j����K���|X�m���f���c�<�?�#�VV�ɞ�km^p��9W��1&a��`���l�Ï��`�`��8ëIϸ��~6���̖��]`�݉Bۡ�.=�_��,%�6A������nך�3�h߳(-"&��)�3-�Ƣb҉�)k΁)����N�|��!kWU�5�{�誵ς�������ަ;�2�W�n���\�_z'�)��Ӏi�Bb4*[�
:�"~N�T��+v��w�����N���ʦ�U]�+�K\:�@d]������GJ���Ov�s���)�%ҫ�+���c���!�v,	l�L�H�'���(2�GǼd��J3VK2C[�:��V��·��X� �����E�m����nh���2T��vR�d"����o�������w���'�zi�1�}t�×�6��"��.*�S"_��<x��Ux}�!�3�y0&0/0� �HO��:��2KCX���C1�J�g��ۏ�|S�5�I�Ţ���,le�/�>SL��r��~&|�E~��q�r���^��������Fm�e)�J��1�ڊ6�]���}����.�[00�]���K���Z���MG��7`�`�`�ߡ��>�����V��x�b��e�|�"�w�X&	����� ��ӆ��:F�g�d9!��}���+2DT�ן��4_,{���� � �x�]'�c��v��O�Y����`��^"V6��{���a��KsT�,3��qWO�-j�ˉ� ƌ��a0�q,��9���f�^��,u{:�����A�CR?W�m�m�ϝ����N������2A�gt��]�ֺd��(1]�����`a`�`8`~`�X�<bD�`�����i��(��fq�'������-$e��bB�h [_������8A����}��.:0k�X�����c̆A��a��?�\�R�E+�J��Ƿ����*���#�&�
��
�ƈ�p
*�؄Ɛ���MZ�S.�VmO�|���ֱ:o0�r�_(ˎ�s>-7�e(UT.Ż��Z�5��6�-au�$��'�x7����%�4���<�d�B��^�����	
�4<,BL�F5�M������lA�������`v``���tE��0�U�9<�����7���O��tn��2�5�����XBן����f%�z<��p7s���|Y�����x�1��u`u$Y\`�i�(��!�"GN��6�H�>m�&�#09060F0&��m�J�y���;�"�*��������F]�6%�50o���[���mM�e7�F���-G*�U��^a�0��3��d$�9��ĉ�ۃ�+~CW[�k�&�n��va��(�!�"�r[B,C� ��	�lL�|$�sYN��y���"����
�z$�	 ������Ԗ�~R���]6��ׂ5ή�>'���.K��k��߆�2�ުη��O����l��үl�Ύ�}���1[j�������E,�G��Gç9k6�\�>ˮ�`j�S`�`N`�`�`�`K�Q�����<s�B��k��*�K7��#,r�x�-���j-b`j�_����YC�������.����a�g-�����0�����Gm�q��$�R���,���:&;{(����`z`�`�`V`�[��a�n�Yӿ�*,0�>�,mBK�VF~m$``�%H�M�筫E�J{�v�������z��m``>�q��d��76b챬N�}��ˆ�����T�Iח���%b�b����l#���A�䖽��&���������D�fmZ``B`j�N�����Ϧ"��}�s[!�*�/�4�s�j,�tEo�~��xI�����L%S�����������e"��X9t>���P�`��1."�]1B��|<'�	`;�>�� 6�յ V~l�c�����C�4)��F�L����f���%����������8��h|��t�`j=Q��R:͍A�D���o�f��x"1v�"�O_t�w\$�D�U��Z$��*2K��`���Q���]���t���"�*��b&x�w�%���D��
���"V�2�t7e�����hkX\]ҡt;Y�y���%�-�,���fu|���96͞A\��b���WB�	�v��"Ѫx�^�i�Xր��#�A�/��y���ά���9�q�6�[`r`d�}�E�50"�i�7��_�F_M�#��QK9�v�=�F��\���|������E��Cf��������4!f���l�C9g��'k�:�<w�s'�Q�J���Q왇e×����(8�U�q�� {��MW�2����"��,#��ɻ�VV���(�4�ו��bO�{e�E�ѷ�+)�u�o&-B�|�/�ɀ�����-��ھ�c\o�-����� �M`��E���tۭs�Ou�ʰ��W`9`�`�`�`�`Oݢ>]�8Oƶ]%x��{�9W�1Z~��5�I�qcu(�8_�'+���9��TR�Ӫ���\A�����b�{6�.���4W�W]d��4���~S��Ee������0�빮�iXօ���wOn�{$&�jc��������*��Ղ����"6[���`q�m��?�}`H�[�Y��$�?V�e�Yt���C�>X�LTG��t\!ҡ��������p�6#��c�����*���Em-�k�Tt�p�]
|�I���r�U���傕�q�} 3��]�~��,�ȕd��ϑ�AE������I��'����KɄn�殤:��Xͱ	q�_�b�<Xv��ؒn�?U�G��yT_�0��q''�^���V<���9�y�R�M;�e*����`.`4`��D����Ȋv�{��`6���;�;ڔ������a� ���/1�g%/����E�b��hS�+Ų?�{/ռ��x�.GN���"�3�|��z3<a����ˀ�ND���c�E�w(�D*�t�ٛ��{F
G�΂%�%���cuE�����hh�m�w<��ۀq3ed�"���Ѱ�
�({��iX�B(������,�3CFvFV��J%�y�����y����0��JR>����4�o1R������X3X�M���.�n�5:0:S���ܧȲٯݲ��n�r�� ���z��7Ξ��$���n��S�U�x{�1�ݙ۷�
��3�K;�v���H#ٺ��~&oU���������X��v�`WWzG�I>�
=��TJ��8%W�����4N&t�e�:�����Lww�S�\�/�E��;����������y�	U�n�ۡ�1L�ϻ�2co�`om��wn�.皂s��`��㈕*`�� �X����9|��ϲ���Kh�V�vp�e���
v�e9���t
��	��ό�~�u�)b|oO��ԟ8��uQ� �i�	��*k�~�h�����x_���{��cSk���nc�5�N,�7|��=���Hyw����=�ɁQ���9�a��T�3b,�-q�W�`�7�" �'��,XX#�X
��R;c5��M�Px���b����ՌW�o%�9�n=�%��~�΂遥��1�р��l$�#a�j;J�ڴ��Ь{X1q/����v�a��Pͪ�v�\i3�d��~����TXss�G�S���UV5��Kс�������󽧉ZOu�,��X��B�lw�."�y���Gq<�G^�ɯ���~�H[�&�6�X�7������_Tj��:����"���`��*�;�_�Xk � [�Xy�������є���%�����ޛJ4�Sp֝�3�X���	�:U�{����:��M����՘�����$�4�����E���Z�h��jlZ[���s;��U��
�O�`�'������el-��s��g���&�q��(�U�GY%�I0�F���=��q8���r�wD�\�N�?��ؖc�g���{x�w�	e��} [{&6�C_�E�#o���k@�Z$�������ՂՃ�㺅,A��)N�e�itt��GLi�4�t���ߎ{��66�3�D�#�co�;飥ܡώ��"(Q�LF�t/�jw,e�ǣ��[,�J�o����'(�zfv�-�k�4T��P�X�#�m%��+���YTU��
V�XRbQA�.����"X��#"�m�dD�����Z�(NI� s��k��>�1��ێ�P���o�|�<{1��ѱ��2�O�\�:
ƅ�,�X	!�5��9�A���w�H�H���Mi�+��X� {��0fM��������"�.��%f�ݙ~����d`�`�(�Eu����6���W_���_G����_�ʪ�=���8�`�FPր�# �h[��B{�˥�sQ�疥����*��K��Z%�0Q��{����G�®���éy~����5�#���Y���`+v}�ǃ$�[��W��4�/J!F�k�u{m�e���U
�����w����<�Ae��?޽�3�&�j��{	�F�+���>f���8hb\�#���;`��X3k+�1`M�˜��T#e{vMa�c�c��DFY̶�X?)X��D�Ї�=�j��p�;�.#7�t����3�[/���
�H/y)u#We����k�F	�Ox9�4�+g�|I~:�6C�%�J�撰& &V���~V��&J�P�@��T���Jw0^�l����$�o�5t��wd±X���G�:�ꏙ���S�l+���8��/=1��
L��eӈ��D5�%+�����`��X;�>�F�F�� F���1�-��q����O�n=�nO�d���,��r�)�`M�l�l�erT�v��Fff�@I��}�w�6_����Y�g���[�}����:\��B*gC��֝f�����5LL��W0Z0�ݝؼ�b�R��آ��4.3�f�sk{��T�[�[Ԁ6ơS���/�&^����2(��B��Jf��D��C7�¢~=����eT<ug�Rƅ�3_h�Y9��`j��AڛS{���Qv1L�,�L�3��� I��9�@*�@��w`T`5�%_�-X5�7��K��Ν�l��}w^aj�gb��X{6������/�44��FE�Ww��fF�\��de���h�1��X4�f�?���|���_!�N�kʦh�;X�X2X�cC,����hY��������nE��煀I�] ;�t�V�.�E�5
�򮋏6>�g[��PPu(2���� �b`7m���y����1}c��ǿƶǭ��	2�+��<�������Ll#Xbn`�`�`�`V`��
q]�令���Fw��%�g��Mc��	,,uW���e�c������	�~t�ʿ�m�����6�����u�opy+Ӿ�z�~#�/_f8���U��{S�_�vx�Qv1L�6�7-�(��v�L�׹j��/�i����������3�X?�ؓj"�����I����&w	�)�2�~�9fm�8���`?�_+4U�9��/�?�W�f���X�6��W���_�N$���$q6�x�#�1I�I�v�3��$�L��J�����
��,�?����<��ڳ��)���q����Bh)G�����2�UG��[�g�;x�(#<|p��9{�����^ف��#�E�֞�Yc˪��1�����y�e�HcVI.���$8VMܰ�^�L�0DY>bF`�``q`	`7��?���x J�O�ۙ)-oޙ�� 1NE�-"��邅~|����~EQ�s��+ggAI�\+�:4;G�]9;����.�u���X��tC�c�}]�����<����HB�O2�|�t��GʲK�)x�V�PE3����ͺ�P*n�n0?�J��`D`Q�=/������X���G|-.z!�z1L_kl���p�m���am.Nd�/T_�����Df7	٪x�F=oOf�
�S.0�����i1�3�Y�܇�t��y0�4���k�8=ۉn�CL����$����3�	&���h�>��FJ��t��=�0;!��*֎�q����6Y��`�����*��|¤�d�imW�E�e0020^���K�o��l����}^��k�6F%dV�z�}�*�+ނ;f������I�Ł���G6n;�+R2T�:��3�
r̀I��AL�k�`��,��p�P�-7�+W9߭�c��=l{Ǉ��`s`V(���ֿx��.v0�5��L��=�q}���-�٢�ӇN���C�^�ϏO��a3v�g�J�)5{���,��!��W)=0>*ͪ'�����族����k�{�9����c��R:JrBwୂ����1l%ѯ��Y%&t��Ls?�]*����Pѐ��{�ЙG����o�76���X�{��N�l1'�0#���`"`��N|<�Z�.=�K�"���u�'�)X<�T�1��3��1�U�r�t�)9��򫎡�����b�[�-�����(tW�㇮��n;4��c����Z�^���n�:��i����z�0���"�,�/���,��ΑWGF�jc|��^�E�=���X�$�b�:�"��/������#�mD����\��.��A�̻�h�e\���ݏ��n�>�6�^�
���6xs��썲�T�Gy8�ݚ]9XH^6��Uf#%6ֳY:���Z�D^��=k;�]8Ƭ#X;��'��	U6=�������O֪S3�`��˼��������������{?�}�+�
�VVVދotDa� �B��V]-��vx�\�2��K3�S�|!����e��فŁ1�m�с9�%g�ug#��Q.�=/��s���(��F��#;��	���!�g�+�Oq�W6�����=ʀ�ޓ���XE���۟���U8m��>�ϴ��B=kⷮ�_�J�ସ���Л�`�2�����5�-	�����6��>8��p��=�-��Qĸ�669PzDG` ����'���$b�}3�'�Q�w�� �T�'�����EvnN[��aY�Q��H5��&)&��E津3ξ?�KRy����t��W���������E�pі6�?~�`W�(�L�>�Q�������y�>�d�M���n�����G0!�0��k�A�1�6J�����MS/��������@��Z�ܷ�͠�v{�r�e-Ɔ��(VT+l?}-V�?����*A՚������*)QF���;�6�|��K��T����{��`�`���Uc�1]�:\����T����ɷ֊�Luz��.Ĉ��b�3��8���F�<�����t�28�:�`�2ӐGG�����?��9�h�~�u�K��!�$�c����
��f���$��*�<���z�Q�i�V�����?��]���6���?^�b�L��,���ks`{�^��|p��f����ֱ_Z�����N�hߪ���*|N�ѝn	�9T�7��d�nf���)	�l���0�����z�H�4����p]�},γK�v���>��f�E��aml,� �ØrRX5ƒ-�j�|-��&����=�������4T'�>��c���9��3|�)%��כ-v�n}�9��Q)9�١l/b�`�`b��K[g��ͼt��}�����B�!�z���|�r�l���i�f������)���.c���X4�l�����%��:W��#C桨�A��_^9��[������4��y�Ў1clL��5��d͌�;����\�
�����t�0ƈG�����ݩ��ֺb���=xr`�X�{ȂG�˔��9�&�0@�^R�d�����z000Q���@K�C�28;Y�.����i|e79{��Q����l��DJ�$��I �
����,����r{ؔ��C���7��_2�|B��ֆ�����P]~���=W���??��:��Hⓞ��͂U�ݝ����旖6���'-uab�>����ͯ�ƈ��~L�-�c:(KDL[*5{�$��i�gw�+�⋆�`o�|����n��"���5�����\�25�Wn~���Z�˰ s�[���e	\X�������:��~J&�h��.3���\���6'����n
N���P�{�k���'ˎ���E���wX��x����~�-��I��L�|���������=I}����>�\��!���6���g��D�x[��V�88>�� B���8����/��&0�Fn;��<w9Q>�0���Q�.�KCk'���c:(�1L�	�V���x�CZv��a��`�A�������&�Z#b��:q�;����B���:��~D&Bq����5Y�u�a���ٟ"���'�pM�w���r�I���i�\�冫� ;��c�(��1�R����ES ��a6p��w?�7�j0y0G0{TG�ع`��i�Y_}	�"�'U����<b��Q��v�>)�M��ٺ�s�p�~C�&F�m��1�m�}n�ib�8�Ů�B�/��������ϕ��cYo_�� ��G�bl`����~�Q���m��b���Y.�<�ޮZ��0����b�`��:1�	�KcJ��-iIp}rC�ml�a�bǭd�0�AuՏsW}/v|�1���{��+t�k��4��k��� FM��N��c}([F�a^������_yŷ^�@˪w1$�l,��b-���[�\��]���9Y��79�}�.%��#0k��(�zsk��%˫�Q���kE�SK_3��Y���X	��ҽT�Ͼc��|�*;��Ƽbn�0Dg�|{	�
��XX�teKd;[0U�v?����`-��X|-֪�>�f����e���d��ca�rna'���3����g�%�S`�`]���0u��,aИ�3;۹U$�x)���������Ȱ�.�m"�	��$XXXX�`�ͩ��~qN4jR\�/+g#Fނ�	�,0f���cC�l�s55�!��okg��-%�cMlle�N*������lw4�J�RT��P��%�E%!?��&Eu����c�Z��9P�Y�$|�ع1Ur�=�0~�0�1�/`_{U����	�>).���Υ1�|cwG&>�͈r�W�2.)�����TM�����ӳ�t�#$��u��Q]d'�p6D��?O����f̻�8#g�s؁=ٮ��z7�o�4�e�	���)�=�S��-t�\*���=qAEVH��+�q+��+0�[XkS3�8q�m#J]ގ�Շ(ţ��)TIgGQ�v,L��N��P�3���t�JC��V[��	�������j��y��>#F
v�	l
���ؓ�S9
z����U�M�mx+�E���������q]_�'3.�Y��ϡ�N�Ǯ�"�{k'���LQ�o7��n��
J���-W[Y&ґȻb��N=������@�-�Lԑ���mAg�:�k�C SW�\7�a�1��`�`��n�Zi��ɡV�+�D���Bf�HN�ف������,�����3���/�.�W���"[��
���s�����	����J^r��&q�p�yÙ/ֆ������4�NM�F,l� lL,l���T�֧|�Yxf��֬1c~�ָ���Z�Q��}I��C06�4�l3�(����*�;��`�`j�-�Qw�Y�[�Y�1M��*����ۿw�]cldx	V�GV�6|��(�t�`�R����n���a�+���O�#g0�D0M��H<����v�������s�w�TLō��R��B�5�������lԷ/Q��pݧ�!�!�i����z�{aD�1�35ֻ/�:�(a���J;�����C^EaZ��>U�km��2�X� X�t��\��L�M^�2F�P�_�O,lk�`�`��.���2i��9�\R��H߫v����6����00��"�f��M�G�p��H��K t|����xS������0��H�n���G�M�E��+c�6�>��ɻ����qqo�".��#qk&`k`�`y�cm)x��GJ��>;_غn*�.k�Oê_����5tGc�o�e+�Yoւ�j�-Y�Q���k�I���Z�S{���r L��e}�Շ;�z��'7%��x! aٻi��W��`o���:�z�
�ш�^���VG{��D�|��o�b��w8@>u�M�b�1�X-�4�Og�����Ezؒ�!�P�U��d~\��Y�v�������`^]s�����'�Ȓ�^�9�����F	���F��3�_��a~`Kf�%�Vk�	��v�k�Y=�%SCۧ���75�Un�l�鄝(՞�2�L
,�LaY���
�?5W�l�8|�Գ��$�5����ר�SG�$b���y�}�X0K�MSI�8�&��=�`���8�S�e�N�a-l�3��5'j���S>��O��[_FBÇ�/ֶ�.�ա�߮�ibm^�����"B�#?i�HL��$���\�F����{;f����Rq�t/��ʺ*}?�$��0�z0�Y0vTw�}�`���s$Y����|���+'��1�͇�����O���r�'��k#5;h+��~9^��"e���m1�hv:�K:�2;�'b�M�3ǫ�Z��OS.�(V}i	���(��10}�e0{�u\��z��I��3!V�"�F�[>�x�X;&
���N��������;���'�0W7.�l����;��/`�`v`w�J������[�=��N�#��el��Y/s0���q�����1]��#�vl�����X��0'1i��n���1c	��l��-*��#�	6,w��=t�|�A�>��kW�xIFw��Q�冭���,֧���گ�do��Q��!�5/ո%�g#2?D����)ڒa�Gu�K�`�lm+}�����h��7Y4V>��F���������+�Xl�nWq��\�IMfi���{+�V~c�1��"ݍ]���ȞB�O5Y��_'bd�_2M+��т��M�q>:��� ��ɘށơ�C��F)��!�ܢ�Snc"��j%�z�s{�� l���R�r���X盺v������"�!k�`�`r`S����^�]��=�6�0rʜA��R�������ݥ4
3�d�G.���=��擂X�x��D��8S����ղcK([@l��j���̫Z�wE���h���H &F�VVv1�#Xk ��&tz���)y�`���%�pG���=O��_-X� ���1�n�Ҽ�J��5��gtX�>V��1(��Yz�R�C���<1/U�n���!�:���!遮�`��������������1<��Ki��ŭh�4Y}��`4`�`�X{��2���"��%1��9/ ����⴦�Z0��B��`S`�.���	k9���
_���̥;v"�+_'�iKk��;w�eC�a�10-�0W݋��x������ĚY�[�U&���������00R\�4BL�`-�P�	��Vf�ms5bK!X���Gٿ]��\��~�Xb�+�Oz�7��"���|Dl&�Y[p�:��`t-t(�����J�iR�+��[t[<�z���l���E��%0O��17CY���bOL7�
3�E!F~b�y��b�دsA���<9s�1�)ּm��d߀��]��M�Xc�YZ�{�vA<t���(<�j*��2�Y��Jqw�����)0'060Z��`���J��~��
�ABR��z���},X[��v�a�����c��ه�4^	���N���5!?�VƋ2"T�/�C+8!�c�h�,��b.��+*�}?��܈�������$Q����3w�K�o��ߚ���j߸"�v,L1u!���逝�+�=���L�g���#B����Y��LSk���t��ύ�I����&���ך���ը�WY�]'bOb����%V+Du���މ�X��-�� ^Ŭ�_v����ܸvl�3�)ؾ���1bMs̎O���˚��z�ܬ���(cM1���4��l:J�>��+D�g/y=�Y��_�u�V�\&�qȟ�S_%�t�Sb��LB���朶Jy�����T2��M-�K��(�F,L���'�0�[���9�r�#���4<[�.ы�Clmk�`�`*`}�c�l�G[��Z���V2�Z�0c�5�C��!J&��Y��ӻ�w�� ǂ�R�����Q��[����!vg�����`0�ol(�@�uONך�ˉX��J�P��qd�`�`��J���*�B�X�Z9XИ��ɔ$�U�c��
x���Η�E-H2��2�)�����c��[�PJњIwv�_:B��<���K)E�83$�6T����M�;�yS������K�BrE
��'�-�ɀ���;Vfƿ��kOr�����(-uy�4�V��`�``��XD�r"JK m�g�o�<�Ѳ�j6�~��ԨL��_#�n���̨�����{�-��K��x���׻P�>��й&M�xj�Đ[��{�O(�E�������g9��\���P���)���o�`q`��	?�Z<�<X��7�w�t��xCߝ��b����eĪ��VFve�v�s��2�;���_��|���7�4ׯ�R;�X��^�z�w�e}�|����t$��Uyw��̃� ����Dub��) sݾ��`w��]��:u�'�E`A``�����kk`-W������֏�/w}.�=[c�,�&�����������g�����V������|��^A���N�#�,�
�-/�:X�3�(�QP!=������"�����U����:��TY�bl]�c�x��4WJ��p�a,�i%�P0�}@u��Vfb�sw,�9�ǚ_�W�ݹ�(�Gq�s5���Yq��;v	eGS��l�<oT9?ڰ�gr"�"�NSX<X1X0�bo���&�����B���ұ�z�Un)�=�eUg�6�LeFk���t�V�\��\<�ZT�؆J�"-�zN��*)�c!Z]��S���yJ� ׺�c�n���3>J��J�f�4LSp��*U�y֑�`M���j�����!�G�E٨6�k�z���豩F|��cD��ϭI|SE�ߴ6���ʟ:,���lě�z2������Eߦg?�4��b�ҟ�u��y�o3�.��'Yf�t����4��:���.�O�yi@�~n}n��ʓO�f��7�J��h�<����S��'h��v)��Y�N(9��x>CR!p,jh�>;�rC�5w�<۠�D	���V'��W���(����,�?�x9h���w<����q+{���[	i��2B�eF��Y��#�*RJQHRVY�ٳ��Ψ��{߹;}N����Ͽ�������.8�2[��E������'/��<ɧ�m�2u?��TD���y���\pzh7��C����Q��Uz�����bB%Y����>���[���J2#:T6�]$�Ҧr襼�{{��1#O�X���Zє��돨0��R�jN��,oZ�B��tY���K����qJ��ݻ�Ǖ���i��%�c��i���|椴>]Sh�	K��x2-|'rҒ��뢏�_�NT�Qu�늏D�`+	����|1?��p�ho�<q^B�۵-;�	�';	F6�U�gW��p�~-��5����B7�Z���#��,L��/��d�c5���x-��Q��R�i��D���y����X���� A��;��9�1)�٬ԵEm��[ ����ӷ:^0�ч'���7<�=n;�Qȉ���=�010S���G����RCĶ|�*c���b|C��p%v0:�0����т���;�m�0�W����F2�e]2r��Yð#`n`�V�����0�GW�FZj���%�6R'�Kv���%��I��[��x�U�i����[nY�S�k��:�bofN���Հ��������X��@虥7W�_6D)��)��i=n��k# {VFF�ZXX��7�ć�̹�38�	(cq2=~�7��-��!	��
'�F��]#���8�;��:�`�`{�l�V����f�v�t�~�g�����=��o�F���f�3rE1`�
^�1������Ϊ����)Vt^�I��;����v �`�y��l��ݹhw\����a��&�GK��]q�Q#h�S��OK�&b�`j`�`^?�rî�����5Ҩ����6�ަu`��[V���>��&F�0x��T��E�w���I&��z�s�r��,ȗS# �K��AWW<.?r漹m���$S�����P;v�N�邽3�1�wn��I��Jǹ"�ť����XX1�5�F炿�9���Ѭ�É<(~L֌K�̌r7�9X5�тł�����c��C��wp�%Z�J�2X!�+��	�X�zb$`�}[�<�!X0Xo	����3����k��KT�s>aX�)�]�N����ȅY�G�U�y<��k'�u�T��g�X.X��.0G0R�0a\Ԕ�x�Cݤ�����|e�G���l/ju`;�f1�:��.����ɲ������M��o^	\0�	v���U.� XX3X��_��SI�XP<��m��h�.Q������`�������0��3��[#V�%	;v����S�yD���v2�A[��`�`w�>����"bg��3���H+�$?�%�|*�	�
L�>�L��4#�c�c;;4�`�^GK������!��``�`�PkF;����d�қ��ȩr����r�cLifg�|`���O?�=�0�KG���墜�"�����8f�ަu�Y�����-��#��=NF�l��tHB�XA���Q��K�D�Μb�i9`<`H���H�X�x�썝�U	?0>���\������l5�0��R��hb����jR[�=�\���i�`���BM�v�J�J�tr�^f��::0���
���������J��/�͙8x�}��P��;Y��W�:^��l���*c�"&���	���]E�ƶ	���:�{O�=����Þ���
��!FY�6[-�X���{�h�V�Ɠ���`��O>�F�l� ��	�G��:����M3��%yU��!��*� l5q{���]X�%���tB�����D�D<eQ�Bj"`�`���DQ���q��?b��J?�x�s*�A|�z��'~7���0FlZ*���9���k�'��;4���N����)�8��/�ٱ!������k�>���nBS2�
�a`<�n�郱��u�{Mk�
q7|p:��C�=�8L,�k�/��}�0�����"���o��m��^İ	����~?�X6�0t�)1��-�ɮ{H�uuw�]O�;��w00�ߌl7b�o�l"�$3<.��;M�؎Ђ�ڋ��Z��#6�	���ѭ2Ag$��{��w꘍�UBę� ��'�M��}İ)Ԑ.�N��Ѕ~���:�Q�P�c��V �����{;��U����կ9�/��繹I�|�p��)+G�D��vۭ��V>1(�x :W��z}�BE
�=��`4T�K����j���ia�Rt��/�I��F-�G�1l/jB`�`�0:Ė�>��j���{ج�Q1t)e3H�랾!b3`��A�`�`,`�`�)[֥%Zja�9�����J���'��+���M�)�F��PԊ����&Ő7���C��JY�0V�T��Sc,c�{��Ll�t�6QS���F�l��9��.A¤���xr'��=�D�b��P�A;˷��H�
&�^�^q��li������K�Ԃ�2�j`��>�Q���߲R�l�v ƞb�3�s�m�&���F��Q�tQ#S7B,b���>��m�ٵkV�����=��Z�"j�t� �˺�e������c�PF�b�H��=����cZ3�dyV/ 6��:c
�����jv4�7-Y�6��M&�ѻط!�f�e������f�
��o3O����zk恹����4/�uUM#�)�[3f�F��,��CW2�x��My�lC	��>�Ɩ*^�h���LQ�� �K6Z���uD2�ܚr�Q�Z��#�$��5>�
�n�]� ���z}�:R0cAg�xrE'��˺+t�!��`K`;Q;��E�&bZ?�QGDe�E�bpr�v刱\�\;X�;�}��i�m���n�� s{g�W9�dw㈴C����2�}��"�D�2�2�~ZjDHw$x�[�(�H/S\��q.M��Y0Φo���mj�U�ႉ�̀in�<KA^��N�{���!�A�:�|�s`����Ղ=E���>���\"s�8.0u3��Tc9�>���`x`�i��`$`��L��S�5|=ՓS��>=u��fD�8���f��U1��v��.�)����(I���]�!%��O���\�|�|h��F�	�v|��Q{v1I��o^��/l{u�|ֻ�g�q�G`���Q˙�0G��we���^���}5�����ݬ}*�}��",��~,,�q��-��V��d�Ԣ���^]�ǵ�OΌg�I;Q�6=щ���/���m{���k�l.�`z5!0�)���÷`�![��Z�ji`�`��pIT?��~^h)����U�]�A���S�OxǃX4� ��K��s��C)�q��u�}�6��Q�V�è-�Q��a�
9�������k+�L$~�vۓ���<�o��[K��k��f�0&��\�o�f��������� �ưn�r�=I8��`a?������)L�l�y�^}�vL�/�v'b/��L��^0^�>����h�Qj�Svγ19�eb�.0F0�`�Ͽۏ�U��KW�/��t�h��s�}�"��=�S��x0}000ew�4$�]��b��]�9V�$>��v��+�:X�����ZJ7a�o��
F�ە��I�>_v��[�R6��	�������e]*�����|t�}�~�����s� ��q�c�Rw��`�O�>������b����ٷmT]��6����&��w3;��nVO��ao�r��.��v�5� ��a�����]�p�F,�l�������3z��)j��N� 3s�-�e`L`=f�����Y��w'ޱ�/��[}4�IEZ?X��mj�Ɂ	������4����>OgK��n�DȾ�%l���񃍁͢��6V@}��`�A���^�]R����w�W{�y"�&��1n�0s0A�N�:�]m��"��Tќ��g�uX��6&&�a3`'{�w0L|Ǟ5o�L��fqQ��BR������ł1�����>lu`^\�n����%���xY����i�o`�6�L�J�1��F�1�@�C�q�n�$��M��ǝ`=`W�D��@�̂h�K�K��7���|Չ�`[�"iϾ
c�	�-�䀘3��#�%��M�Lx����"Q�쉍O�v�%GL��-���N0:0�v��Fo�%����̷<ybc�p�l/X��,b1L �KvYqs%�I����X`�����l�k�<�b��X�#�~��[3�\������{JE���	�*y`��W$��Z0L��W��&O�W�{��������b�;�I��r��>�9�%��2��iԽku7���
�С~d�6��j�`������K+ ����>3�4�H�C�,�N���k/��N������2����1�{����l���'���[j�V@+b�X	�;�>0%�T���Av+��I~��/E�U���΃U����ֆa�`ш�?;�f���e�%Q��7�x����c��;ff��%�@gpuF"����i��3�ԒC�
`�`�`g�������ú�m�{����v��¥�w�w;.�3#&F6�>�	�]ع������:��c{|5�3J�5��z0L��^9��V�4�p��3DzJݢ��/��Vc��t��l?%�q�ـi���n��m��)�z�>��v��BQc �E�\�@�.BOlC��C�}n�u���e��o�7��[�3�~a˦X�ߏ��1j���>~n��5:^�r��_��f�е�����O]�Myd3�3zɲ?��!��[X<�;0�:�g`_���D��.Nu�>����鋇��n�M��ʙ��!]yu�jo��W�\����Z�|���d׌��ȅ����ϳ.�zo[��eC�T�����wQǌ2g6�]SR`�``�:k�H�T�p��.���t3{�Y�2DBh
f6f
F�Əl�]�yp./1��|��U���#X�s��`#5[�i�~��ΠC���c����>��������'�dZs���>ȑ�(=ѣ9����^��kC�������lQ]�cym��*���k���})J�F|~̠:����Ϣ�My��R�)3pOn�\�j���$%c�܊�M�y�&8�[�|d���i�8Ӡ5��yg��ᕆ���O��[9vE�6��/�ls�?��}s�(�T���A���:�7���V�ğ�~_ȯg:_]O>��|�C��^n�\%�T-�&�qUW�"�9�V��c�&U�粈�u�3�T7�"�4�
Q��m%�F�E"$�{��eG'��%�񐢣c_Q�v���D4}�W�w�8��QR����h�U�/,Ԕc�OSeM+�S�L�iS콄�{cu7��K��џV]�DX�(;.��g�4oF>j�q��?l7��2�H��.�:�x�%���ƒ8�g�϶9�%�X�+�Uɱ������~vj�߬�,vx0�9��ǣO�|���S}+%��� [Am����.oK}j�g�X��2�R�X)e��A���KD�������U�X�KQ���;6F�t%����bE)��ai�X���K�����|�v��H��F��\�,"��w
����Osq�Vo?�M�TI �x0f�T+;sM��<�+�"�Ya���w٢�2��-+C�b��Ö%�5n�r|{���M8�Y����O�XG�9�Q�[��6�����Y����8g'��-�~�Ӟ�F_WM���������>��S��%��73u���3?��^�ȊY��;sS.xN<�b��l�aM``���I�"�6�>�=.x�.Аj��\���W�JU�ܫ���*������{?l��/��m�/E�Bnߗ��8�e+4�ݍ�ȷW�$�3��(��⤿I�o����fk�`�P��-C:�M{�-��ޡ�q+�{�!��0��a��E�W�![fT���T�|V��{�s��ֵ�W\(�������Y������-3������������]yJ��o�v��qSdi:R��T�et`���n��iژN3:_���e"����R3c��ٞ���w�푭�T8�<1|)*5�o|Oe� �y0F0�B���q�=`�`�`8�uD��j�*�"���PK��j�vIk�O�&�*����'�˩r�A�"	u��F�&�*���ܟD3RAƃ����uᅳ���l���sy�Z�z������m�f�$�$M%�G��5�i����"w}4f��kwI��ҤU��=�S���C��:�&��'`��i��%}Gj&Cb�а��]=���1^ı:M^q��D�����/G~��3�=|��0��i��F�䅟��E��v��7'��/��*���:s��y����>�6����4���u?�y���ﰭ���yI9���j�E���͂>J�N*��81�zhXp�]���ػ.	���b�^��跈:�����n���3��P���SA�(#�V�j%�gT.�W�ac�js^���v���x\�$�.r*�/�����4~?���f1�5M����.a�\�W��~���"�Q��s#�t�?�i�ۛ�;\C"88����Tݰ����0�M���LY8�WgC�$T��<=��NB-�?�y�F0��w���㶙���U��Ջ�
�3ؘXH��5���K��յ{)?��'���a)�el:/�o<x����3K�ٿL����2�-;v���/cy�4I�4z=��v��O�4������y-�L�:�wg۹G��C��:~���:f���3�������n���H�G<�C��s�ꏝ��cwe�j���NC�ZY��j ���-;��0V���at5[v8L=(��Dn�F`����
�7�ؘ�C^�ݗs�=��Kܷݵ���G?��N� ��M�8�ȱ[�β�;�{����u� !~��ѣM
v�5<�����_%Sm
CJ�^��tDs��_�|���[tf��*�щ�1�7G����������m�j]7ޮ���
t��:x�'��/��>�������i����<)x��d�����]_��U=���4>��$�V��2���~��ZW��y[�k�MH}���=fRYκ������}GM�,�td]xZNv�+F~QA�n�ϩ��S�Y���c���,~�5C�Tؓ������9�	�p�����?�Z��t���a�]�Ą���������z'B�����1K=j���Y��>$���tv�m'ד�����Z���qd=�a_+X������Mk�y˟�Nť&P><��50R��`�M�����1-�ɌQ�{�~�}�?�JY�����?�%������·��5��N*1�U�wJ��uC����1�]R85EmY�J�I+�Y|�<� ���������)�b��Ȑ�<69yh�����?ٗ�?LD���~(#��Uq�y��ӄ�E�P[�w:��r��
�2XFw̐��F�b��gӃ��ܔ�M�+��`q�ﾮ�&:����n�W�}N��y��N��Ǣz������o���>�,.�gW���Xp�Z�,S�{������-;W#_�	6����n����w�ޣ�s��w�d�b�_�L�[��RJ�q��,x�eo�Y��ha���Ĕʣ�:f_��X�Rcͩ��l�1�7I��V\��o���"��Q��A��!}E<�h���X��c��eFi:*�ʔߵ��Fg���C��BEMn�N��Y�}f䗉n\�yY:4.�_-�������
�·I� �/�c�,���p?��E��ա�6a�_S�hd�>�y���u�E[�#����{%������q*D����D�4��6��B,�s������g��Y�k�=�wn�D��Ƀ����AML��:�ĺG�-����3�v��ԏ��<Oi�߬vO\�!U��H&Ko~�2v�[�T����T�:+3M�k,��r(8.:.5�jos���w����}p�D�-�Mf�ǵs��0����V�Y�S��k�F]]
��ִ��F���=<�j�wߴ����R/��Ysvbc>�J��8q|��gq�mg�Anm=�F��E9�K��$��oj:�(��FR<����2��לU�����ؘIm2�#e^��=>�q�x[gj`c55AYWiRm�:�v�X��d16f�X��n��[]�$sKZUI��{k���βΏ��r�)�����}l��� �%�H$6�W����d��`lL�kV���&��S�a%�SW�1��u��� ����Q\��3��v먃$&�����&�t6����X�v}!�9g���Z�9E��x�|��S�Uy�KL�{\�/�~]��.!{��P�Z4[C�l�ʼx���q[l,h��Bh��z׮��fQR.rŮ��z#u㞰�m�l����<Q��S���5#�)�\(��!�Iה3�ؘ�[����-��R�p�o�E��σ,~篘-Ue���=쀍�^�rLQ����H��h�Hc
6��X|��v!K��=�-�AG��l�+9��A��Gx��K��I͍B�3�!�p|����'1�/[v���&�X���B%Q{�p}���w,�G�acD};���Iǩ٠��u�7�H<�����dƍ��^˩oQ�W�1Jա#�k�cm�Cwjy#��\����{�h�X*-���b����s	66�����A�,-�P\�n���z�����c�F�A��	��|�R����X����&�,��YȺ�J��ac9녴"N��Y?X)z��<=tO�;8�j�$���Cb�m�-�{#�갱��� u�������g�3/����
�F|�?+�N�I�}���D��}{�R�J�F�|ź���ɤڴؘ�i<�RE%�E�՝��T5�����d�kQ}3>�4��cg:��bcst�2WK��m�0cj<���z6�}�Uý�2���R����N[cc4����i��}�+���>��"V&�}�
O���Q��K'��	5OacoD���?b��{����\���E���O�2_Wv+ *?0G����.���]����5C���l�v�ͥ���\R�Wˤ��݇��bc�DI�����2�����Y&��`cڵF�O^���=�(�h����46v��17�ӏ�F|�|J���vJ:6��v��h���UXV��aD�I)Q@ZI�N�.i�;E�A@:�K:���;��=�Qg���|�r%x;ϰ=_emU�w�O�/�.� ��_�fN�4�R?�TJ�9bտ b�*ؐGv2��B��!���ρX\]�����xH}8W���\
9 �1.���m�U(�a�3�DxJ
�1����Fb��H�N�
(��T�E���r�wxp�eA�T�4@�u�����k�vp�ýC?���* � �d���0������ZG�d�P 	��UaK�%�G�b.�ȣ��u9�0�V���wL#XRH��� byv����$���t�-.�:/�� b���(`'͈�^t+{���G 1�<%�O!|��X���ƞ�w��1�f!�h�"Q
�Evr��Z@,�1j	˝��b��t]�����U��p=j�ƅTS����0?Գ�;�h��]����x��p
*ͪt��i���g?�e��a���ej\
bi�2��������u�J�X^�U�.�����L�fEN� kV�N���-F�8�tOH��zĸ)6�L�7�H�)X��S�#�L���nό�d:�i8��/�u�W+]���T9�j�����7|�~R�Z�Z���T�o��|?I�ʖ2�/���������A��_���x���7pS���$N�����h�7�_ɧ���c�Q�w�P0�K��锾[I���L���+�lIΚ�=���Vu-��h�96��9�.ʶ+��g�����H�����!:�ҼAx�7[�c����4��9?��f�}���jvA-f;�l?�PM�O˯F��Ѝ+xžu�|�eOAg#�O2�j4�ۚ"{��#���%=e�)�t�:���a��Т���S���^ۋ��J�)��d���'�~Z�]*����G���V�5��Yda�~�6���e�� �mB>��s.'��^���}�Z��D��k���I��zn�9�+(�T��䔦w�(��6[J˘����)J�g�����pߗZ��k�|],57��㠻�'�����\U��8��<W��6y�ȋ�Va�m��6�L;7͖	ݑ2��9�c�T�h��=���fNF(S`Go��G�ǍE���~X�̄F�� �o
|֯��[��P��:x�~��i�K�{Z��Z>Im-0��?�z�bP��7f=c������`��+�c�r�*D_��j|���<��G�Q��}i���
�����≯�@;��&��
gw��q}���O�9ie���*����V��Q���зhv���A;�T�8�;�t�|�aI8��b�Ag�׺F���9�V�+h���+�Ty��x�s�2���������>�n�.���LD6R=�_�渒i���U�/���%2����d�ShWp���`�~��0�]�hR���NhIA��RB�P��XJ��}d1�2�.9���f����&�/���(O�P2��A) ;���Vs��R@�;��l�EP�bM���f+v���Ϊ��c��H���\�j����R��}Ʌ2�m��J�i�j� B�E}(3�l'J�cw4���W����ã�����/�ը���{ʟH4W�~0��h�!�m5��>����P���0톓ao�O{�����`^̮,�E�K�]^R�X~�P¹�_Lb<
esa�7�Uو��'(b)ъ>�<=���X�jp���F3U��v��|���m�����Q}�B��c����v �W�n��EA�:��?�_��ĉ`�%f�r��4h��=b�&��뭧ڊ9��V�=>�~��]�Tr��+q����?:�j	��H�w˭�tG�|���������g�'C
�z��z�jI�c�o�
�C��a��k�4�+���0�u��4L��?m^����"興���� ���?vH����
i%>�����߾�Ni��֝ք���#�[��Xj�xSG��Ba��V5E�Xf언O�E�����W��g�TN�Ǘ�bx-���Sv�Y��e��f�b��7��v	��TΆH*�n�v
v�:�%̊P�4BRAs)y��O��]�>��������q�R��Ic�|3����΅�����JB�%���htk�98�� b� S-�6��3�Р��`��s��1ί�!����Xѳmt��B1p�d[,I�b�,��E!uR�~ò��ns�FȰ�>�
1CD��������}ގ�������w�c�N�u*x�'�������
��a�p�쎶���u�Og�f=�!BY���i�:|�e.����'���SzۻL��{x�)?�����z7s�x�Z%2z�d�k
}����ZJc�BŭQ,��L����*�4:7�>$%=�>ql{�쪑��|1��Fr��kא��p1Ss�悺A�-�crbj�@o���Z�%u��$���N��r���[�N
�����$KK��KY��j����v�������X���1._��P�2����Z�>��U;g�G�ۣ�&Rx��� w:�4���	:��"U]@sﻝ?x��ME(ǫ�s����ܣ�
GO�a.�_��϶���E����"�:�X�`��w���4V+ ��A��gx���ڏ�/�b���bO�)���KcQ��(�>K'`�T��aF�O ��qYc�vɝ|��vM���9X^I�&m´6J�����ӵ�#5�d���P��r�=��zOpHQ�G��Ղ�g�i���(�)ۜ�?�g�����~����˖k�Q����D��@��c�������R�϶�$)*�B���'&�3�̿/ю- +ɗHc�z�H��OM�P�I<Je0�:��e�U�oō�j�+.��r���7!�}p��N���?��{�作���6γ�W����&[���AY��A�=��B�o暴�/��Ϲk�"bxt���T���SuBvCf<Hf��a,^~5���9Ooʅ�0�M�}��u�d����k�Bɢ�C3<_A��Z{���.S��3�B�>8~?4���7�u\tؘ�&��`�>���>m7�X�]\�Ɨ�d�9o\�}��bd8%�U&q���|�&�5��6�dx���"_����a�"*Me�˘�;@~F�9�X��|*ۖr�Mʲ��cHG���7�)J������<�����-�"ӲS����n��|�X�'k�-��eA�%�
�a���M�Ɲ���+�g�v�y}�)K�!���ϖ�����t�MG/�bu��/�����*&�h���xJ��V�f�J��rv�a(��Z�K°�V8#��Z���f��Cv&]�ȷ�������f�A��dl�-�G\Wm��<��w�(Rr�Q鏺�X�	�ʸ\�ܮ�v6FN�R3sڈ�[�UP
�v:ڛ����	Ͽ��kp��bb���P%�,�YZ��*��HR,L���H�l�%_,0�f�
o�B��鳵��:���T,_?h��ko���D�D�.�_��'�����.X�7|My��Sf4��2��B��5{�F�p��8�w�_�ga�<�Y��:[��Os�L��oz��P%)�����zg�y�条r�9��}�
|j
Y�
3�v%�J���/�����L,�1�'��K��fZ�MfeK��3|�ϖIg���
�Q�V"�{��RB�l�a� �蹎�6�Q@0lΞ*����T�iU�.�Ȕ�a���S޵��6�2(9�5s����o���|2J�����UC�`�Q��f%�TĹ��LrD��/�r�]��!k�訂r'�Nt�2����j�J�;�J��t�_��TN%��������_̓��� !�M������c�/���5{�ǃ����x��/��������r3<ns�ׁO �7����/`ɉ�ˏn�Q�?�l��o���NI�Xy��MX���fߙ�$�������MzӪ�$h��A���0�ضYĴV
e�,�9<������P�g�+��T��V�Y��~�}1h+���~�F	��A􌒨���@l�	������Β�4��2����5� ��Q.�����Ql#O�pp#�?Ss�7S�����>�_+�儇��pYt��]�	�,��ъ`Ke��dja�<l}��R��+o]7����t��OBz��urVE�U�Y��A�Ńt��D�@�Je?g�Ἃ7qA9��]yD����2ͧ��I?�w�g��V�p��NM� ��T_�[O b���SZ2���ع��!m��l�W��YW�_͎Rm/�J��G�9��6��z4�ion�/ްq��JZ�<,��b����|P�6�(�ឩ�J|����L���t.��l��pGR�M�����贆��
]��ʷ����V/��n�	�Q;���d�6~�:k˭��`��a����dF�h	���y)Ü*��o����ME� 1M�O�(������ŏfʞs��`KsGAD�!��N�=xQ{� �9���C�+3�e�������;A?�
{�� V��7�"Ď��z̄v�hb���_�g���n�E��M#<&�Y�u�< b4����l���\L~���|^�@��)*��,cM����Xt��m���ѷ"tE�[�Ar����Ę�po�?H�
Ԯ��?W�b6ډ��ftV����,,��X*�9�RՈ�Tv^��aS�6�)ot28�@�Ԭ�-I�b[cKl��ov����(��1|)�줕�2�,���7���@l^L]�w�|Z���fX�vC�5����"ت���g�����ut���@c�1=C��STK�>�k{
���h^�?��~��M�_?�)aĸ�?�J�x>��\���/s��{�ܷ!��Ή��uK�É^i~�b�V5�,ie�<V�uċ�Ga{���x�N"�](+K�b��?u*x�L_ĩ=Џ+7q�\��;�L���qם�=��P5S:��MйilAi�$��l���IY+�Kّ� 1cj=d���ȊM|�aڛ��0���Vt��D�4u.�ؘ|�!��&�dc^�:V�5k�b��a��b"5��}ጬZ(�T�Bc�@L؋1�,��ճֺA6���lE 6����Ȏ��L�sT�P�F4'�����6����3�����'�籶��}��<�4\3q5��%�@��|l�3@��A�M���ǆ�S�-{HD��Z��?��[��ޞ�`��}A&���0h�(�o�F1o��8\�2й?\i�;�P f�P}3Ld�/[�F{�t
VS��'âX�xc/I���C�#:��fi[��<І���d�%G�X��� ����g���T�Ӻj � �H�1>�h���#g?]�-��6 ���0�i~�B���)����e��T�Or���mg f}=���R�$8��j���Vt3x�a!�AΑ�'m�Π.�۹޷�ye@�(�$C�ŭ�*r�U|����[`�@��+���~b2�V_[�Q��au?���1{����I�D};'4T�o�1d>�	2����e?2��8��Ip���i��o�q�����Ռo�D������ �� ��b�a�^�k,Bb�¸��@w�$�q�ٚ-_H ^���11��p�}�&s.*K�&J��<�B�Vl�W�x&] ����S�π�.h8��E5�%��y��Ƽ*k1�rc4G|e��a>��ݮJ���PJ�����v՝�|���E�5;��&�[EH�������>C ��b�UщM}c*�P �i�F��>��?�x5rs�ᖟ��،(�8�,�<b��9F����#b���ı�oG��XcC{���'�1Bí�b�cA�5l�p��OX�O��ȝ��xK�����2浨Is@l�ՠ`X\�c�a!�g�b[$��s�>�d��tD0��I
Ȇ��|Č����?F���{]��[�~�����A`=��=�Av�����Đo��(��j5D�E�ˠz����+5Pg�C��	�5
"z�?	�a'��k�w�������^^��uc�$�O�q��O��Bjo��ɑ�� Z���w<c�[�h_ZU ���w�1w������T-��v��wV5ϥ��G�*^����[e��(�0���j��Kd;��OD�gL���ɻ����؜c��pP��ɵ�A?��!a������Z"�ت���Nv&�1�	�q� ����C����=;vW�($3����m��i���\ڀ��f��L�Z��jk��������rѹ��#�յ�u��g�xi�ԓ>ky�����a�><f�6��갇��]�A:~����x�k]4SĆ�K��{M"�o�7��S�L1S�l�Lw�b{.eC]5��3-��Da2ǔ�f'-�s��Ue�M�l�E�e�y��t®��J�bi���AJaɻ��f�� �.^�^�ʕ1�H����K�̇�L�bڨ�в�PI.7���RJ8�Q>! ��9p����N������3�����)/�&1r�Fh<��G�;h��d2m��և���L��߽#^Ă�f��|:��[�&&���~�Jb /�7^�8�?��d�t���W�%���-�8R��m"A�K�u[�B/�j���]�����oV�"Ԧjeʭ��vi�ض���%fȏ���p)�c��R{��ݬ~�<��|{B#6�U�Sp�G�v'ʾv��7��kZΦ�h���ßA�����3�ut�W���>�5}�Z��w�;��=��I_d| 1�p���Bj�C��b'ܬӏ+L�?�
 b�!]�I���f���ٝ��t	݈�y�ߺoVq���ד�?)��R�� xB�n;%tS���B]e	3j��,;"ُ ����w���Z�u-6��X�'����zCk��س�wʷ�L�'.T��-&t<.6�x�������,+���+��K�f;���.�K�=,|�+�l�P�\�d����}
�,�%��)CJu]�A섒3w�y�xڍU��~AUA����-���Aky�f~F���x^oX�y����)����Ћ�z����m���:���	x����WJ�T�r5��"��,Xh-M�5,��H}�!�&�K�w֛�D��f�	$$$>|a5M�/O�<�|t��+⤤��C���b7H�n9�'��4zH����py��D�����s�|i%������$l��"��Y̙���~c��"���p��	�D��Ɂ����>���o���"���7B\Xo���8;S&�ɟXrȠ��(P���av�f��������j�Ti=�wG�<�x��E ��[��P�+[���F�"��=�׶ �r�m#��]3Qj�T�by�KqB�w���o��o�2��l�[+6�J����no&XI�I�ot�����~j�0�#���ݣ�/6 ��1����A�]�$�q��Ά��48�p�P%unIȒ�\����Ǧ^�u�nvb�b��'�khÓ���)S�b��n	
Q����'43��3H�A�d���H6�dĉ��56�yk�����f.ƃW�66{|U!�v'�>�I:��UK�����y�f�,%�̇�z�a�t�5��Q�D#HY>���f�/���4P�W� i^s��pt�bN�y'�Bz���21�B��f��Ӡ҅���Z	�=��^i`s��c�Ӵhe�!���M��LT��c��K������r'�g[G9t�)hQ)jqkw��I�$�k��}������F�	A��Ҥ�1�Z�] I����R��,����{fBo��Bޒe�7vD�z���x�ͯߤ���1�h���UT�a@R�����F����T�	����ni鐔�T~gMlg�3��=���=R�[Rs�bO]%�Z�5���/J�n��d#uE���˽�f�:J[/���!���0!;l8%r���c�N�a�gk�M���=�+����pʂ��d�E>&R�3d��0�B(|a�����6�Q4ӥ����f�y�/S���[�(��Jo����wP�@���@7ܡ��$�a*��?��l��7��M����j�V���Ɛ�)Q�Y`P#�_[��>%R�Έ�\r�}n�ÀP?�x�� �&����7���[(�4�R�&"��{��i�C����_x�ճ�noFw���?�s����5��"�:����W��s��X�t��>v��ɪ%�/v�#�)�B޷3ޭ�{�H��:]�O�2��n6$Uy2���ؾ�*ɘ����h��2�Z�ه_-Q�vT�|f���zܴ'|>�~G�� ˿2VIr����e1#�K9�F��b���62tVÏ_�\�b�~5Ɍ���bS��_�U�ύ3�j�Z�X�T��4�p�� �*v��A�''{p�y�joY/��$�rR��Fd,�$��V%�����
�b�O�������e��M�����F�]���}Q-�1�4g��hp����<���u��;\u�,��IY�9/�:�B��f�WhĊ����a�����͠�#��]��#��dAW��oЪ�"N�m��j��7�I�˝����0�J�DΞ�F���U�E͵�����̪bn�`Jq�P����У���Ӑ�\��@���PªS��[����uď��͘Cg��_;牃͡�s	̗c��Pb}�r�(�!��3�P� ������
�,����S��A>��h^�>}������X2,k����X�K\���:���,����d�t�"
�;#o�X���9��A,l�H�74��������K��a�b)�6�ђ�*�<��4����P����Ϧ��J�>�&^BH	a�[#�;�(7�(X}Y���옜yZG�>b����*5R�b�&DG������
�d�B���n�t�j�Y�3U�{�����i~3�h�s/R�B�M�9N�
���]6�z�E+#f9�`��\  ��H��ڔ�^[E�[��脘E���X���ʊQ���$'X8?u�J?���䧣���'��mR\R����T3gu�ʫ���ؼK�"��3��a��q8��?��gE .�GL8�@{Bc�PfoPw��%�������j�l0j�$}�毝-�
3aA��}��3I�C�
�} ��9�	U�Y!��Z���	ږ��g��S��͖�l�_w������H���gR�J�d �m�֬ď���M
��q�WŽ}���W�
D�g�������e�}�����t��"�·K�j����N���5 ���Iˇ����ud=t5-J����F�}�X��wfܑ.�1��|l%)��		�>Q�;�&�����e�q�n��.pA^pXq\��vMz���Ű�6��>�֎��߸���u���}���4��ݔEX*T+9��0��/}�?w��
6��"� '�I�9p�� �̄�-�J,��u�͗��L�?�v�^ّ�)L̟:m��-��9���7�d�n�V����mw�	F����/*/���+p#�Ac3��~�Dd�ʿ5�Q��!$��!�B��L�M���0!��?�$��OM�����^�甆0)� q"��W��Ձ�,��6�n�O�����ٟ�
[�D�ՌH���]��O^����V��-�R�a��G��K��h��!�$p���(+{����_���=��v�:�1����:l��1�oĥ�2�X�����^��?�Wݫ#V�k�Efk:�� �ǧ&�����1�d\�w� f5,':s򫡽m����o�#�V����B���A�T�X��z�m*s*�[K����k�����8�,�^��W��� v/C�A!U�re���'����77f�x*�Xu��Ꞣ�\W|�������T9��;�}3�32���d-�q���m��~�!��҆o����:��nu��1��a6a��<�bt�i�b�VZ�r�e�{yF~w������C����m�K�á8�jc�c�QCʝӯ^��$^.	��ܹ(N�t����N�u(;%��n� ��-�77���9�%�I2�4��eFc	xQS�#8����)n1�xg��s��}�ҍ�G��Z f\���o�hG#����4%X����3��R�b	q��Lpi�X�:�H�Ry:������a�q���9h�
�Ψ���EbT�%�0��7�h��f�P ��LK&B{<a���>���cV�� ��`�+H�d�PDF�H!*Wπ�*�
�����}?F��+�٭���婍@����H�=Nuy��'�E�ۚZ����	�lݜ(с� Ń��פq���I�%ݪ�t ��sa��n��(�1l"b�Dтm{�T�:�dr��h@yǋ��^奄^��g�#}{3����b+�L w��U �^���(�ڥ}�/�'Bbau�	�>�X*	IP$�!.y{Q�XlA��xՊM���72�IV�aì=w�/�aFz�r
bO^~M8z��\9Ѣ����Čq�B��� xP��31�ÀXH4$A��pW)u�U�E���1�qM���f���}A���uBP(	b���%�����H.���-�A�v��DP�uߟ�y���-�����}��޿Kfl��Oͱ�O��=�����>lC�'#YwŖ����� ����o�Dە�����r��� Ė��GN�v��1���5��>1M�6�d=��v�pZ6{iї� 揱��&�F�~�Kݽnt������{�'T�V��sЗt9y���@�J>���Mf h*ֶ)�����yu��}��I�!u�]�.��5]3������/n��R�[�ю~�(1�i���qZ��(~��*p� &Wx�F��
�8˯}��-թĮ:�WiTUZ�#ғ�!�#I 6�Q��4�[��Ƀ�,^�خ�D� :׎>*�ǲ��\� F�I��Y���4+i�Rc4�j?�ͺ��~!��ʍ��hK?�1Vb��r���̆^z:����oc��@̏B|�C�%˼�p��yJ��*�O�귃a&g`%�?Q��:����3r���v_&�����i�)�]\���a?z��"`=����aP�zc�Dӂ���������%����,=��;�i4lW�����Ǯ4Z۳�$ؽ�*��$��5' �x��lkNqT���h�Xf[��g� �l�u�>��lj��5�~�� Yqί��C/+{q	�� m�.E}�rl^��s�Y=��V�31��+'�!�wsO�Ж<�A��{�4�4�N�J��BD;ĸ�����&�������d!/�ALAgK����%&/�+ݠOJ����d�eL}�{���z�h�ؖ1�9Y"\�p��v�){@D���!{Y2�G+�6o�� ��������n��Z��b���%�gZ�v;�Ms�t�y&=�����2�|����|���V���>�����3�&֖%^�ø��Ҷӥ�1P�y2l6j����M!N�,_n��>���4�z��e�B�b�H�8|���$#߹p��8Z=��X§qk��2�;�hE�4,+6�}r�^����
�^_6�uP91��p'E�����$�_C�Vc�`��Z�	�(#�k���Oby�84�|4e�J���/0��ؗ��Ѷ�2�J:�c~�Scw �6�J�Aԧ�=(K�hel%g� ļk�g�)� BʨD|�Q��� ��d���ohǟ�� U���3�ٍ<eMm��]{+'�9���̚�v!����W;U.<�lxZ$b���� ���K�~��)��_7A��;�����(?Uxm�s���rX?�M.�����S�9$=0x�����bC-ܱ�n$�a^��/���;�Alo�|�g��!d= ��t�:� Ē�����?�籆!�ʬN����Xnk��/C�t�5��mC;26=�YB{-�:��m�"���7>��ZI���d��ߔl��SĴމ~_>�[�!��v4�_�B1_|#��B�QVWg��;���K{|��ǝ�|z|�A�^	�ihp &�� ���!ʷ��.�(xxb[�G:�r;鴦|yXv��Y &tl��@V��� Q��6������"�y׸;����5dڋ �=*1#QaD����K'�7ft�� F�Cm4�h��r�)����:[b��|:b�\�r����<��YbAlR�ME�����f������ �4�5%�$�4�Z4H�NS~bJjI�p���A�xt��A,�2��4��Ӗ�/��_O�چ�@�v5EM۸O��~3-:*��1&�a� -N�R����d9�<|Mqbá+<ְyti���Ĥ�Kn1� 1a�fK���:ŔE�Xo��^������a�?r��'¯�R%�w�&j�����h����P�ۯ@l��&��HU���.>��h���{��׶���q;f���iXTy��Ks��������]�q��LM>�� ��p5�z�)/��G��`:8@,Q�Jz��Q��Cw2��blB�fv�F��jr}Kd| D,M�J	bq�����ϖ���}G�E�@���m����*s]�@)�=>�v;z@箹���6�I�k�<���3�5^��\�������
b�����G"P��ݛ5��� �\��Bdn���{����r�fĄ��x�p\�H�lw���XVA�*3�B��%�� ��0p0�U�8���Q��,B7!��R�X*���P���:�m�<� �y,����,V����4GA�j�Xo7K
߽�@�;�d�wT)� ��@U]�fe�ZoU�(���9�Ġ4z�p���!T<�I�d����ؼ�q����D��3�e�����=㬪��O�rAـ�T5_i� �,��¦YPN�Ċ9�Y^�ʁ�?�ƒ������3B7ߎ��G���UDd���0����1ԫV�t�s�?�#d�*1)_�Ԗ�+$�V���b:�����:����]���[.S�{�6x��}�{����1@bp0�9.3��%FEb��ϱAL���������T8 �Z����x�JC����\X�p��lΰ@LH�]㤚�T��}���&� Ą����Y��8�!]��
�r� 1K4AN��a����f��RC���Q�9�+H_��X���T��[�o�"?�t�1���H�����?zp����kX��X�l�j<-j���m�c�ԑ5��</;��:�P��>��'/��ӰK1ӫ8��^"6�Ч���}�:���A�D�#��l����Ene�X� 6�V��]K8��x:�D��bjl����K��1)�Tw�U��I �ѳecٌg`a����|m�+�*xVK�I���;N�k����c�r�
o�kG*1�׵���T���{k}�����Β:��Q�7��m������Z�ӓ���s��beA��y���+|��jc�gF�J�xKB
�m��H�]��k�{���8?a���nq��!|�'���%���vԸ���s%^Q,�߼v��ߖ���}예��0\��ZPde�7��U1��ٛ
�c�lR��c0��d�%@�;x�pck0֪�� �Lu]��*�t9�K�:���_-K-�������$�>9*a�h���XS�]b�nSx����	e��9l:���P��9F�31�|��6/�u#}���ʔUF]Mm���U��V��Q�!����V�+�C|׼�bqԙ/�"��v�.pW�NX��AL�����'�j���"�����/ �r�(̦����a�����)�!Sq���I��A}��^نo
��U{�f:�%���;�LiCoƀث�ڕ6��i���|=�ױ� �(����Ȑ��'N��v�R_���ŵ������N3��l�-�Z&2�k�8����+.	����ԕ��{�]g'Ll��n &(�O^|L�g{[��C�5r����z�"d;����Ѕ�|�����pu
�p�=HI��9*V�8@L	�u�\D��Co�n{U����ElW)Ha%ix崻�㝲g�@l��~��yt����
���B9:��[�{�{e;��Cs�ƾ
bHፌ���d$��F=��U���*7��vH���T�_S���.^�8�7�4�6�-���C�'��Ď��WQ���EJ;��Z�P���h���h����7���q{d�-{f��d�l�[!{fWd﬷M�
!"�22#�gF���뾿�|��s��y��8��Ia�\�������;���\.� �?M�Kt�d[��'��zӜJ�k��Id*B��[���:%�,�1�նr����tLT�5�fp ��8��w��C�ly�U[�%b��<[r��E�7�P1m
��A��8�ӯ�4!~������Y�!R$����H�V��s{چH%�>@�Ѓ��Q&V�����]�����������<�H�����\B��n]�������z?5(��%�5�ׅX���'�9�
;yD��E�,�$�Y0���e���ݷ=��p ����3�#x)V��U}�����$��ɜg�K7�;z$��V�)tA���:���H2���	f�M�=�b�q���&�yk�|E��ƚ��9�X�`���,KZ13�ȫ1���y�1����m\5�9�?d)��1�Z�G���f]�b�I��: �:�˟Y#v�Q���i��A�j�,������=�G}Ҋ3}.:��5	1k�s�y�7I�Z�Խ�s����l�RE�uښtG���B��!��{f�DX��8ݷi:���e�$h�Iu���$
7��U�51���;�{?1iN�1qR��d�!��Yw�#��k�\�.j:M<W����R%���|��߿�W�������^qQ�;�c����JBL��&N\m����6�Yh!F�YKĞ���<yͧR�A��ة7��1�;��Y����;l#����#\!�H�8��u�R�\����lL�b�3����l������u���Xy���6A�]\\*�r��|�b��=�+�O����Y$��4!V�&����.�QM�9�&S��������-��;f��4μ�Y��|� f��5�e�¿�w@<}�o4W�1���-�<�S�h��h|Z�W���u{�i�/N�|,R��tN��������qr�(l.U&Q�:�j�B�S�ȸu��s�̠�������n�=��*O�Z��2�XI�ô,b͈��y�-������������5�9kR��<Lf���#��ЇX����+�����x_Ǉ��f������F�K%k>�r�1M��[���I%�w)�ڑ�.{q����$-G�`��XI���]���c�,cGr��/nUp�ɾ�Xْ���颴�R�r2m)��	bq�F��^z"�)W�Xo�c���[A�^I�0��-��=W*��y�ٗ��S��S����QG���c��~1��
dV�6�C�1UM֯���%���1�����t;�@��w��m$�aar�~|�O"#�����-��`�$Y�>(��KS�%e��U����)7�п�+7����Hܘ����u\n��7���Tt��/�35���R9�E@l�/�/]�1�*��{k[��	Ą��%����bH^孲o��@,a,�/���S/嵆Wnb��b���3�cS��	d���N���K���������.�4�b�e��
�i��a�߲ûi��9����Џ �ʋ�{�ҳx�t�b}��)�B��/=�8^�?�Ɲ!�X[�Ӄ���e����ջ
O ��Qk�C)���Q!��bQb����ww�_�ja���`�%U~����;��ҏ[�w�j;im��A��D�^^�n�3�/>�dNEz�k���z�Y��KX?��L��}�bkI�mu�i�
���bl,���S��ꐃ����1m�"u2Cv��,�����sIΖ&����1%9ƕUC��O7_Z6g���*'������+���lm�h���~��C,7qEX�u寱��`�SYł��HA�k��|[��r��M�����5���u�Dm�����J���2b�O
�����:�i����w�/B~��}�-!��XG#�f<[��ќ����~��q�W1xE�W#
�O>ي�y��p��E����ALVZ��$��q��ώ�b5,�	.�/t\)����	:�ڞ�$ֆ�㐠��恺Z��܋�����G�T��������rQ<�ҀX����?7�u���Ġ��k��0j��m=���Lmݾ�.?�����5c�_�9G�闊*k���qQ�UU6_+Hu�5���y�nh�j�1���E��#C�4+��k�B쨒�曔����Z��Lg��$����$�hVϐ�nϓxC�!�������/ߵ-��t=��b̴�ɔշѱu�#�d�v8!f���J���y���c��"Gz4�b��5��G��N{(hq7Zn�C�]w��e��*&�je�����O����ߵ���Og�>���V:��c��^g<�d�S �$�fV
i��5�����I��O\
�ZUB�Q�����۵8�������ml��|�s�r�>�M��]��[C{1G��z�bOF��ҁOk��^ �� &�S�]���n1;ǞR�<�7�K^$E�6�Gh?:�c�W���"
1i%nB=Fɦt-��Q5n�%$�i|�Ə��h�4Ǔ�^��b��l3�(6ڇ�
�v%>0%��O�B�[�V�
�Ȱ%^A~�r���F�FG|Ò�{˨,��b��(^u	�ǢGb�n^���!#p��yŻ��Y�(��5Uo[��5�t�l�)\���F��2�z�����5S^ ��ư8�M��dF [�����kQ1Z"��1��Z�B�}�|�a;v��yEq��������f����?;��~����
U���%���"W��T��>�T}���`]?�}��������M�߻�<����.��zC�=�Q"!�;C�N��(��[^C��=����t�zʉ�E�z����E�֮��6b�~�`��4��j\@���Ę�U�O���Ȇ0M<��/� &��E,V#r ya���b�y�n�˯I=�-
i9m��^�@L%�n���O�B���!��fa&q��w�l�a$ͷ0����������C�8܉m�ۂG��N��H����
0�(Д� e8F!��u�(LѢ�nU2/0���^��{c��Cц���3��L�X��Vo��e������7��Ń�F���̷��$�&�S��1�7��4VÎ��VƧGS�iV�7CW2�N
$h!����q�*ŗ��aJ�+�b�?ÿl-���z�yW��7�!I�V-%)�F�و��VJF�����b!�isu5hON�7E�L,���!�3t�%�z�Ƴ���&�F3CCb��d���Қ�侜���?	ǣ��k��N��%��̦Lj�Ī�
�?+�G�O
u�fwފǴ��n<5瓌������+>�	b�
���0g҅[1Ԣ�<&X�������B݀3e�Ʋ=U^r#�~
����נ�jEg�=���p�M�����b
E*��D8����xS�_4z�U_Z�s6� b~���P�?*3�A�Kzz�\
b1�G��!o,9)�-ͼz�'M f���4��b���*�X�?�b�X���'d�\ެk�Pc��nǅ�u �L�,��r��c���KI��!&�V���(a���:�wT�|0�M�X����6��~Rߵ�9�c�;?ǐR��/��8�K���"bU����!so������'�C̷�]�Дw��V�����T8�n�
7��R�X��1���~�A�tڛ�/���e$��O���nUAB����� ���z���&���	������ʹ���6�����g���."��ŘA� d��p�{ņCi1�+�y�V�ڿr+}H�d�z��iu�`���ZF�}�6��?=F&��G�����2#�o~	��/�P|`R��d
�N[���膺��5t⟔�Z�o�5�MYmqI�:%��V)�焘��O��.q�����K��� d`��$��V6΂���Q�r�bT����>��9_1(n~����b�tt��L)e��
yM}C�o,' F�?Yo��CN�l%�<�kA}�1e��+	���_�~tr�C,�X�q�\G<V9�%�G'��8�L����Ӱ��f�q�{S�5��K19~�5Rc'�p=L��{-�i��V���i�z�3��l�a)b��$���X��B�mk[�Q#��ѩ��p�i4���
1���5ơR��a�w�qL���Jæ٨Z%����c���-o��3
�1#���?��_�푴r�%v�!��A}vc��g�n:.Mtk=3b�����l�HR���n�sں��BľX���i�u]���c���Ob1sj�5wN�U�방>���XdX��>���ND�:����}.�M�r��]�~Q@OI���(�	��2W�N�¹*�;�u��He�}a�ڡ��ǔ�H�� 38�^
bW���B1����.dދ��$��@��:1�T��vU�e��ݳ">��]�e���g����`{8Bw�� ���U	�i��TSU[��~v��f�eY��}5,�'������F�
1'Q��H���k�7QS�hmU;Z'gI:J�(���g�n��N��+����P$�_��6���iWC,=$��޺��Λ�-�鹁��Ĥ��O�
J�����k��A��ٺYF������̂xE�Y�棪�b�]X�}��c����19�66��)���1�	��!�tA=X�}ï�uoH���B]�~~�=f�N��a�4�]%�I�|�C��'�a�\C�ÿ��Rb6*\�>���g���p�n��F�@�?@��gXB92189��*=������vD��f�OR溒	BL�Ҝ���ٗm2�Yq�E!��L��G���^�KfS�3��?bW����s?]��_9�nmA{���cT������u����M�y)���a��M�bbk�uw1i�|�ؔp��c�g*ė��f��W�$�U�ͱ��vl���7y��=�Z�X��[��.޸%Ć+O��_�!�ֻ�*��
��0�{}�C�!���Po��*%�`�uj�񣬯b�f�Gef�I�-�׭_OĽ�Xv:����S{y��Ή�H���;�����c8\Jy{�s��X�J�����W��;T�>C�d��C��p���dZ6���>���ɵ�X�և�����2�v���Yl!�x ���{���6�cªw�! b�����$��g��XմK��Sz�&��V�I.�ϛE�Q��;�	r������Ҹ?ȧ�x�~8c�%����8U
���-�5�B
Q�VAlj��&��������.J}GIߡ���b�y�oq��:b;X�s`���/�q��e$���Dc��=]}O �g���ab��|�袆���H�������o�/D�9��G�ӣ�cb^��wP��6��>e5>����|G��́�)������(㼽�B��b\�F�c?Φ��k�����b?��.�ͫV]6A�"�܁Xt����q]����1v7K� �$��U9&0ϡ��S=�r��1�wB�W��B<Yp��W�6D�� ���-�ֻnG��k������@ĸ	O���������@&1xTA��/��{��fq]>�]��Yy�^�eh��7�Jo'&�܃����dmd'��v��z��
�Ia��wg�Gh���ePh� `$�i��S�.��n�Ni$E�;�>4ȡC�FB$�3�3��~w߿�<�D�b�Eɗ��M�.�izLa'�*�I|�V0�ǻ�i~k��f��h(N,�^)�

�|Xb�X^���=�+�p"��)
��y��t���xȴ@�6��U�ʲ�ݧ��x���KG�P��N����zQ�gWF+9%�0y�*; �+�+�J��N(�4�p�t
%���� ����F���<�l�� �}��7�n���ċ=�o�s�?bd��;�N�8��%����5�o����ݠp
)�G��L�[|����d3T�B�X%��Wv��b|R'�l.c*������-6[ v�y.?�Q���#u*;�u9p��{ס8�Ϲ���a�j����o �7L��L�H��v8�B &�=�gc�6)�1/<e�]�*��O�^� r�|�*D��X�X1tդ�a�z����i�GTJ�-�Q80��τ�2��ذC�,�s�]�u<�d�v�}�Ƽ瘘��j�<y��^��J��C_%C�3���������I�Ŧک�	��'�k��֭_d�
����w�X�d���[t\})�����,�h9#~�򺍍��O��QaR{�G�IS�ci�M]�H�)`o���U1�zB�o��|{'>�ȵMĈ� �ދ��ZV??ϓ^z���(����Ҵ"�h���@9�A,��L��s���JmuW�\ �e&n�[aQg���{�G����J���!uQ���N�
[���|x��/�&^��h���2�}BN�V3�N+R�˒�%GV�B�@�I��#S]6'Y,�j@���A�:���J+]���J�Źj�����K1O�t'�����.Ź�B3n�HwJ�7'���xFĊ~�M!M5���	>��z)�3�J�9<�� �1ݮ����8N�ƛ��	u�� FZ{@�5Զ]�*7qP��u%P�b#�1f�Ե��/nR��&� �j���l����	]��K��e;��3�t�f4dJ�?/��*>���E��>]Qxvm��-1�����[�TkN��VF[v�+���1��w)O#��c�=WT��/����A��žLOܰ�:T��ËИ`{~�f�ͼ�́�(�ʈ��%���9�<9�>��Z��Y�p�;� by%��O�J�d�Qy$�r@��Tu�U�خS�D�$��C(%�aɦ@6�8�H���g%K��� �W����fU_Bvf(�2�������<�k�=Y�
\�d��=� V�_��A��n��>��������eu��#���8�ßOǀ���9Զ}_�����ސ<�b&��f���a&�����Z�ط�$�OcV�2FK0s�L��5AlF
?��7���t�@�3dC�)m�Y23ඎ�7(�U�{���.Č��:�)�����N{=2�� �LʝM-�"
��%���8V���~ʇ��]e�4�� �� �.�����2��&�V[��P9Xch�����./�ŕ��;�Û4K�]fH�L�`�@f�;M��&��>۷yU�~�X�a��*����a��~�*���91�g@W�N�-�9���TO�l�_:wun�Ͷ�x_Ğ-z�c�W4|�ڭ��#JP�g�1N��+���M�Y_��S�����}����v�?�el�-�b�R����Pp`��9�KI�= 1�p���3pcc̚",�k�� ��1��z��z[�6L�ש-�$��]P�K#��Gۉ\��r���`#�Kl*���~+F!C�K��X�3B��okF2}ܵ�
bl^r�&A�:�?��K�v����vd�܊��U��qS�i˿!������n���d��.1%Dv�f]�U"�^f<���^S�>@m!'�����4#��CU�bŭ��aNn���?��ߨ�@�`��y��({1��ᡪy���[�9�QL$1���
:��vpv�?J ��
���
��T�o��t���c��_�y��dn���
߿
���F����*�j$o��Q�Ǳ��ks����ף����p͗S��JĲf	�ȕY�f��H䇫�Ը���sD7'�çl4�ف�p�" Vׄ����^���a�B�R�{��{�AIi��C�62��w��IyM������%�:A\�oFw�ɐ鏛�6��*��%��S���clK�ށ~�"Y5Fݼ� ��k�LEuR��g�%��$���-���矒�e�8P}���;n�b\ظ��rFv݋g8yh.L_�AL_RE���������6G���� I.-&���/]㙎��)�9c�7#�Ú�׾\G^S��r��o��0�c�Y��׻yD�K�DuɚZ�;��б����=������(l����JϨ@���a򁰙݂�.���	ڹ=
�}#��,]�5V���h�É�@��$.������x����,�{ �(����f�-���Ј��u1��]���`�x<c&�f��G#��^���LX�.�c��o���S\@�!L#�CeL�n�;bU�O*�[M!�,S=�ڭ�@��}������f�Q���۠���8!~qqT���23m�O`-��G�=�l��ZI�q���>����	�n��:,6B*����aY��?=4�˦X�hd�&�����wS��~(�����%�R�پ�%��q� 6��Ƿ5�Xb)51��c���2��tV徙�x�Y�FP���zb%-�9Uz�4{�o�C�>�l�e�w�?��o&�v��*��!ݭ|CVHGH��E&�r����&M��.�v�jEb�Ѝ�5_�94U���4Ͷ�1�sH�9��F�oo��,�0�I�j�ħj(Ŋj�1�Q_���A`X�7��}����6� ˷� F�$/�k�?���𭴙�5�	.����>U�;��N�i���Y�
b1�.����9ջL��V��� V��k�n)`��l*�	=%�������C�e|wj����!���� ���B�(d_�x�(:�򶬃6+ �ؼ&���h���}#��Ƨ�·�0�^)۾��� �A�'O\n,��8��3^�78�tSo)���hWU����؁����y՚R�Hw�|����Mz绉u%�ЙS�cG�Ds��j�l�H~�U�XTԿ����N6���]�w^n�;����~�,��m�IF��r��ѫL��4߿2�"*�WS�c�jz�ߵ�ˎ�V�V�@�ꛚZ�4]��c�� �ʆ9�#����֑�mx0�R�?��ͪ�^oJެ��z�i��6ꃘuA��7[��w�"�["=
_u
 �� A�" ��c�4��6�����b�\�᨜{�ۛ�*��X�����3�FqG��{b�BG�ALY�0�M��M� ���s��7�5 fyXOod��p���6����'��Y�/;��^:C�8a�w�B�I6g��>�I�k��e�֥���l��m&�X<S�	m���.��@w���N+SL�R�2��1��~�:�e&� ���ڲ������8��r����c��'�U%�&i	����P>*����:������@%� 'M �b��{�Љ7sy��B���_nA�#hL���gT�C��IV��8�ډ?���v3oFW�`N���U��NO�z�ZX���Ix~�*�/��N�2�t��5��v!������|�_L�o��o��i1�i�zRm�Y6_Q1��؋�m��2�U�p�C���)��NB�"��&$�ű�iӠ�8G���4�W'�6(���{E�A�������{���� ��H�=�����T)f�:j���$ă�x�k�]�&���hɧDp1�������-��YNa�.��y2O}Ҫק�����:^��s�㳸�����:�0x;�{�;>�z��'|�u��z �x#�����$6�߀�:^�bDV3�zeܪ´�x
W%��r�v���E���W/����dAl���Q���ӫ�����N���l �y��Z�j���]h��`/}!�%�Gh��/A�S}�IK	��p��i"w�?��_JM��j�l.�j����b��sh
�*-7G�
�� F)��w;$�ז��W��;�:Oa��3$sQn;���w��ASC~U�)�d��� Rk��[�b�VQ�ݴ��9�>!:.l?ʽ@̖�E�"?���g ?<�
>�<������y`8�`K��rowX���˾��|�c��dQ[��ݟ	��sK &�fϮ�|�J�hw���,�Lh'�Q�d�`�r�ٺ; ���CS1b�k?w*F�tj���j�8����;IJ�|"m��g[n��b��_���Q�@Z�tI]�q��f�߳E��l���� O�k���:uf�+�t�\�{���GɅɧb�o��''Pb��R��h�"�j��
˞x�% f���l�������\���Q�����:i�{�!�3�M��H �B�(�8|����'pn��\2����������^��rz�����X����}�>�u�9�������#�
�,;���~V��rڼ�4bJ����}XO/k��T���Ќ@,��!���g��C���{��-S�8�b�wל���lEz�]���1��J�+>�Y�2͖���g g�9��Irj�!xGg��@7b��X����T�yb��͕A�ʵ;���%�sx��Q�̦��?Fp���4�]��w�y�6�~�q����w�U�E�!�n~�Wn��OAL�,�� N<���#�*�y1�R ���:҉������@��܀ZD���Y.nRqcI	T�=��u
�����)n�ę�I�p��!����1b��[��r�BX�x��z�[�ov���F\�$v��UF&x2Nzr���@�D^m!u�3I��V�UT��텝*L�h�E��� [a(n 1�A���qZAG��YX���Uu4 V�Ĝ���Y���Fjp��;ܮ��-��4&�zK��gr�#���1x��띢n��R����8>%��'|����%ak�˿�Ԋ����ܾ!��y�	���w(�B�A���K�H�y��l��#�P�Qc��;���I��6�4�T���i���p��Af��:2���xɋ���-'6Sfc�֊�4]c�4�h+�Fa �n��`'�Zw��_�LD㮟Y��n~_���va[C���	�����<�I�M]�za|��V��$z"���bT-���0�)����-�ZR��a��_v��=��L����u`�	��$-�I��,�^��~<�9U?�He����zc�B3���y$�Wx��Q��U�o�|�ո[�4���5��C�x(���Ubj
DGCt�dI����_	�������=_���4S�I4$Ś��ە���7�K˨�Z.�?5"N23cd,�n"X��)	;`�)O0�*4�MT��"�����9��移iF�[Z]�b�aW��j��T'�V,���ʯ���;�7�|�ҞN�\a����Ǘ�m�ib����ܙf*��ʗ���E�C� f'�a�Ȓ):� �B�#�1�j�m��ZZ��D���b�:�X�t�����ǳ��p�#]2�7 ���Q�z�hDl?�%�U���E=b���Q&��Ӥh��Mu��J��2�y�ЉC�f��T�tj!b�[4+u�5�*��ێ
��/�2~b��;�~h���eS�aa��Jw����KR�n���Ewww#�-H�t�t���lg��q�{����?�T_m��4�#�Z���7�h �[�����A��E�:Q�&��I�{7 ����� 
��-�n�4y���!�I]��"�7��ȆmC�>���d���f`
JD�8��լ�ǅ����+�N�N*_�mp�-`8���� ��Kiv!D�a�(�����;�0Ov�m`��ҋޗ	���^��Y� 1��H+"�r'�ϝ𻔸,���DA,�0d������?�J*_��1��:�ͧS�w�qGW�)�=1h�5V9�a���n�ͮ��=��}�i��*I�1���A�#)�Ķ
~�&Ju���|O�'4�1��2'�	�j4�/��ʘ�* ��"S����\ϲ�K�t҂�Vڐ	[(BԈ<Yo�Zi�G�m~,<�)�K����4A�3�! � �V��,Pkh��45�wc�b~�t𐱥�rM[���z߀X%���Y2"e�fY>��Fk������7m\2��e��Ա��YVF-P�����Yi!�@ܶ�1+��p{�p�7K��o_8�߃�![�h��WV91Iv�w��� F��ǡ+%&[,G�8�Ɗb��)"n���-��	uN؏�#/Ay��&$�;��48I^}����킥E�������ėNmV@,�h��Ru@]��;{�H������f��;��4=)�@	7�4�ĮݗO���4}�,r'�<� f���е�䨏�� ��]X�����_��@ZI��7��K�b�����؁w�1�r��ź���q��XR�G�U�*s9�N�u����A�1�}$��J�z��Xοy�����%��i$">�"D��E���XQt�oê���=�"��3IFf"�Ȟ�P��_�8��:����/��~�E�]�D끦��Π�N�E��@��]K(�:�y��ё�����a�[��o�34lE�;Z1�A�ShՈ{w�����b_{�s��4:�e}J��b�&1�]��;G��9;��zJ����%�ˆRw��}ǲS�Se�=���_��/+�b=�@D�c(Z�� >/�,�i�0���(�W�ܔ�fN�9Fi��H���U��D���P#�o)���P�n��	��h�+im�GXԕ�n*(�|�*?�,?T���q�;�N��4��>�z�L�: ��0��.�����1�C%g�������ώ��%�Y3鶆)�w��&o�	�	z�u����f4S��d����:T	ĪX�rS,�?�:��7���"�H����� �N��#����*��	ڇ �!�l Q@��N9J��{ytb�q��b�T»�y��m~�l�X �Y����vn���R�b�'jF|�A�����>��ٝ ����Lt���rGm�����Ci���T((�C�D
�Jv�G8gG@l����WG%�������Z@Db�w��T�hjw�n�Q�K�)� 6��PJ`U���J6dj~�ub�l)1�ʗ2��"q�x%@�w���N��G��4���*�0��Gv;2)m��a
l�����	]��z�Hd��Uv�)�5�5ҡ��O�5�$�2Q�ܮ�-� v�R_s�W=�O�:	O����ۚ�:� �70����ab��z�=E������S�,Z F�'�W�����E��;A%�]b+���Pn�>���웶
)
ic+�{�m_�2GU?s#��=� b=�&a$�{��u��X��Y���+����ğm	��TOl��j�TAl�٘߹!Eq3�3yx�M�ĸ�;�i����4,��[�;�X!/�I�����Q��ӣ�g�1 ��v���[�5r&-W��%Ĥ��KX�0'��۶�>1��֑��f�C�x��U,��{I��8�P�M͂q�q���~ca��Hb9
��-�o�g���CfN�@����E6|��hx`l���)ǈ�/�k8�
��evs�������b}��4O����������-a�9���~�Aw��[��j�NED0�>�+����h�&pI,��ʘ���6��'I�e��������AS�)x�y���������i�S�x���n�Я;V�=��=Ķ��+\..��k��hm�����G�t
����rA��O��;�rW�ݰ'�ef���9ZS� V�L�@Khok#��cZ� �} �nHJ�^(�s҇�s�dy��q7�X��ӣCq���7^�߬��v��@,�������ྜ��>�5WZ�@��}r6;]����h�JV�~���!N��B79v��Sd����S ��{7&�HM�g��,P$����^��j��0��=]A������>��*;
���㮋����׏A�]�^�Õ��EةC�����(.��}�0h�X�QڴR��D��A1_�^����5�K��;��$+�_��F���f� Gs&@bc�oM��˴R.�X�Ǯ���Q@wyqc-�>Qz�&�<�'u��f	�{?3V�E�R�ޣ��U���ةvDM���[���c^���k�!�<X6�b�|�E���Jb�TD�b�gE�y2'KІti�x�񚎯 ���ȴTJ��od7�`�?��1g�4]׆���!��ȶak��/ Ƭ�>ԭ?��-yc�kܾ�1��xw�����'ԡ��5�}%�1�f��G
<{y��:y�)b�+�2�iI�*-ԕ�?��Wb��Z�*_�q���7���{��ZbG f�O�9�=�cKo'��^�H�
�UU��Dh����KϺ�'���c7����;�Q7��^�w�) ��T�ź��J�&�_�<S�*Č�o��d��9�N�R�h�XI�0S��}!��{�gfX�kc�T����Db�}.zo�Z�`b]C�:�r�1\�J���_hI9K��n�_���;x�%�8SG��^�!W4��^c�����N�Ĳv�$�N�G�*
P��mrA�>_��%,���=;��iI^�xF^�TX�6]��]����� �}��S&ƨ-�$n���Z}n 6Jj�A)h���d�������e�,n�:�����f*�B
�3@�Y�i/��"���>�6���b��>�7��s��(SS�0�|����
��u"C��ʮ�O6�u,&Y�V�G%��B�1�J�J_��F�Y˕ၩ�s�_!��{p�� �oRĀ���t]A������������<����`�}5���E	b>��	�a��u.FF��1(, &&mP�xQ�������8�ז��曾�U��u��lY�����1l�{�INr�FW|��ot��2@L�Ԏm�+3Fz�v\�S�,����3�M���]�l��{�O@̼X^e�?���A�+K��6�h���*����ǆp9<v�(4�ʆA��۝8Yr*��!<�"'Ą/?.�Tz�$x[=��}g�����Ӥ��K�@/��&�&*�@�9��ǧ*�R��B��y��,�Ѧk�W���j�8��m��}�b��V�2�n�=R/e^fI����1_yx����K��ʕO��x�-C��zo6���RAGAz����l���Q���eH�h#�N�A�EvS׈�������a#�V��%�;�xGj?�r�b�O%Ŀ��b�#�ʚ�y=���K�g�wG�P��y���`}���#��/�;t��� �~� �>�܋us9�Y��`	bt3���],�.]���z�Hi���ϙwA�wO�X�U5�=��e@��8�ߥ
6��y��<&��s��Ĝ��(`d��9j���T(�k��˿��:�XsT"�y�{#�N4+bfd��;��.�|��#�H9A,��$-���X"��7����wF�7������MF�������F����O�|b��sA1����]�u���{�_"�Z\q ����|�>�����|"J`�1q�5v�M٥���M�+����歈\����3Ie���z�Pꀘ8�h������5B}��F�#!5	�{���n�#��"�"�I�]��(b���TT]������nfh�A��G(��Iҹ�K�u�.ȣ�T Ɖ(���6N)�m�_���=F1�W����<��ގ0�Ac��N@�.3)�s�~SW7'�ASZ���b�1��>��Tɣ���Nq�f��kA�C��c�Y3�uy*��	7���5])�b�j���x�7�	�|�k5qy����
Y����,Alәwp�sj����R%7F�kn����f��s7I���!���1>V���i��e�Ԟ���RL�%ZTh���2�LdNW��v�̦�X�D�xa�0�St��,��I���9 ��%�D'�É+n����P$�������g����W����{ ���q0��;9�3�=���Ý��4���$��
+o���ZA,�s/3�Ј��#X�1��ė�,�!�jݦkt����Xu�<P���+�R����/�ׁ�p�$��UA�mo�3GB�Z��p�L��� CI�ߌ���3��<�+_`����~# ��ĚG4e2	Wޘ�D�O=c	�Z���]��j������F��&[#�W��f�g@Y��>�j�O�^�A��*��9z��Rx�_�XQh{���ݓ���0�����<� �a����%��S̑^�P����:�`��}��8ciXПV����h:�4:�������-����N�)e�T��=�69% b�\����|\?��V�!���~�	l-�9�R��'��`�N �c&-�M����O�����&ں��@l�[	M���Zk/�{���`
�ʒC]c�E�@�;�:&�i��ߝ��+y�;e4q��ݏA�T�����ls�����֏�0���3@�b����=�3� a&��wOni���������䍃�M��$�@�DS�U|5I��5ӡ�F�b�>e��u#��Q��Nc���X�@B��Rr�̜��1�%_�^�o+������s�מfz'�p+�6U���9�Ð�c��~��!R|ko3dsNp�$~}j�D=�
H��#^.��ʌQ�X��}͕^Y�m����5C��m�f�mpN�%�����{٘�4��6�f�)y���jALpo^�F���y�l3'�eǷ{L���~�:bU�?��y���O����'�}N�R-y�<u���y��%�����E/��f��u�+�j�X�,}*4�^n�0�L�i�(i��<h��Wx�Orr���3A���R�C�v�UŋL;�Nް�f�l��h�B�o��|�q6r@�?�;�,S� 8�����d���&�/���ǚ`�p��r��KХOֆSk�
�X�呃U;31�)5�OH8=$�Ĳa����,�&8(
���^� f���G_�>y�q�΂�dnbW�%�{��H��Cg��aQ�� �z��kM�3�p�Z��� F2ݶ̟��_:���o)3Z�i�.�9[���ki���`��n9��h#�;�<��OG=1��֬N}�m��#}p1�/���@��!E�qe���>bp=��3�)���5t���U�K��\����L�Q���Ci�|%��eT�����?���MM`P��O��C���;�C��/���?�^Th���eP�� `���A:�$���[iq�;vii�naA���[��sf�q�w�����E��P�g�w"�;���������N�asI8����E'��j����D��Q�E��ʐV>&oz33bF����p�Z.��e>�݆F��؊��֐�9�1-�������a����o}Fۄ�s �c$#R��Y���y������,� tN��sĉ=�c 6{q�q¾_�/�:1�q�^����������?a<��B<v�2zw�7^�b�'��t>�����m9Fo�Y1֝Ү��=Y�����Y>b��f�1��El��	��	� ����CS��߃l��)�g�:q�V~7�?�?Ϗ��B��NA;��-�fm�"�W�߹�  u�[R�|~8�Y35�o6��Q�fZ��[���W��XM�oj�Hr@L�
.�O)���e"�m��|�b��P�����X&�!��Wc�������������>�x�Z��v ֥���
/�41�R2���ab�$u���58]���)���� �������4��2���K7�ˬhį�������y#l�]�w`k2l���!�}
��z�,q�Rs̨|ߒ�����b��Y��{�hk�fu��/����s�ˆ�2Db�J������\�K��A�i�g}�ґ5�hhs�}��zZ���U�?6�m�����Ŝ��ȕ��g5�A�֋�l��P4?s1b �����~1�ya0���o�&���B���� �}�ۀ�0���2٬M���bC���n�"�r�����<���XLl�K��(?g2|��x�Jd���^��yiH�j��-��DM���)�n�%�|�628y@lɶ��4����d!N�a�[��p��`z�֗��a.ɨ����c�e�<� ��M����ĄL
����~a� �LxT�%40vFdT�����ق@L�J-O�4�.����c�Փ<h �aA���(H��u��&�]����b$����~�k~Z��m�@���^��ev��(�"��k�TY�2�G]�]�ye��hؔ��V�r�V���Z��'���'�Q�D��|�-#�F.��	��z]F{8������Q �Sꤌ�fժ�� v�\y�~��pA�ę��
{�S�Z�)h4_$�	5q����Em1�j���������[��0��z0�LP�-������%���@����7�]�R�Tl��e!gۖ1���T��J!c�����1���r����f-lR��]��(OʦM8���]�L����Ħȏ�8��P��E�F#Y�����;�f�2�Rwn�H���?���x�{ZR���d��������t7�l����tчX	�6Dh��1�U�!k�����41�z���΁�S�%!䶉 ��|M��:{�,co8F}����i���B�c���� �m1p���kQUA�u�H�,w1�0	�;�	��D�HZ��@�"G�=ܺ3�98�!��b��3j�� �Ba�U�]�s;���4[�1�1^��j|�>jP1����p������!#hR�s�$�4r� m� ����f��b��1��2���ꬺ�|���SIcCf�#^�<.C���95�	�9y↲����U�{D݋�1A��yui�a!	�ȼ�y���2��h �4���s��x�O�9����G�����D'�/�����} b�n;�{{��h?���'^߀غ����X�����ER:A�{2�MV���b�������u�}
��� ��S��%{_`N,�ī &�w����Gj7anjnY��+K�gnѳ�J9ˣ��R��;����u�!G�y�D����<�V;�8w�	�J��N݌l����������m���"�]
]�<����K{E��Lɺ�X:�0ףh_��P���/���~}W��s\jO������W��K�$��� ����BoGU ��I�û�<Ħ�l��K�`o�>��N�#B���@�R� ;�M?�&/iV:�	bj1�����?b��xT��@l8=�����@1ڕ)�%�1��AB���*�L��k7u�(Gڿ-����e;�}��B�d�P8=�h�S�b;�Dߥ�hh�*���5۪����CnL�9����!��'�� �W�,l��?�J��
�|/;bR4��JK�j�Z_^F$���=�1��te�
��I�g�W} w.^��=oOe�ĦT��?��ǔ����L����i��g��D5"2�m�w�C-�	{�<��B�����sU�f�XA���iֹ�������{{�U� vh� ˻P�B�"8ɪ�A�J� c��c�YRR�IE���Ěr�%!$�g/C^$h��e�u-1������Mk�Y�Pf�V�yO@�ɱ�*z�6�6�a��J+�	b)���)��N�luCdC�+�Q@��z'�J^�t^���b�k�Z+���zk;d͐�u���ח��]q1���[�K�҅O��-�AL9���x�xc~|���mT���������[������V��h���m��Fi(+G�񲞮���N.��AN� �ad��4��,z�)Cb�ϚW=��������o���E��6�	<s7+�JZ�81�@���tksV`m�Opb	�m�����K����b�����(#r� ��%nsD(Ì�J���6L!o�����n#��^�Ar<���	��1/&ؼ���ؑ;M��'�M�U��oO*���-G/;�w3����a
�g;�_��H>a��1�0~�#�H+�)�NM�jtֆ-�0Pzf��W�oU� �2���XV;Ut�:�Ǐ�_���U@�ˠܰ�h�%O��>ňLA�
�A��s�!�� :�s�9����-�H�o��
q��>��gҾS� �92�R�<��Z*�g���������({�O�}`x)���Ć7���%\�7A+��o��.@���#ŝX�x�d�=d*n�Cq�^If#f�����Br~b�98��L\�ִ
M����Ĕ��ƪ���v�s���Z��7
�X�u���n���ۥ���lY��U$H����SGo5��E8��lU`�U��<����WX��Ģ�Uh�g��.�F��[r���DE[+���7��V��J�oP(�I�>�y
A�A�����?��b����nEJ�{�t�=�vgc�4���Q0�ț.��
ɲNT<�����s��]l�<�[�O�x9>��oAl����1�ҧ�����u᷆�X�6������0}�>$�4'E�*|z�����T�Ҿ~�ڋbrx�gD�x|W+�Wz��z� 6 ��r�tɟ^�7-G�E�x2b�!F��#_F(+��v�o�	���ɶJ�T���-���t�X��1_'Ӿ��^�x�A�P1�I�R7XFʲ<���^w�2L�u6?��F��
���tc.�3���~2���s���d�0Q�pxe�B��J�}�Q�'(`���� ���GX�&�O�%��l�S[��������!�%'nM��x�b�޶�\y�s|Y��oH��	��d���Yr�g��	C�m3<��� f��f��l��g��]���O݃r�A���qh�I����	��^�o�ֻ��=ҭ'	�K2�3��ٰ�����>����Ah��y��c7��Ѣ�f0g����?��W�Ŧb��u=������#��V����_����FC��Z�L_��E�q_�	�!�2?�<��~�ї��KI��uSb���X*�.�V'�0
lA�.b��������R����ݑ�eA̠<L�ck�UK��-�!��P��Ģ�����+V�\@fWS'AL�"1�Y��/$���\;�x���{�H+��}Gl�y̯�M�& &b�=�(1��rΚ�e�R��5Ďq����-e�Ŷ1GةA��@��H}#�h�\˖���D�ZO
�r������!�S,�\�����&��Y��)Z�[:]e����X 1t7D�h��Z\�U��d"��@���Ërޓ���|J�d���VĀ���������ŝOg�˅@L��v�6Ks�>��Y�GQQ���xb�)���WW
Ƣ�|��RNb�b4>;P�LS&�����0JSW{���y���AX�F%{��� Vg�"�]E���Y�������)qr�����ܿ%xq�;?����1q3����v�o��<_�h�1��k͒��Kh[NG��=�=��@,�ԼIy�;5���&�ɰ|�3S}��\�~�)�~�k"�C�b�3s�Vؗ��A
m����B| 6�}DO\;���R���1�U�]�O���R��"��A�ŽS��G��:0�E��ި�s�?s�@,�x�@�[n$��b�lk/�)
Ă��3��Y1&QQF[�]}$�߅����H'i6W�Y/̂�v�3��7֡�>�&��~�j��u�g%Y
bbD$o��V9.�G%&$�BL�A*XK=�@Q��5l�Rz2�\�b����Ȗ	�6�,�p��30�%�c�o��mv�>U�q?������(n�|��j�j���E��ː�3jFϛuK�6I���G�����K/H�W}Kb���m��25 V��έ�^#gO�y�b�����|kg���`�~g4��u�G1�"rl-�1e�C���$�~(�X�g^/v`����$a����7= 1�}�P%+�K� �!��eEzӬ�=�Ö�ʹ�kLk�5���1��D��ܓ��j�Y�X�Q|� 6e��z�c��~]�@?�xi	bW*r�l���Q�B��"XP��1���[���$���dI�<V� -�`|;ԓ1��$�q*b���9/Ͱn$3H��K��@81���k����=4��}��b���&�^Z�՘���ݸ������m��T��=�
L��|�U�����rۧӏ['������rd��H*Ɣ�n��v�Ps-�1ԼzF~�q�[ScsJ�L��	b��FH�&n�1H��if���u�ꚦ��^�����^b;���@,�����ɋ�h),e���]b�>��]l�VʟF��ľ�nǻ�b��,�}���"�iWߥ�����~�NVθ�ZJ�����%�,�㮶#���(�@1G5*3j�b�#T�c��_z��,�K�_F�X�C2]��t��2��-Y��A ������_,U)U�@���+�b�Б��[]�1u��]m�� FqSO�͠]�d��`O��C�L%b�乱����켞���d�0���O�{�`��y��g���,r�1�f>7��ńZ�9CY�1273�3�NI���Ḋ�`�g�Kb}XM��t�J-Rs���Ez�u�Al�gU"2Qյ@�Z,!�~���a�������O�?Ԅ�����A,�^梱h�������IEH�k[���O�u/A8����0u�u�ib=J����a��R��=�	vC@,d��W�p�wl�H�����U����L����a>��H�fj����wØH����H)oūcI@l�f��������~����� ��_��R[��IVS������
��߶^��c)*�"
��8�|bW�W��u�B5˨|?-MK�I���!vg������'����l�:� �{�5@h���eX� `��A�;��ip(�AZ@@��K@�$������Ki%w���sC�����2��\��5W*z-�TL;�`b'Z?l�4�{���~�� �����4�|����愴 ���j�^%�l�'�t�8�lp��X�DzX,g2�����4Xą� �}��F8���;H��qx
���>j�ԁ')�aZ��ɪ�~S���%1��ʧ;�O�O�h�ъ��Vi@��i�ӓ��ˤ���t�:&�;�=�������2ΔWs�M�S��>����w� ֏u�Y�X˷�ܡ�{��S�Ix�Jwŭbۮ�!kA}��O�M��r\N 6��,[�4�f�<��lG8�)n0�3y�d����%�m�%��;́X��
rƥ��ޔV��ˈ� ��WW��F�ߌނvZu�m���ʚ,��o��1��u���������@�H
S/��媯 ����%z��n��:���8mĨ�[:�Yk������i|�1E��7��x�Dd�hO�^�0炘rԀgÓ8�Y�l�'�,;d��� V�qM:�d�@��C�|�<.v$b��-�խ���XW�$h��1 &���MNq�����Qs	�^��KK�|�v�%l����$=h��f{���p�'Lc�m�*����]���)��#kJ�9�X֢ � '�U�QZ��`�{u5.��RĄ"ᰫ��&0�GCF21KXwA���V�dV	TBEhH|X-��~���v�b�qh}����u�|�~b�=h2!��JF�jf���@�O	��u���n�O���,*����CTU������2����k��v~*P�a�i<OQ�|4���({�7e��,�Ɛp�������5{w,D�u^Ѷvw�(!��?=g��r��A;h*��k������5� 湁@��C�z�N�IZ���b�zk��!����V+|1J V}{u���6��4d0��2�6b�FGu����X�cY��,�Ӵ~p� �G������G��\,P	b��\9Q-9�QK:��1/|5z@,�B��{G 
$��~|����6CЬJiMY��-?uM+�0c~h^ bq�:�//�5��uy��T�j@̩�i�]p�ݨ�W^��Ї(r �9���j�������P��33��=$�p�����=�~_��hb� "��cH�O�'�ל�%X��Nj�e��Ff��yC?��$�v{[��7΄����2�Ek:���Rt���8�Q�!�1�l�ܚb�bZ��A���*�ٱ$.�� ���qԕo�@���\ZX1M�����b[n鍧H
d� ��g��(B��8|���v<���7t6��9~
�~���}*<�
b]z�����vv��Ƈ%}Z�O@�&�&�;4����cF�&T����b�2ɕgVU��;3$ ���xQ^�W��Q~��\��i~��oۓ��otI���(�5"�9FP�_��wc��(mRF���`A�s&:�k[5@��r�M�~�Nt���7K��|#�!/��h�,R9�������
bN�J�dJ���u��R��lrA�6��|�$Ԏ�(yQ�%8#� �P+�Xr�����j<�/P�U3�CAL2T�;l�TO~���H�+A�&�����.7g����g�d>�����L�Y�|M�3=ו4�xI$�2t�ٗ���ߗ�D#*�YNQK�zC��Gġ8,�C��C��B�Ϙ~�h8��mCa*{�E���>����{��iG��k��~�Ќ4�o&,I���k�e��6���wY�w��8��m�d��i��=�oP_;�;ǡhB=�c��P�s��X�ڬpA�򣿵�V�?�����O#��g>�v���'�D����a|�}	��U���X�\�����G�W?��/���.{�g��@��D{oJ�X� ���3~��?MrԶN���4�I?�7�$\������x�o��ل�sa�=���-
E�z��"7(wo�r�M���b�����`���B{9=o����F�a�����3$�p���űޯ�E�v7�a� 6��{�6լ���0WR��Z�]{� {�]R�r5�Q�B�a3��J�F� 9,N��2��?�m��O`����Q�TĚ�A���򈸯���D�8���*&�=��P�4�'����&\g�a�^ Ʃ�7I�y t�O�O�cX<�b1�O�c�y;����\$P����@�	����8w)���P�n(�B���-x��171-�k��b��~�S���$b<M����
HۼL�yny쨍q��[M�5�a�U6���>O��9Č$�I���g�B�&\�����p�a5��_�s�WO���G���B�vؖ=��b�UN"[q�+z�g՞01������J_���-B��yO^��ɏ�K+{�K��-~��ʯZJ�2@�nvN�&��ַ�75���U��� ƷvGMhp,<c���=a1.FLz*srX���eNv������p���5�_�.	�k1;K_��y�����Q�{bg2A6�"���>9���a<�LQ�bĒQ6��D�.7Ͳ2���&� F�F(��蚁(=�ά�ЫH�	b���-r��{�{�(��V?�1���%|��|�8ND��I ��}�q�f��F�yw��C�/�ԏ�����Ϫl��ݺR;���ԯ�����f�pwTէm\�UVh.��ڀ؋��,��jͪY�r(&u��� ���Z�F��@��ݲ�֗��o���V�ztמXhvϻG�Cf�1I��Ĝu����XY�"�!�,l~�-���zףd9}c����-ɧ
�T����_��Ve���y'�W�����bϗ([y��M��E6�)�%{Dj�n��T��
�c9
��f��x����·G�x�Q?�HA���p�=Rē/nc�4ㇹF� �h���'��H��t��%n��)Qd2bm�%Kh��.ݐN�qc!����s촵�s/K�f�x�b��V\Ik�n��ܘޯ)�/LH@��ַ��ɯ�DĬ����t�ľ5��e%�-��c�Wv@^��,��������3B���Bp�T"t���c�[.8TR��W.�l]����*���Ͼv�X�:%�ҩi�:A,�V�B��]R�[��&�b4k�LO��vZY��[�v���1�̇D���sST�Ǥ-�_%�!��X� Ƒ�@M���5%L/߉���+���sI��~��_�2�H�1�A˙dL-S���rg92�i?�ɵ�J^9���s��xQd���:�ub��s��2=�|a`��j�����>��pwu.��$��b̬���#�Ufg?�~h��2���P"�6�[��;�^�W�� �� ���p2�Cٖ�:��&������ǋ0Zͺ3��1��rd;6����V�8��5�|s��Y�:��Qh����D�7
��-�'u\��Y��B�'0��%�@�ZZ:3�{ߏvAچ�s�y ��z�+u�u^���Fz"��X�-+��&c��'dY_%Y[	Ć���8T?�q�&JF��e�s1ϯ�ꋯ݈nF��Q(�@�pQg�w������z�;Gg� V<&O "��0{�m 4����b\_ʅ�іS����ŭs��F�AL��gB��ᷧ��!���gP󻤒*w�Bk<�ź���4�� b%�e�JZ߲��X�v�ۘ�U��M*ZEQd�U}]�2,�K��1��a����d��#t)� �7���<$b��P��r�T56be�'HT�%^���!���un� ff-��a\�N�j����rw�-�V�ZN#Jk�堂)ҖƼ�(� f�Z� �;�����E;!��Y��-�\x睐��;M[��~Ȇ�z�G����7j�� �vHI2"��x��}/-F^���!����3X�r}0�����3��ݮי�Yj|�n6zVL|ki�6�Qh�(�%�j�n��/b��%��K��|�K��pC��E׮(@l�ǆ"��bo.J���m/���������5@$L<"��hZ�Al\h�,Ğ��٦q������󛗦J������t!E�Y�1�-$*|J?$y�I$�� &t�r�b�|��*���aiW���E�{���$�"L2�9}��Z� a���T�w>�� �+���o��7*�F�|��0j��;�f� �0V% ֿ�ba�)ރ��{
b��w�zq�4INxއb6�����R)en�e��nK���u��z��6��4�<IR�M1���a݋�m��
n-���(�k��";"SY�J��u'�� b��EQĚ=u���aضԒ� FC�`] �`�d��8q�Ν��b�	���>,���sf���� �^G������Lk 3^����`���Q���dS�hE�}y���]��Yd$�x5fS�����4(2��!�$D�!���-W�%ʓp�&	��%�%|�DH�����Wa|x�ō�a�Fo�(;�]�Z�s����}���pʫ���P�ͲE�0���>m=�T*1��6��:�[�G����Ⱦ��@́�q(��l	��ndy~�=?��|����#�Мڍ��p/�E���'��V=}�w������";�B����K����	t��N�l|p1�a~X��PY.�n맧�������*�r/�sZu�\W�s�]�z�&���2�?&u���7��l~�\�JD��9��S2:�'�n��~ �75uݾ�2�$�d
�����z�������-�4�e$I=I�ٜ@&��pe,���5%�i\����&���F���)!#�4����G�)�Ě�C
�P,�ջ��yv�O@��u<׸tT�xs.�?��%n�D���:�U�3���n�b���$&vJﻱo ��#2u	� f~�T?��{a58u9e{�b͚x��V��j"^ӭ�=c�<n�tiH�M�#��]A�x�}�f��:����W�6b6ǭ�˙s�ӗ�y|5�b�vK�-.�5V���E�v�'9�b;g��R�����Аq&�'����m�?����!�Et4����w��S�ϖ��Cw��Td�xw�;$u�Ob��p��r�ZR��}���Q��+7~�d�mx���k}���������;s�e�2L䍓�ЦĲ�����Y:�(�ݬ�g�;O㦻U�b�dN�h7�����֢�^f� f|K��G�93�����Q�ݮ]r��l�������V#�l�X"Q��B�>����V)���ncU�����T�I�	խf6�Ҫ�2b\3_u��n�9}
�\�on崃�|'|�s���$N~�p��4mH!�V���mꮧ�E^�?���j���A2ڵ�Ԑ��^V�����vFf2�;�
	@<�}���p#�-� ��'����(íj����S�P�ߚ�?�VH�	�?f�a�KM+nu?��/���&\Ah5�vK�N��2��;�Rן����;͑LRU�g��sz��~Y/0kbb���$m�wt9U�����m@L��X�>�� q́ާJ�c���jsI��l,�x[�j$u)Em� b�Q�V�T��2
���׌���"��f�q`t���(qZ�]����Rm��g�E ���3{d��5� �����D7��E��/�A(�����/���8��h���w<j�a�,[�U��{D�&ee�G���!+��2��ʞ������4%��<�^����|ǤyM�����Į�i s�5&�V�r��;^1o��^�K b�a1J�E������\�%\?H���E�b4E��VZu8�Z�@�MsV�}K�����SGJ�z��銒V����~N�1�f�S��] ���}�n�_���4%	ǳ#!o<e���o��ZTs��f��������s�a- o65C���?�"��;��^%�bǅQ�s�0�wƱ_^d�3Y��^^�;k�:�,���К�k����`
� ��&�_�3�3�Z�;��K���o���ڂX׊K#��|�sP��M���q���d����V+�/<���}0Lϰ��G�}��α��ۅI��t��Y^�=����&�g,�H����j����-�@���Je�B�Q���y毻�`kng1S����������J��$1k�4��͠o&F� b��[�0��<+<���z0\D���g-��޵v�rb�g�FGْ�P�Z�����-��A\J���z{�Fm���d�˸�s��հ�{=h�f1����zNAP�/�w�,F,v�_�Bq���0�Q,R��1L�[}f��{�hP�Aϒym����v������#�=	y������P�t�����T~ؕ^���÷#��).+p�$��gL������B��ĳ��y]��Y"8l���d�:�ٗ�H3�.� ���"ҺI32�f������<��2,+�e1e)W�S$1
h遘���,a!���˥��Qط�A̛�x%��q�C\��S(7*U��ߠ�B�5�(�����%M	��B�'�j��C�G�v\=
!�� ׎Vm�FY�bǤN��]�1��$�%�!�{�R)���f\��/K�|�KD�r��F)���D�3���Vϊc�;!��^�:Q�[)@���h�UҐ�t�{�S�p�[?L�?X#3��;�{b��._R�S��&��L�c?"�p�^(>~��e� &1�fX/��MvD�gN��ӻ{���7��tM�O�q!L1���أ� =�%it��$[5n|�A���ڕ�WOrŶ9	^G��lΗ��RD��=�9���γ�^��K�X����s���+xC�&/��	�_���;�3ܨ)q�\qau~�S�l$��U6w���������{s���|��s��.�������v,:kʹ��a�'� ��Ԍgr�	�S %���A|��/s��&s���*�h�LKJd�e�v b:��<�h��5
; �DZ@CÊ�w��g
Oʤ5�O��O��c=�~����*k�Y�����4��ժ3���IeϮ�e6�ʸ4]����՞cߺ��6֊O,�*ˠ�Mci�' �x�#����E|�6��],�-���U\%q�/��Ev�yb,I�Po��+�u\1��M�S�A�u�E��Ao��E�$��%9�L�i�����8i��B�4Ӧn�)������i}�:�����T��}d�AVՅ}Kb�3����+�I�o�`�d�}�6z�U���HNuS��#�YES�ye%N��x�Ӟˮǧ��Қb���lџ6�vx~���7嘛�nSW����w�zӨ8��_&�m�-jV���֖��7;:�����o̞���Pn�?�����M�a%�;��D
x�c�H�(o$7tĿ�9�G7^q��Q����AN�_��s�_����i3g�e|���S���W<`%������cjI~�?���Ю/�mFY*.Ĕ2	�g\��S���r�&��A,��� RRݷcu��]�f��kbh�WjDJm�v#"uV���p���Ϛ�9������F���2S��T'r�
�$R�;�$�B�5��?Y�������ǋ������I+�2<�1L;�(��v-%gu;��K�����_:ot�a"Ku�ώ�j�Pq�Q� v�,��f���ᶃsT��^?Tޯ�������U7Ǿ �}�o� ln��� bpG&������,���9%�� ��� �*�s��M{��j^)bCĺ��p�s~֘\�N����b2Eh�7��F���Gqp.g�퀘�ϖ�xgI��g��c4ꛄp� f3�E<@o�
mS���I�I�b�w���9y�)�6��G����1B��6���B�<��x"��"{���x��Q��rPr��Ie�D�qU�E�Vs�W��yc������1run]�w��]���ɬ�2�A����g�T��(֑雷��=@,#F�{:n�+{Z�H{;������5G8�o��(�*�E]��<1����8U��.�J56����q�YG�D��ßo��M��´$��h�v�d�hYo�DJ�ڝ�
b��I�0Uْ�0����Q?��G��oI���G����*�9�yi�tA�P5��#�F�đ�-�4�Z��.���~w�v���@%�15��ЬSN�t��j�;Rf���W�kK����d9K
)��� �����4��b�H3hN�Zd�1�{]{���B/	rc��ޫjN�n�����7��!�ឯ�ר��A�޽̚A��mjp�;���� cv��[��'�?��z��+�9�^*���<ٻk����rC��֞t��f$
Gg�V^�'@�ާ/)C:1d�3]��L�kI�AL�$Ƨ�{\CJЮ䁈k�<�mA�t�!��BTn%iy_���1���M����ðu�>(��T�XMl:�&.3���p|2�6��M�\��6;qf�Ѱ!Lw��b������ٝ�lB����¶��@�N��!ow0i-�Y�:�-{��_�a��3"݌&��9[L-���CR��C_?ZVe�Pqo����
B�w������U�6�oo��p;ʬ󀹉ps�b�oS�	�*.���0/3F�.�
�p
���#g�b}U�;}�z//�_ڏ�ú�b�V�%!�{����nz^D� �!YZ}\Z�&��7B7@@��N�b���3������B�uX��rW
Ĵ�ף�[�?x��\~���>�Čܞ9Q<}��7��7?��Vb���a#���{.���?�_�b���ג�'xP��}��ǋ@�o�T�9�P��N����X�A�&[�Ggf�s߇����$}  '=�じO�����w�^��=/��S�t*;�c>#l�}�-d5���	�md_g3r��N;2��jƐ��l�1�|����6w�@�"�` ���U��gQ^���!���7
��?|t_^E'kM{t�"�0;�> ��iS��x�@kfb�v�����W�)��ؐ�k[��Y�Z碔U�ܢ�en�H�=!��Qq0�=����}�		7��"e/=ڔ��lBtV�M����^}�11���[-���t,�� ���k��ꙛ�L�3���g�v F���MA�my��D9��"���d��a�VD��P}�iB ����y�:s7՝��S�vK�@lO}*n�+t��2���&+)�Q�ѓߞ���f|;ס69>A�Ğ?�	,|R�:o"������U'�R4��H����"!Rl�c��P1Bm����E'�>m��W$Ϻ|��@l$����Zt	��{f��kub��i=.��[3�(}���
��	V����OkaZTV�E@�7I�b�=V��&{�od
������1���ι�'��o��I�W�A�zE���g 6O�4k���D�/�qa�S	�V>�(}{[I4y��Į<6}X���e��S]�#3�Ҽ!�cp,��/T��?�,	V�;X�1i7���$����Kݧ�3���d���ZS�*���>9�z��~;fKQ�ѥq�e�gR�-�C�KiFSm��<Ba�@}{�֭,�뚤�� v7ׄg�v1�[�y?�:�Ͳ��?*�P`�+>D�Ȓ���I��AY<�Ǆ��a[�D���9��In麹�{O�؏KW���Cs"Ay��J!���� s����V�6:s.�:h!���j�f��D�aW1�ƈB���o�T�8��[ID���(��K8<鰫fq�����}�A��c�+,���ȇ�#F%��{2 F){�z�������QEC�?�����+v��65?�З�ݕًu�Q�۳
-�b�e��G��=)A׍@�s(�ɰ!��@Pa �d�g�$c� |޷I_rG2�p'�]Ă+s�ɥ�/o�\S�蚧1�P'�#��|�j�O�Ğ�,^Z)�C���y�z���{ǫ�Ro2��`Ǡ�?2m�X�҇f�c�Θ�������# �K���4[c?t��yT�l7�N�X�l�ȖQ`��MK�b�٭�@���	]��,:�GfK�I��, ��^��8�X�M�n�L�p���b�tҖ�AҕK�|�[�z.(q~̿Y���Z*�!���U�V�oGP����B���9:���[kץ���������&J����f1퉋���8qt�����[Z�ňJ��R�v�۱���s3D���jAy����H2?Ԧ��p���8�+�|T���>�H`�V�M��T��2��͝2,�������jlU�,Dz^��+��u9�~�W4LSP(88K~tg�je$~�}AaYQ�W�Uyo�!� ��T:e�:ћ��#�����iXƉ��7�J n� �([_�yO�0J��܂r��F�e�s�\��(�r�Z`�(��f��������e����X8�_����Y4��Vh	�g���Tl"��Ufٽ�>1Z�H�����i�:!f�v��:Z���hܚ�-Ӷ�[H>������D�?����<,�3�_�	�7���ѭ���e(H��t�fSX���l���%H?���X⁊��2���E�ݫ�F�X����5�4�Pg�Q�1ͿuJ�jg��{H�-=/��+}:�p/4��^�{��t�p{�'Ϡ��� (èz�a����tOƖrpFΜ��{h��u�}9���E'
�E�3�瘛�G�����Ħ~���V��5f=�)�b������j��:.��ن�6�v,�:u>7�����l���[�k�M�5��\���[�/��O�WP�g�cD��n�6�ݭ�w�&��;$�C˴��#�j��\F����.�-S>�~��_�6ひ-�Z��w���V�Z!��U�iw�3��sB���*���l�nSnt�j��a�=��������o�<��kW=���c�K��Mb�Z[F3�����=c3����[t�Z�`�Pm�h��R���&}���`��K�D��_����f���KGN��1gMm%��UL�!)��Iܸ�k�-�ŰcʨU%�7���-3?l���3��rp��]�\�_�j�^�1��n�+4K�+��M��>揂��]W��y;�b��M�v\�N���p���\�;�7igg���2� qG�<�h���>�j�{�A�M�z�?�p��FM�/�U/{��>ֆv0.Xc�j�����ʻ�����+�XF;0�[;C8�L{��k����O,Q��7�Gp��Gc=�HJV�� O���-\����%�����o�}�G��R�.�4O���v:�y��<�+�B)XI���kA�ã֩u�H�$RG/����c�o�mMc(;<��D�G��p��Oi|��}X-��D��aQREq"����Y ����0"+��R	-���E��e��%�B����.�����)�;o���LP��b)7���!7>�`=(��埶N��e���5?��������np&���SdA6J�xx.�e�h�7�j\̫Y�5���h,�5��q	�;���WrvV�Y����Ɨ��4!8���)�!ܤ�6!�,�l9��6>'��s�Q��iب�Ј#'����:_z��ѰQ��5FN� )�v����v�xV���]t����\�$�l��f����N�k~���}r:��C��T�t��<��9�ŵq�ѱPg�z\:��[��r��vO�Y��aJn(�.��+𖻈}����b�U�"�85E�k ��
f��8�*�D��"��/܅f�ﾼ�İr�����L�%bi�{���7:ǰ���$,z��H��T�����a)�ŭ�9M�y�Ӿu\G%�O���e��GmtF�QW�z�cy��1ɟv��
�S�^l���m3�w����]{��x�v<F�_L]�8!��M� AΕ�p2'��is#.���O�y�|�*dE���&���ށ�����P�n>��h��*���R����>oS�m��j]�'. ���L���>	I]*Ȃ<���|y}!6<$���;3i2�s��7�W_l����f~r2]��2��`~l��,�d0�غOo����w����<�u5Z��bX<e�+��Y���~�J7�?�v�;e�_la��UE����S#Y��z+�0e����\�ykͲ�9ܺ�U$���?��Ų?���5��mC���m��05�x2f�+Z�e՚�r?L�{Uw��^EI[�F��k���_[,��	�/��4����;�ڇ;��X�`�LH~Y���~ӵ\�'�N4��¬��R4�p�����њM�/晢���9Zu�����6b�8�C�e��D���=D����Ӏ��/f̂>�F?����\w3~�q���oI���zN��n[�$N��B�Wc���c�x~+i�aiP@`����^�h>��W�@��yp��=�bA���{�5*|Ʈ&�BGi!�\y7�b�G����;�����,|h/:���`�l�����]"�Kw���Zu"�J�wwҳЯd�^������fT�o��k�0W�3%�ɝ�
�$�*� I��4q�	�=���?�����7[W���G(��Ḅ�ˑ)7������c�+2�� g�Hr�ˮ�hO�҇�%k����L��i�E��|(K�V�Q���X^��-~̳��+�sh���eT�@Q�%$$�CB��E�)�R@�C������N�iI�zzu|�8�|�:�6�~��ڜ���x�HD��Yo2V�~�Wy�9a.Q((f��X�g$��'��g_�l�u�n�<�I���Y�?Y�H�H��5+�
Uѷ���P�����q^��zAD%+�Y�Q�-��;0���
������M�Q�i�Z|GF��H���îs�_��ԍ+�~�|���{E��#�̾�ƕΒ�)D;ē����i��������<A��Sr�{��*hK�_?�G�+��\�w�6�l�!��h��8(	�p[�~�de�s���:���j��nl;3:{�H�Y��x�P�X>pg����;?c�{^����rC�#ZZ-��˔�cG����h��Q�0Ol�l�j�/�Pr��#w7���h|�eW��ڽ����p��d�~��y@�*��n{��b~��U��+��v!��8��w���SQ��Ӕ>�k�Y��C?,y a�'Cgrd��[q���./8C�µJ;��
��LR�BqnH�j��_�w�W�Ł%��y���ض?'��47��Mx��P�o����a$�$���A������}�a��o�p�����q3
�jO�U����E-��דjH�A�n�*��v�.�b4���67��|36���7�~��@_Z������
Xc�J�0� M6w��yȼ _Z�C��#­�8���Q_�D�g�U��ޭ��v�Y�Me�f����J<������/�@'>��~�̨����%S�>Q؆��r�3�F��LS�H�����^ف8�v�*
f�Y6wW_���̜:�;,ϟ��˞�6?i����`j��N���N1�������Ydqv*Ƚ� �Pg媗�߉ul�0�(g>�j�>�0]�q�2ʽ}i�����j�*u��Y����(��^[��j��fY���~q.V>����)ůV�@�2=��YZ��Ff��l=��NJ�d3�S��B���l#ę���vM��"�d&7/u"fmZ�E	/��+��>�������\�n����iyՒ�PM�}���.5�_�*np�<��W8; �p²����1tAUn���H�L��ٵ֟m$х�Rcd���u_���$"�����Volʭ8��n���Sn��b��^��c"�c��of�5b�̱�G[շg�{t�����9��n��I>�����99����~����fg �i�u�04�Ό�6��쪲x�lb�Z�c������C2Z�nm�r��禈"�!5B&�Rtʳ�'"~#E'�E@���}N*S�R.H
b�kMma)�'�Z!I��d,�� va[���#D��$��5�{��4"#�zx��
���=Yp�'Q�dokH���=2��v�T���*t�r �M���>\��e��oݠ�q1�7}[��g{p�)�ʓ�'3 ��#x���eL�G�d^��BĔ茕��b�慨�ad�"D�A����y۶Nz���}����� �̪�y:�}@���Ȏ_��� bu�bo�����-��P��*���Ͳ��z�f���8a��#�=���}:�FAV^$��1s ���;ׄ��j������.��X.�#��]�2��>��� �����ܵ������y
�i$ ��鳭�y2�D>�7�A�Z2rp v�r�Gz��o��Ԥ���ȳ����K͹�νo�*1�q%[Nڣq1E�i<�A��Y�!��q�:F#�r8�����9�'���a�ED�ѱ�C���st�-���v&�:��9�z��X��O�
�v����P��E*f�I����k^#^{��p���E���)���--����
!hH���{I71M�_����9aµ�8���SZɟ��,q�Al�����m��`�-���{!{v$ �i܊ȝ��]vZO�L#�y���Q2��U	vtY��)���L�&AL�/]D���3c�c��� �}����Q��Lt�cR�qH�))1�ZG��۾,Iy�iS�kp�^�Y��Bo!��>t�)E{w!�]���J| 6�귡j�%e 
b��l��+�ʱn�ҤB	��B��Wސ� �ϛhM�g�rX�S��A�8�	Bm��8���N�2�E�szĠa2q�q�o
}�!
f$C}���Lz�1�Kt|Y���/�|�F�bAi����&<y��=�G�p[ln�8(���G����B�1�����c��`�lz�ٷ�}�$�xE+ ���6!����v�� �fwo&�UN�x�%�M��	�J�w���������9�`ݰ�0��Tz�bAf}�L@�
�J��2هp�d2{�Os;t��X���-f���A�.�CJ�~���1<������Ě� v!����M_'��_��81�� A�(ڬ�3/[E��E�A,�j�靎�qF�G++<X���@,�\v[���UJs������j���8�;3�֝+{L���I���#�9D�CA�*>%,կ�1Zb�jv+����a��VX���O@�ܕ�C��%	s�D��0�E{��)5&�^8������N�dA>���af(0�����I����Q�Z��Ӿ������e�e� �=\R7�^jd��}
):����Fb=��MZ�b�5L؆���-����F���Tրbn��;�<�	�������q�����L#�����¤׸=J��.��|����!��ae/t9���sE`���}�ƦBĨ]K���N�;xƠxp�$6��@L�X\�y܅��i2��Xݒ�
��%�-���b�̥/C�*�)�1�BG
	�d	,��|������@��;�l٤z��K���i>5�R(t^��V?�'Z����t_�1��W��Q]��Uq�nC]z.2 �߉�+���(`d��S���b+<������P�����u�(�� ����ig����=i/b+A�1�7qSMK7���A��DE?�ө+'7v�c(�T(�)���1�We�����C1�6A��Cヘ�Ķ�a~���+C�h+�K��3c�W���t���}�:ӽ{4Ă b��0"��E��8&�$��߁؎�(Kw�9䙃k�-�������j/=�_Sg�m�����׹bwN�=l����7�l���7�`1��4��3Ҩ�Z���σ(A�@0J�Γi��฼;���8�
8���?Z�������
b���������͆r}�~Қ f��
�coS�ɲ#Y#�hAKb(�z��˛�CqB���>͞z v��:G�/硽9�-ՃR��b9k����eP�כ�z#��3A��bJ��s�؜2�w���&^ ּ���L@jj���ԏ�qQ��	Ī�]t(�(+��`,���jѩ���$;��a]��܍��jd�2�Q#}��_L4�Q���el9��D�=׾<>�zNUL���@�0C�oǚ�4~��9׼%y��=�'�[gm�]��yO�m:+A�ݮ�?����t*�O&��!�ޒV5��YA��8�j$#��&��-�j�������[^W��QԤ0��:y!��t$���=�Þ��c���S�d�:�pR�1�h�T��@�d<���e�5�����[��*	�LK���R��J���ڡ������F��3��y�1�����Wi���(��,\a����}U�_^�5��ˑ�Q�~�i�;��a�Ր�6�$.�$��ܫ=�#�����n�Zť,[u�D��W�7��Z��|���h���A��_���;�8sDh���?�
ʦ��ńc���Y����ЖnUoO�&`<�Էߊ#�3Ֆ�V�N��@��%6��Y�K]���^9�B���~B5z�ʚ>�Lam�]����~@�׎���Y1.֭%5^BW�֜��D���0�$���9#m
cT�f�D�1\��sn��t��X�L���FIQ�'j�-"�&M�<���A���F�,������j!�[_^����N�u3�x�@��7;�rr���de�Q�2c�V���|ze���n���='�Im;�y��J�c���
<��'3�Em3���(�My9dt��KH�Ŏ��� �C�]��i���%�wKk�+����9ᓯ�N9���̂Z�s%����	�j�T���A���N9ܗn���5����T1�:}(#ӣ9?6�`z�ոw��Du����g��
��Vr�_��e��ZK-�o�����;�$���U�ػb_-���Ba����3��Gׇ5�/�FTb9͊�5���̗=�?�BF�S���nH#��A?}_�$�0)��<s�ȯ����\V�;>)G����bk�g�'Y$�8'�M	<�I_��5���Av����n����>�� �������s�:�*��r8A�{a&k�;뎪Ȱ��+��ݤ���JV�ʒEg�y�����(�3��+���,��c���H�Q2j���j-X$$� B㵾�y�G~d9II䠟:���r����Jt�Wid�6���%�^�W��,^&7^�����!��H����5�iu�T8�7�?����wUr[��`ޥ��B�/���D�?٩҄���߈��B�&�Gq�q���Y��y�[�_����0�G������D����>��7�s�Aq��e�{���	)�*�S_:/v�d���u�χB�?�I"Z�'�/e�iJ��zQ�?j�+�34���
5}t'���P�B�4)�Y֌�_�($Q�"@�}x�����Q��C����Ův��I���
�������'�˼LAL��6�W��0��2�rO�\}K�\E���2���T��z^1!���S�d�N���~dx,�W�ҙ@�����F����&QG���e���-bvp��lf3�o݇�����x]�)�s���n��_��|�����հG�~7|(V�\I�=�F��a��XD���̎m�!�i�F+Dx�n������"ϛ��1�&��j�����Ҥ�oO���`K�a��i��Y��_���%ן����Ȥ���:Xul�"�<\�bᐭ]���'�KYY�`���;t�I]��x���-��5R�W��^�5·�;���JW�s�t7�f�U� b<=�T�� ����s'%C����-y�M%ﯲ�����x=Ѯ�^�n��ڒ'�X)������:�W��+�A���3ߨ�'���T�@�.��W�.�/�H�k�W,�]��	���g��c��8��@O�$C�o��"�3F��-na�.1q�ցj�ڙ���j߾�:	��Ֆ�O>��ƴ�b,J\<�"W�j���J�&�}���-�t�4�p��FJ�.�<�O_��Ǘ�"&.���)�\d��3�ͱ�E�<:�~��<�?���l��5���421�����ҽ��SD3*#n~f.�fD�0�U�1^)9+����/M�䥍�T<��$o�}����{y��
���.b�*	TH�@�{ИW4`v���ܲ ,��[�G0x���f�u�'~}Ǥd�/��l�ðu�A��H�<��:
��c�#\�".�7#�3��r�0�vB�b�ȤU������nil]Hl�.�3�l�^$�.O�/&Y�#z����k҃�+r;ct�(�1��HԜ���+���#��jeZƩ��i�ob��c��h�=e�1/d1#��P�zb��g�F�7G_�G{@>���li�V����a�ﾙ��R�ta�V@ZP<���(�[Ȱ Vf:F4��*i�|��MO_f�|g��w�M������!"˳1uB�S���W2j�lD.0A��R�ڢ_l{��n��A�Cѫp���RT����O,���t� ���7�0^1{�:q��@��u��.��\�\����䵙��A�7�eХ��k�<���Yk��[ٷ^\�b�뾚հ�U����B���,����x�n||���?���N��rK<M��6%����$.�����NO��sU��﷽G@r��{�_"'KB�S����br�tA��$�"h�33���G fuxI�.5��&#���&��WːxI0���h�a���q�#�NC�i�A���=���j��+w	�v��_�~�5�TP������h>BV����j K�*Ţ���e �i�U�tV-�ͫceD��R�ѡ_�L*���VH�U��%���i�}��6sk�h�M�Á[&p�gu*���]-���u_M��3�!	=Ř�C��0H?Ek�����Ȱ�d�f/�bo~��^�א��zl)����f�����y�R�a��k?7���n�&�2=!���1���wuTS ��l1V}�^�!�e�ms�Y�.�E�O5�G;�,��j���)Ň�ɦ��yW:q�ȸ�����h���aE 6	�'b1,��)b�%��:q(2�G�tL�����b~C�p]�[f��)1+���@,p!��f;,��d���]����oCp��T���G۝=���v�~���A.�E�;c�[�6��{&�!���$�g�ћ��Ъ	����,�D����XԨ;$��k-�jm,¦6���L��#�E�e�&AA��E�ܟb�S��(��/.�-@�o�����#����*�K��;e� �����.�v�f�G�B|f[ F���eo��T����̾?o?���k�v����@n`�5�Ʀ�A��ȱ����Z�-�O\�s8�1���?��s�����$�X��ɧ1�EH�,��O���p�9���H'��><)!�țO[	X�� &U2*Q�q���Zw�Yu�	�M��֔�������?D�V1� ��''��Ɉ���jJ��G 6����'ks���+�3��b�Pt����l�-�l�3/A�ч᮹�u�J>~K!hU�*���{��k[l��V�Y�|7=�¸�O^�#&���__��I�����)�:?{���^�1��X���`�K����<�.�$1Fu��:��ڡ��`�.ce�^�i{�m�H��ۀ��<�t.��q��> �c�i���K�l��(z{�IC+�eB`���Ŧ0zvⶸ���1�a�0W�\?��;��j{ʏA�� )ȳh���w<����	�����8������{$#;�{KF6�{��^��eS�C�~����[w������+V/H�Ȕ�Ë�|�OoC�ݧ���fv�k)�u)��Bg}�o���s~yM����)�!��\s�@�J�����u�+���;��i�h��`��A�^�Қ��܇w1?�gSp�����"�{C�F9���I�*@�\ݜ�kU�js)]�{��Fra@��I�l�$�k�7��q���Q�A�═
��媟�[���qu1=�����*�s=�T���J����5$��~t�_�'� ������#�焕�+	#M\'��p*��n�_��_����cG�*c�� �E{S�/�j� [���m�٬�%�$����{����?|�����x�7x��
6=b��-4Y `;�O١S�G�׎��K�`g5�#_�02�"W��7Õ<�z����3�a�ԕP�M��e��$�<�5�7�%�����h �3s���[wﵞ��a��]���S���2L8Z�F�tc��~�I6�_:�?�D�MB�	�˻�#֨
����/$2H3�KV��P^>Q:��Θ�B�A��F��}�]9"�-3�
A���Rcs��wE��o���c��u��Ł�=�����I�g���eG
��`��x���[���(�J�=����W˛v����r�a��?���A�N�x�K��~��wCi�5j�b97EP���,h�~��T���ƪ�f��cqeL�_�Ň���ƽ�\�)8w�g�[ISj(����w+#x�8�('[�6GHf���8����I��/�׮����TP\Ǵƍ4b7���א�MT���o&��W+�{��d��v�W� �l�b��U��_!����φ-% f ��}FKz�D�o}�ᠭ���� &��U%�b��[?�_>S���x���?5��&|d�~�ʇ��.�g����������[��J�"iA��(eg`)�����oM)�WJ@,�v���ތ܊�ڛpU5�����X1d� _��k,���-��+5��=�E��Zha���Ս�Cm���1,�C���k<��fv��EUoU@����1���5C��!�iQ� ���? p��^�:�}�;�7��X�x�"��&'2q�V_�ָ�Q����=eRʅH��xn�K��.E� �P���:�O&�)�:�q�=>��.1S�j"(�<�s�d�<� 1��1��f��~��9����A̰�f�=���PE ��w?�;�=�HO��Z�J���_Cҡ��!�u_�vM|L��e�t֢�y��.�N�/����v�~�x^�q��b�r�#��ɐd+B�5PY��&��Alt#��]�FdX��뒉�o�b	/"u�82���������1M���ը%l:�\9�=f�נ�.�ƅ9MGYvo��hJ�
�zЃ�*��Rw�Ux ��%-��[~ 6S$I��t~�,`���/Vق�1���֯���1�w��A̦p-Q�h��Ѿ�L���Ky"�=�bvz���_�S�Ƞss�*nĆ.����r�>ʖR�?��rt�	��${�?7'#Jkٳ�HE/1���2�̔29��#����B�J�UkQ����Y`7~����,_|
b(\_�]y���a��A��s/�Zl_�{)EsZ�Vٞ屯�ŀXq77��z�i�hc���?����ٖz"M{׈������r�AL ����Gt�a.T�	W�{b������%�KQڇ�|Dw�@��	��SI�Wʆr��vX��Dc���g�5�3�-*��2h� �b�/q&��;PQ�h��#6%��� �l<<��tY9DF��2�E�y�,���y�טn��^>b���������\"SYlT&�'���h��o 6���y�K�e�ڀ ��YE��/ F�=N����+�'�P$�)
b�	~捄������+rE���AL��dĕ�����&zE>�G4����E�(���.6���Xr��p?,<���׉D�P ���=c�콦��Lnl����c�N�-{d�ȈE��4�	]��[jhb]����0�SU99t��p�������u��#W,Of���%;�;3�) �,ǻo��z���"���_��'�sPT�3mbɳ�f�7�z*�X���̺���*9C;���QEA,�k8U����b�BV1~U���_��E�-�
F�A���3�
_}��wx��4������9����=���4�Q��m����
�R �'<s��Y�����OgY����j͛=���0�hh"�EJ �c�dw�΂�c'}� K��]YĂ�յ(qS�!k�w$�&�@�-�l���cSJָz����	+��b���bj�?��0��gOwO�1/��w0��*��2]'f��'1J�N�qz��F�������1�g vBry�	���9�Y�K9U��a; v�:�ŋs}���z!��N�����W�i��/�$�|�9�ȳ;ӷb+2�ۄ�]�(������K?{��N#e���$���Y=c~H/�5�I�{��N��S�+��O�&b���ۑ����Q���xka�-���M�F� �1Y���Y�uĬ���P�5�{߶�Y�47����N��y�T~crM�������^ ���m�$$�ɐl�W.)�S f��9(�"����o��%�^��bλnO'��qEfѝQ�6�&$����!�W�����<K�pAL��k�����A�elրyh�İ��S�T_�mb��ojT�<�����<���<�	���}�b"��5��~���%����Pbn���2�b��7��1�3�\�" �����Zz��']\T6�����.�pQ���Xq�t�s�q�L_�ɂ'���B1oN���+x�)mq[��� �A�$��Gr�nB�]�)��4�S[��$�Ə�	�����;Đ1�yWR�hA��m��`Ȃ�3#;����-�,������<��2�� LX�yS��\��I̞� �8د���M�+�|Q@�8��bKe�[�ro�I/5�Ӯ�G�X�#�c�+2Us������� 6�v���Z��R�9�T��zC��s��!�L��R�L���f@��h�1G�V_�9\�D��C��ڶ)}�jWd��5U�P�p���A�J{���G^�7��:�ذƀ
1�ɣ���`vB���@L�Ζ���u���w��g�T�J������h��Zt+e���9?����3h@�j}�ʮ�iI��Y��'��wP	at4��gG~� V1E׃�+���'/����E���!�=��p��s�;R;�Ӎ����w� V�S� Z�2ydТ��|�h>�!
b��*d؆�z֚E7�ϡ�Fj/A,��
���	L�H���S�Ѽ�P-o��C���￀V����\���IC�k��KbB�(�tj�\,o�l�:6Q7�͜��䜚9�]1�,��.)A�݋�����N@�y���;}�hB0�*a����ݞ���U)����8]e���6�:=���&����ɘ�vO�@̎-) 'kÿ&�z���1}R���&G�qI#+�r,�|$���AL�7�2�?�A��Ĭ��4����_L~�0�8R'M�C�~��b�ݞM9�C����\�,;�g f�Ɂ�ם�,�(Sv�r႘�HV�9b�{���6�.�U���p�zr�9���ǳ(���[V,��$|/,6i$�](�o�n��=�g�!�A����q�jH ������+ީo����й	��X�Q����̴�d��]KA��x�w#����.;Ly���̜�΃�j����������|;��'�@���f���\���M�[n��� Va������x��;�d���R�Y �f�w����R�|�ާǺ��l��@��B��| M�qV�Åjs�h�P[����[�2�BB����� �J��m�>1O������C�;q��)7�"��O��`�������g�k�	�aRǩ�!��:#���$n�)���c��_���Q}������:�8���NB`iq|͙�Q
�M)���=O�,�Μ���LX&�(�TF�n����/�v�XG4�	�캡���9��(�x���bsG6n�r���nSo�8�|F�@��(��Ҝ�fV�Ȕ�3%�l��+�9N�f�����8mF�Odz �'b9�dV���m1P����З� �{-� ���Sw9��Klu�2��U\�q��O�]�|5���)������$���y�3��b��ƀE<i���(3�g����B���*f]������*�1w���4ǄvNN�1�Owm��ے�c�X�䧷٬�yY��0oN!�A촨Of�ugI���E-�J�d˸S撴'P寸�J��iK ���s�����5�r��E[��5�(Ҋ��I���$��f�ui�X��e��h��UF�\�u�kkb &40ׁsx���^�A�]|~!b��o���8Q�.�9��$�:0Q��x`�R=E�⼅��8���d�jCu��ju[�A�㖅mGl5��ĥ��Y����@�X���ӊTs�n=���m+�bX�} bT�V�v���Mܖ����*�A�$[���Q�?J�.؜3���Ăk��.�y��m��5��Z���zyu����q}��̣i��X� gA�w%�Ė\�:E��G�R�����ͯ�U�	����U�jp�� vV�ت��|R��u����1�mxt��Z�BK^q�d*x�����V�w5��m�0^Ue����c;�A,�`�?XŝYC�K�B�LkF�>�);Z��u�oN����t�d8o��)Ǻ��۰����^:ܠa>�nS^/�ͶJ�����J�<�2+Hb5���:�/��ה��d�>�|z	ĮGu~T�+u���~!��۷{
b7��l�V������4n������Fh7���^g�����oQ� ��|�ߎ�3���;қ�[g�z8?̦kP�֐��'t����Oܾ����!�FBB�NL��w%��3���LAtt~��i?�I(k�)uEMW9��Kw�}�1X(g̾�[�Y|H��~���A��LR1���2g��5%���>H1�d��QG��f9z�=��9Aʤ�2��3��y���S(6=x�rE!��Xnf̜;/�7V�M=��f�4���i����g�b%�YU�SL�B�N�N[��m��������K�3�b&�~��x��[��<Z��
�Ā��=S�0Qj�*����È�O���<�@^���y�v�I?҂���ؓ�w��w�5��È��U�MɷE��f�(i9'k���n�J�,̯񏴭��M��p	F��F� �o�M�l&�VX��n+6��A3��TF��u�ܐ�C��礪4z�e<-�b�dtHK����9����2U\z��w�%�H�W�|��G"y��]Њp�F?���$��Z	�q��_����Ҷ���S'��WA�"��^lT��q	�����u �i�~�PRg�H�֥��O��C~�
�O���[c$e�.�Y�Ch~/*yux&�{~�Z'a$��wc�a��Ɗ��HK���cg����gM�~����4SLj�I�0�u7���d�uǭi*�|�gB�)�[�#�8���pŷ`*����f����J���=�fX
��{+%����-_(iH�3���4K���w߭K�3���N<�+��ܷ
"�{H��a3�m������[�/I3E�]��n�fT��iH+E�L��6ُNi�Z����#X���-�=_/��T�z�$£ݍ�v�4�I�d�u�
�A�r~���*�1��|Zp�8h�F���Ͱ!��W���/�vH77��bC�[�]4k[/��7����)�G�HU�p�r����L���rRʏ���GZҸ~2�U#M�O��6�>c�7��'��w�~0c�����~�m�$$���o�~;'�a.�����,�
'AZ��D#�k�¯�m���s�|� ��n��c�	���EEZ2��~�ߺ#���e�$�i�o^�н�S7!�`�\��+p�o�r��_	�Q���,���{}�~D\E��γ�n6�\��9.z.Ҋ�ƅ��8�#S��&�[H��%�"�?�i���/��Ū���+2b]r�k�����RGKXb���Ѯ7g�z�5�k�=E�k�e���vݶ��s�����]�C��]��1�Ȅ%�/�YU�G}M�[�R��u�c'�'KFZ���h7o�r��Cmv��CG%y+nd��v�5d[گ���������Z�ד��I�{�ے����_�"�i�H����}�y��PE-f�%�/���d�;
��8����|5Q�Y�^����Rh7I��Q�����
�5I�}��W�����ި���J�#��z��7�Zun��E����21��u�0H10  ɋ JJ�P^
>��g �Gdk'd�9�(tm��)��Ma��Ma�L8�kawh�d7M�8���)�܃��KB�_Fʜ=9V�w'�_����{|)���}���م{�_(7e   �  8�{���Xq#{�T{�l��=��ݔ���b?<�[+�*pl~*��=Tݏ��y���>�=�*�۫7�aʥ�
b�?�z�i-	���p��g����jҦ�˲֝�f��ط���S�jfN��.�<3]�msZ֌�_�9�t�\�1E��y�I�A����O��{=���,0���3���~0�:�����"��k�!���,���>ݦ*{m~qT,,V�ٷw.\B���-a�<��X*��P�,y����gJ,JP�S=�����fR�\���TsG�����t#_Ͽ3��lŮ���=}��k��G/���"E���7�Wb�iUk��-��:ݗ����M-���̗}��e����\v75R��Ny��Ѧ
�+�W$��?���-����L�[]�3������ƴ�U����2s����G�>>Y{�Sq)b6�b�~^Ş�e�E��S���"Vc 4�^iWbҾ��ign��7�7)b�4�,��i>����}��i-�[���P��j�+du�"�d�\u �}u0���몇{?(�U���S�r�b�؄!��1�n&�������y~Lʓ2��y�\?F��Z���]l�lit�Y�+���[�Y͵���R�y�򭤈����`��  ;��%�����z/ظ����   �  "%  h���eS��a$�E�n�V��$���A�[��ii	�nA@��A�,3�ewv�������G
�Z�d5W�*�3�(�����b��_~��N���"��Cl;x����d풯t�L�3���孯�n�F���- ư����O��BIO�e^f&�tH+y*t^@uY�"�.,c�b��i�{0��k<!uQKJ���hbu��6�l�'#A���e6����3�3֮�n\���I��'Ą�û���h�ad�m�nS������^���y�]L7\����L�G�k��Pj�K�[��7tdϡG�R�J�q�[��O����q�Z��pL1d���E]&њC~�7���`�qG��J�?x]�V�F����{-� {��I"J*�c��՗4�����<���'�#(�����+�2+� &O�Tj5�t�B��W}�b?J>gS�a{�B0z��] ��N���%����Я��ʄ4��l�igkN��.�׎eO6��᪔���'�R��q
�~�Z3���Bܹ?�9�4�Jr����8�I�9h ���zl��}�5lK�HA+�M:u���KM� N�7}� f�p�-~�Ĵ�!:J��Z���ĸ���zS�_����B�.��k�14mXq��Ʌ�X{o�k����!�쓘QV��D1os��R-�1Q����O��AN��Cm�*e� �=?�4-�22Hs��$�
oG�i�Җm����E��p���ļ�H���?�eܢW\Ah��A��{7̓���|Qi��Tct�b�~��s�Gx��IgO��a�E���� �ޑ���<�>��2��E�$�MLn-%,�/&i�����؆W����MHc��OG�eB��3�AlֱP�Ķ���*ڂ���4�r���A�yc��_�-0j@l)V�����#K9zU佡�n����P���-��R���(=1-V%ʕ�nc�F���C�v�p ��;�b���KGw��L��-���/��%�!�EKM ��$����J��6�����W�u��O��!χ��Vj�Sd،�ۤ-G�/l_��0�CYɤv���ٖ�
b��G��=�X���j�)��Q�9
�E1�%T�V�`Ϸ���?:���<m5���6�ex4qXO�z����WR��g�׽�� �q�c��+y,�<�[����[���#3YL�MH�ir\�^��h�s���9$�E�F���m^���I2��6�յ�PwtOo�MR�l�%�C3G-ԣm2�N��]���
��I
@{�8���s���"� ����䔁�C��1/�+Zv�"b9"�á�ހ��A��h��b;ҵ�2BU5I�Ws�mg�0*�4��	�[�b2x���.zo�Rn���}���mQ�oC�h�p�a���Km�M(�!����a@̷Ĵg�<¾ɸf��D����kb��8�{7Y�*�I+�M�h�z.��!c|=9���ܛ&�R���?ńV���$���t�~-�n6d��A�6<��L�D}�iџ]���_�O|�1ߣ����}e������0]
_��tk�F��&�
�9)���t`g��.yü�����L3�	�Ք�?�㿐�'�<%��s���p��+t�DK!��"��U���������zʆ=��)�*�}����m�BVǇT��fJ%V��J��������������T����G�{�:�_���1����}�r�V~�� �QY�4ĈH�c�'�H��>�4e\�=�y��٠'zN�
�vO,���bm�S'�7��K,��ե���_��C��uw�늯�|F�v)k$OЂ�6���y�gg����|#
9���<�Ŀ�{�!�Ī�u �f[� n����?���k2��\tƯ�Ewg>j?�X�І�&���mR��O�Qc,O�!ec�S,��]��)S��3��VЊ����,�@�������~�j��h�ʌ�u%_yHa�3�ď�1Uc��ؒӥc�!+}��Z��pNȧɭ��l;�m3r��0{����24�/*�/�0Ҙ���kHb�2�E �?��
�ϛ~��Pj!t�3�)�2�H�J3(EO���麧t�λ�j���a�(�T�p��s�΅o�`��s�_��
�~-ox�⒚�h�[���4�3d�qx�#.�6T� �23x���T:��{*�m~��A���PRx�H�?�*%��{>1��������K.��� ���6zՃ�T�S��s�"������Z��f������M�en��Rm���bu�|������~:�7X�������x�yv�m��q$ǍA�k{�}+�*'@��,�R�f�6&�z�������n��dS�S1��أ5r�"���@�y�0�)�۝e�U)�hJO���&��-�D�\�^����9S1X��x?��Z�S�$Vi%W�6�����Է��X���΁�(Qң���W�O&��Χ���7�G<�T+���[��ۂY�����kÕ./cO�[�2<'�%\1��U̪�}b�h�B�w�a.��1��xCn�
 �ը�w�d�bEdJcV��m^����5�X�Ub�)h�yt�u��د���
[<��
��k�dt� �~3��@c�`�)�4j`��E�
b>R�*�J�d�XH>-�V��1����1�A�4TD� 7��! ����ýB���l� �lVbDs����w�k�체�y4�A��+��xm�d^G�&��*��:�Qj}��nK��7b�~|gb�)�v�|�/O\�<kNKd:�Al��H���°,��hR�C
b��U�L��4B)��r��A�!��}5���*���F��L����aC2�$�9$d��h�,A,
�w��-<�e��o]x�YQk������G��\u��c��a �XKu]��U�?�ޢ���������`�0N�q�XɌ�o�9� K�J��ԾX�f�,|g��Q8	b�N\S���,G�&S	w�K��@��&�}��R	~��T�Բֆ9�����2E)R0�8�����耘tNe��&ұ��wM�ω@l9�`��ʵg9޷#�v9‐e��3��\^4�f��H��n�D�1��w	��_U֘���+�m��XL,�׎�\=�K�(<�["SL��q�+5���yx�b�%��oWwc,hloH��z�6axI�[�Q���2�e�$,�%����rKf�x�"�76�vCK�	ľ���,[m��)P/��_ă�{b��{w7H����bhf5�x�� v���?*,�jh]!������� ��7�deHq���F�9��CC31��$�g��ab�ġ��HEK�	��&oj�ָ�}u�;�YdX��*w~��r��cB�\3�'��>�:r�ߝ��Џ9Nk��D��>n��������~�P�Ğ��R���G���:�����Pf�����l[M����9�����H�K�|}!I�j�Z~;#F &1|/��k��{Wm�,r^O	b�����OƦ�x�'�O�@���b�E�i$�~,g:Nrb��,ŷE<{$ƻԶ�y(;� F(ZZ��չ�;1[�"��}� ��)���	���P�r4MB����j�*���Z���M�Hk��PF�5l��Z?��`��}ϵ�b<o��3U�3�����+8��@�ی͕�x��F*z�1���,��2�z)�o�7�.x�L�$">q}����Z!uI#�tg��	��G] V�_*������7�Nx`��3�!RÍ �=�zS�dm"�dӃ��n'u�����,�|����z�_8��c:.6�w3k�*u�1⅟k�)ϴpr��e�����y[�No8Z�cwjLYFv�uz1����X��/=;�������8ĺ��X}6EJ�6�5��������(*�٘q�PR6.iRkXv�"�	e�<Q~7d���Ҹn���%39�qȜ�����:O�O��+|#�0��qx�@+�rڗ��(6�I�5@LC!���/Zene���m��� �밠g���+��۴F.����4<k��e�-\>�	<|�?��	'�t�?�b䰓�N%�
��%Z�Ŀ�㥤r�b�]i�a�.�u%k�����@�@?�=
M�ԛv��73<-l-��B]���t���{
�8�Ӷv��A���$%)�@<�9P[�ӯ���ĸ ���{���0�]R���OA,{Q}�1-J'[�aq�0i�E�v���R�R-�e;%}r�
-��@�����e��kz~�+�N9�i�0���xń�th��*A�HC�&v�^Ԏ�2�'~��� 1��}�%�r,[r\T�)��J�_x)|h}���Y�)�S�xJds�`1�i2
�q�6x�i�<���jN�H��<䟊]r.��leZ��] ��X]��p.s�uLF�Il�7�p�vG�Mbz��`_br1+������V�� �q�u/��@b�]��7ݶ���m�k)\��k�C��`�����m:�WƖ�<�����W�Dl��{_}�;�A����I��Q��.�����A���&�U|Hb�x�a�Q�����y���D�����>~9��`�l����EIv��	(�8���5S���C`�#�f��|�f�q���f����'S]���%ќ�`,y���t�;e���kVNL0<����1�Xr"�<�$��� ������۝J���u13Y�o�L��8@lh8uT;�ޠ��v�X\�9��b�!�vǯ�	)e�M����I���C��t]ւ��Ȓ �\�������V�R[��Ӌ�� ���kL�q?��,�N��O��bG_�=�CWH�.S��{��S;@k�͗I��7������������bb� �aι��Д�m�XU���6e {��m+y�H^[y��o*���BP�r?R0Fq`~��&��󞠹�9�4�l���u� f<�u�$\���������P	�VܙB�1��81C�d��:,@��ӽK�/�i��v��� �Co+�¦LS�$�F���W�b܅)���8�j����E/�E@�Wm�O�w{��b;~���d�P�:Tx��N/��k�����`����]�iC�(k�߆�nU!b'�a������_-������?�����F&9����{i�鎻ch�7
O\�Z�Ē��?�8_�}o��|k<��b�~y_z*�X��Ό'���o?1j{��o��_�OVR�j&A,�kqh��AE�;������p	�h�u]��0��o�D����ALHb�����[�����rkL����Ҵ�ryS$�z�23�,�-�Xc�<���%E�����}�I�� �@�����fHk^��1�&�FĠ��/���������l$|��J���i��-��儕l�`�"v��k;�����nT��`�dC,!l��Ĥ��9R�8��7�,�mkAf�mḕo��n}}xZ�[:���]+�H-mZ��^��Eقb�R8�z�1>�7[����i�NFD�V��>�аӥAMcb�ϯ*~�Ֆ4I:�F\ǡ��q˂X���k��Ye	)Vy*��� f��V�M�:�a�^�&~��Ns^[,�)M'-�cN�Y���BD 1>�=���R'��P����/{E�@�Qy��A>|IE}e6�,]� FV�Gg�b��x�&�kb_gbj����'������{��v��� $m`hh�)O���$���X1#?�@�d�\̄��������N��脎�ڳ�a�Y�+J{��o1�,r%")���i9��7�c� ����w@_w�m��#�7�,Ĉŋ#3����9��]�w#@��p/�v�!�&R�M�1�G-.��$Q"���e��'�}b9����� v���z�+���vj�;,�����dQ�}�P_sۼ���e� bk�pU��*m�aP�.��;Yk vd�����_^�rFg��ݾ��(�7̽�>*b�c�7{Fk�ԁ�%�`b=����׋h�4��Z�E��_�Z�&�@���j�M1X���!��e�$�SO�Tn:㧂��-��d(��-��A
b��8SN��e۞p{i{�5$�z &K�n��ԫ�n9@��:`���jc<�G� ��F���ȩ' 1X=�]�IJa'��c��P^�GH &�M��j�RC0��#�,i*O~bo��I�/Tqn�}�~�m--����@�sQ��KY�ooNl\V]�@,Ϣ>A؁�Xi{��p��~#6�q*��&?��k"-�'�g#�����T�-	r��穉P�9
o�@�S���;��XWc��o�V��D�t �����
�4
�9�>�f���z���h����# `+ٜ-#{$�JVo��Ȋ���u���rdfd+��蔽
9�8{���2���{>>�yEd}h
ߥ��lǆ�Ԉ�����b6�D=�1:��L�PЂ������J�OR�n�U��gU�u�q��ykœz�M��~������p�4W62/&R9��s�c�bd:���N#�Pj�̥���i�f˕9��;�%�6Z�??�ϭ���V�[ōދ�fa��͟�JF�t*�!׎�j��l.��wsE=����0�a3uė�p���M*.��Y��w�d���f���G�T%���a،N`K�0��2���5:rU�_݈�2�n�u�ܻl�Fȕ�6U����u4��6+�L��9�`2/?K�w8��👱/� ��T�8���R���[�T�x��9���g����M�ޫ�G.�R9�[��>��%���T[��rg&����M�tz�=Y.��vU1�Og���r�ȟ�_���aR��ȣ� GԞ�O���XO��#d�Y�jB�/'@�u�t��܇{�����&ȅ]|���(,�8�G�fO'��+ ��4[���EL�������vVT:����<;gC�r#�|�=\���\�!$�(g��Ul$CZtr��b�e���t���b��Z_�C�y�q�}=�j�қ�2�f{ѻm�C
=���fF�۹�h�.o�f�!���N��#�B�#�N��}�]7���g!�=7�����v�O�y(�'�sn�uy���6>�hb�0��B/�'�O��r�\�b��I~&�"����^a�\�`��#Q��sѴjK��9��d���if,�*anǵ�S"�0�-bQ���-Z-��jK>�����ͫ�%�aCV��j��F�����4�J���j3ߺ��qe�7�?5��k'�.B�����>�w��;����2S}, ]?M�2"~b����Nf����r�"6��G���)*K�c��lW6!���GE!KT�Ӵ���V�B�8��*`�bR�s�h����~1�m���DP�Pχ���Z�c�\ C�PK��d����9�q��r�©xo߀U��}��~�2�e�� ���8��(�������^>���NB�3�Q҆QL/�:��J��_Z�[Z?�֓sx(��%����1���.���Ag��9���2�aMݛw#l�
�hH��_��X3�0
�i��x���9�[a-�����o��)��iC΃o��X)�x���ڣ�u%ܣ��>��s�5��!�˙��w�6A��-_j.]��Ѻ���kZ��J!w��a�����άRփ��u��ȡT��ZQ��A;�����"� '$<��i�^�˗ٿ��DQP9�xD���)-��fk�Z
)�bH�M��|y��:���E?��E/��%�96�L&�G(�����#���d��t�51%:�q	Y�(��9� �I	��k�A�����{s)MbӐC����t�n2Z2{s�q=�)���<P��>�h!��[5��v�E;�!�����|�2r�s_�3�`K�ES�R�֢ђv���e��軏�� �g7��7'T��2��զ�Z��]�ܤu��ZKO�G0��{����ѨCN|�կ��i�s�)]Q<}Q3䊔�WY�>��M
�٥e�{�I$sT��
�����Ё͹��r�lm�2	�v�ӌV��y��M!����K�nqS����i�����7�g8�V:��;�xn�o�Bnĵ �l5eȶ�$�>��ziߩ9/��gJm����W�LE{9��
��tڦ�+�����7�~������9ٚ��K�j��F�ޤ1K?�8!n~�acO�A{;�>�?�	��:�^�B�fG���~����(�-�!lߑ៺�#+�0Z��>��\G���eѡ̃�;y�R)�4�BO �^��S���1�[O�q��k-�%�vŜ��ڇޑ��s�R3��!w���`O���ӯ"�>�w7�rX���t"驦M	Ꜵu�*�rO�&'�YurZl�-m5�r��~�1E�l���繘n#���J�9l�i;G�J�A�;�d�5' r-�ϼ���ڐ�-�'f)(
�!�+e~o�yܩ8�rS��b���p��m��]Y;���o?����r���̓�a<�򃔶�ǘ��I{p�4b�,M��Y.s�!.��JB�g{M�+�S�۔�-�_�ŭc�W ���c]+�[��6�Fa��Q� �E8
�3��
������^<����a�8Gq��0�A,�0��C�i,ɪ��j2���(����d9������C��\��S�5��ʻ�ǌ�ά��	n�-�\�=N[µ�X[T��a��_<�t^ab��f�x;ޚ��1�n�[h��jk��Z�w6Y+|�O���>��>�ыy�Tu¿��L~rJv���D$�Nƽ�o׌O=���v	څH�Tg����p�r���+��0���k�g<��G�ۈDk����7�<�mڎU�������d���˧����Y��!wP�t����b_e׏����AN�(mq��W����)!Y��s'�r�"e��v�U�VA�h��\Ƚ�/�$������P'aL��n��� �b�}T������	���$8�O">eo�Z_��2�W���U!�@��S�-E:mž�C.�럷e���*��ڐ�D��O��܀�_&�����:��$�d��Q���܌�����z�8���r�~�����4uR�7_�dM�q�b��*�2&��zsp.����3"�nC�����[��7�O�~0={!�d�Sё��AZ�e<p����&>�Q��E3Қ��!TZ]��)'!W�n����<lv��1
9�z��~Z���Sr�����.�9�[?l`�;���s�^��V����Sw��0O%���&W�& g&�g���۸
FNšD���v��l�>#�:,��u�M�ړ���R���lM�*�&;�'�Y3���c��~�6]n���)g*��r]�d���! ��#��Z��-Ƚ3{�d&���[��|D=��ID�*�Ҩ�>ֲ���nѨ�i�B��~���WIɫ��f�*i+.0�]������mZ�A����J��<�T�E����������*x2�0V�B���0   �  B  �i  $�  @�  �  j�  ��  ��  � K h���w<j��q{�̔�Q��g�U2����!eo�{dD%ıgdό�e�=#�K�����\�~?��
��C�o4���*^�}��ӗ�V L��K��hH4�׻+w��Ka̯n}-�M\G
���������0&�G@�T������P�4�`G� ce�s�ݳ�>V�ZJ(Ԉ��e�>���J��!�A%���e����dXcFߟ���2N_��F���}̵P]:�3?�U
�G�`O��X����W�b�S�q�/��C�|Jp���V>�Y��q���0�~�M`^�/aDՍ�"��@�#��������d�����+1��>�0�@���!g��JQ[=u����T��b��S�d���ãr�
ױ��F�����I�2y7�wc�o�|T���\{���"�N���E�X���-�V|7G��P�=K���Y����0��5��F��(�a,�m�V���*&�oB	��_�
�P&K���>0�Z?,��'![�| c����p�V(��&�rp�?���X����{o8�����K��ݒ�	cƗ.~�MT����Wz�8'R�K
c�����L��g����I��ˀ�����h{��.��!	]:/ӝ`�:�q��Z�D��>2б�<��ƶiw�5��>Au
��8�N�3c_$��ԷP�
����`*�����v�(I�� ��� �'+�ok7ka��D[gG�G��K�}"��SU�P�����$]*��p�,���g��"n��0��I�#�\��%
c�#����(�^�ϝ�K������T{�i7�D8�ї�8Zx`̂qѐ�yM١�I�q�y�
�2˗v6��>k�Z R������M�X�I�#���h٩>��0fնf���/F;�7��Gtc�V�%9[�*�	n�0,!O�߷܁1�f��k�z�?�߻12c�N��h���7���"uq˾�15��5�o��W��*4�վD��X[����$��Ԭl7?͙���X�n���#��O�������.q���-����{����UÚ`l�/ju���K�]��C�o�Ϫ`̕��� BР�o=�%��w�raLQ���!&}4.�?���x�ݿ��^u�C�����邸(0���r-W�˞����2J��!�
�i=C�����*���ʖ�8c��8���.�]i�w���s~����@���i�4�cE�a��_�e����xTc�ԱZyN}����2,�x����8�����[0�WL�桋>����T:�5�{��
��[�.��j����u�N�ϕ/`�F�b�z-����&w�kŀ�0��p5!b06Ĺ�}�Qr8A�����S7��y�g.-w�;���^�c4��r����o�]|����aLcI%%b�c��gF�k�E��0�s'z����a�9��)\m�F��l諨^9¡���GPQ�	cŴ��껯,v��eT�Ձ�����ۤ�j-?����ῆ��rNbs�8'^(f�L&��D���|3c=C�]�z�U�فL6�;H<0�'ZF�ER���*�E���t$&���5H̉`I*[�����N�6��'y��D߼�T�# �x�	�jq����0��"?D���PLVa�ب�ЎQg�M$҃�1�v�$M����x�us#�;�����'q]2Ek@fy��L��Ot�.Mz'P���c�`�E1��݀�JƁ�B�M��{�m�r2�ald�y>.�ԝPuZ����39o�a,���R�
)��<���%�l�#��r_�m�j�h���54�̼ci�k���/&�ި�A�!eZ��6c��\�5\�����E�.��c�t҅<�����Xƞ�ϫ�d����'�R{����p�tDd�`��f)�c��\��kT�V�])�0a[E}=c'��a��?���(����dfP��'�X�-�ص�TO��=��^_%G�f�_��X�9�BO�f�ϊ�vT%n�y0�%2$$�=�쟔z�L�J��c&��D�Z��²9�p׏�~������.������>�2~󡙷�1���Z��U���	�K�Ual�9��᪗�������[��Ά0�w0j��Y�y`��x��%�9Sm��`�?��'��fYa�����㯰M,�R�R�7��d���x���4��y���q�l���[�h�+׭E��ַ�e�Đ~�􇱾�T����,�M�,q��4�5[�!n��b��6TW!B��NL�Ď6���B���L�I�Ha��X(�^��Ǆ����g�),�'�L9��_ğM���Ѣc�Iջ�%������rX�����ae�W=窯��ȿ˧�"�o��W&�DT�y�*�9�����Õ]0��p4���{��Q)��]��%[*��4rq+��6��N��S��1o�U�L���e�	g��~�q.#���τ⦹���Z�<�U�v�]s��yg�~q"glg���eH+�]R1����9����5[�/�c�W��H1��CG	9Q�6f+��`,��:{�F�v�ug�Ĥ�Mw�S��MM%�/al61ђ�)ߪ�H�1��Wf�/ܑp�ve��Z8mFaL��6v}�p�Q���狑z�EU0�N�t�03����CC��m��_`̭`M�R��R��Ò��O��f+:��װ״��2ڲYڐcn�1JJ��Cם�؋����k��c:7�קl�}�����G��I�Ø���㡱�IO��U_��m>T��)�sxb6~����Ş��s�C��E]�C�ʈ(�>*�a%���ٿ�N,#�m7Je���w� �bM}��ԉ�,қ�3{�`�}b�η]S��ʓ(֏1f,���0���j�a�yHc�3�*�&�1�:*�`t]si�ߪP��m��ǰk�����:Ge�k�b�V7�*�g�k��[C��&�\ܿ�*w���5��eڗ_���lU'g��'�Іo�������?[���:�.CMpV_Juz鳺;\2+ȃ�S���[T8�[�?�@�#�ħ��o�o�Y	VZ�����Sc-�����\r�F�#0b�)����ƳM��չ��9>��<��[�1�iM�w�E��z��K�3K~�1[�����7f1��*�B�Ҥի�����wӈ�:*gӫ��%�8���E>�}`X�f;�',��Z�Gh�=��_��7v�k[�x�oz���5����o���ݛPF�\�^Y��*�l�#������?Vn���@p��ES@7
c�U�NV�r�+�)Ƚ7��������u���M��G���`��8n���i���bQE�>D�"1��c���{	�5$�}{�p�,�`,�����}c��y�7������0���m�!*˻/|A������o�;|�u|���ڳw;�ؗ���`Luvq^���{ʞOE8�S��E�>0��^��>�B�ϭ����ڗɽ�0&��k�h��1E�g�1Ii_zO��v���x�;��?��k�XcB{����N�S�撨�1[���~0V�ON��b�Y2���ÚD��Ɩ�D������J��"L�p���ܘj�[��2����^o�R�X�F<�uX��@)�t��Q��:����Ч��0�,~� L��� Rχ1�˼��:�,\C9�ƞMKl��0v+�(� �혎�fD�
mU/� �y˜W��b�k|��n�Ѕaۜ��-歖����*���*���W�ڥk��^�P"��xn,�H���["�*r�,9O!:�e{�[�nߩ�mU�eA�n|��3k�X�4_�O~:�=�����䋧�c����Ju������W2��΁��:�[�_f�f��Ze|KK˰���>��>E�V�9F��Z������؆1>����S�^��|s{���,��m�C�e���F�yT�r0�1 n���`��?ףF�
��1�ơ�)���!��<*	b�9W�f�����+"��$q&W?���P�0%����P���_v冬-T�0�L&җ���DJ���h�&�r��������h2Ff���f�$z�[�c��1�����S�N?j�sH�RcD�w�F��o���ܚ�V�v�����r�Cz&u�_���4�5���#N1���k��S�:b|J\^�ӂ�JU1-�H��=r��KL�F�D
0&�	i�f���g�J���"�}QSչ��4�Ck���b�T)Y5�M��+=�R.��hI��)�<�\c5���B��Grfc~�uL>��(}c�������"�h��$���g#�a�0�f\Yl�5���?ƃ� �@[�MB�}�*��ƍ��/`lC���6ۉ_�0��r�M�ŗ�0V�/�y$%\��-w� M��!�0��q�0��-�Y���������� �F��%`2�6�9�F L��U�M'"(sk�A~|��Ǫ����fL �F`���q{d.��9���Q{I	���:�c>`������ �	l�20:`F�D�M+=��㬟"3�¨��t�oAkFl0;`����S�
��s��+¬;M/3U9\�q}�.�3����t`*�<��C���
�:������(Km{����� 3��)0E`F������㸵�g�!S����'�A� �)�F`��qsV��C`������d�tS�����	�L�i�n$���,X���l��[�����~�Ã�� %'㹬�Nks�D`��� ��,�,`J��E��"*��y��˂�'�q�"��4�+`�� +,�?0G`��"��H�{��XR�����/CR����"`���q� V�0*`"�����m����y��Tz���(lX8�X`n���� ��/�)/�����d���7S�N��ׁ�6 �)0i`~�h�M/� � &���Z���+����g�ׅ]�OX����~�E�k�k��/�eƂy�)b��GՎ-���W(b��0���,1g������e�d����`<~��`׀ŏ5F���6��N+	t���?	���6������h̹�9����=5����D����\���y���;b�c��|j*�$��~:#���q�X�"z�����|^�q�v�ñy��َy�����wڎ��q�nM=������^���6wlfV�p�v�Ǝ;S`��"��z��vú�d鹑/�[�u��W��ݍ�`c��`�ה�t��2z�$�^���ȟ�04`O�M��:i�.����q�>{��#ߙ�����K�%	�!`�9�%��� ��wG�I�p�W�ɘ���S�gC�S�;�^`�_�v����	o�w�
��E,&`7�Ol���ڴKn�aǯ�Dn�ǁՑ�Da6kn�i �̱u�V		��T�����w!d���-B�8����\��ؕU�F��)��q��50'`������{fW���D�w�ᬮ�Yw˩�;��0v`���t�x��:
Ȱ�_�c[�Wz�W@vbπ� s?cg�7�e8��c�?}k�zU�p� u�!�]�`���8�e(gl��~���8����&ݖt��U�I�'sq8�#`1�۱8֏*�0'
�ɜ���c�%nU��at�'v�.�x`*Wü���_{�\n�*+ ��uv�k��C�m����҅����3�2x�z��mn�=��\?�CE����ױm�K��&ͯZy��B_��rQԤ�`�X0c`�C'���3�n�9cr����\�����4o�!����0�w��b�\�v��On&5X���-�>i\��7��G����I����H{�Xܩ��a\��	��'�#T΅oe	�i�'��3�����rm��p�H�b�W�rg�����vb����՟���u��&͹�qgԘ4�-�"!������w�;�w��qǤ��Ş���E�y�SPk�Ds�h��s�73 ���7���ש-J��0?�5�isO��O�%lU��'���&O-)zU���;������_/�;��+�"���~45	=5���z��~[��O�{g/�}O��U��s��k\��#"�y����Fpj��`�n|Uy-60�e�OB��'o$b=�~ ���GG�'�2���&��U�i�i�.Q�pg���ڟ)��<;���}�O���D���G�E�?;6W�û�Q��K>��S�c7x�.���Bǃ�c�%���]����k�	l�{�5��I�IV���m�a�Ꙕ�aE
'vX$��3漷����T��j�{�ß(�&��YY���C�'�	��:�%!|�eN��w�P�K�������<���h��3`b�Z���M7�WO�;�U"̯�"l���A�J7R`a'������w�v�rF�]�|���=c��'W~!�����+�X�ݒ��H��v�gPNB�k.��փ�J����S�$|�]lf�y��q7 X�M`���/*�î}���p������a�S�R<1`|�ց���x��巠�?!�<+���,Oe��VƉrb&���!����'��r`RPu5�u�L댸��:F8+���~[��4�G�K���Y�Z�G3��*�c4ާ�.uy�G���������츋:��['� l׃h�"��3��f���E:x�k؍���?���"�1;~=�Ō^�O?�z�=�=�@�A��ݣ������&O��.� �Wq�{���ZElh�m�w8V܀q"�lEI"{dgDY�!IFDRD����*d$dF���&{EDfFvFIE��t��^�}�߿��%�f�&[ȷ	�]Q?��.!JN�2��:�4�.0e�Y���#E�R�����4��-
���vL��j4���2�1�Y��Mm� }����qؗ��ԃRx��,�#��ce�y���֩��X��<�Ha��� ɪ��`j��}�50g
A�c& &v�X��V�+$�&I��I��5���R��3kE�������bU\�][��^�yZa���z�<#�d�v������+^��-�ظmު��[�_����kV��mq�fH�E���F1�WmX.^X�5����G���%�6�%07070|w3�&�GuF��Li�tJ��<s�1g��`�?��v�O���\�E�S��\[�v7*�<p���՟`;��~Q.��$؎~�k#n�:v̲%����r�eJt�J�{쿮�f�`�``�`~`��2�n��Vg���G���(SSG���-�m�A-
�C`���
,Fx�,����d2��h���r�jdН^0=��8�w1MO���G �.��U�b'A����J��.�6������`�3�g8c��f�J�����[۫�l��Q(z�&�	&ƌ�~Ԏ�1�%�}{�-�?EE0�!`���j����KD�����%��?Td�K5;Ho��̥1�Q�'#�`tv���.��2x�q��ώ��6���1|����5K/���9���A�h0S��7`��9����۟|z�����ʷY���b�Z0�,����9&���"2�5����a�N�%_L���B�����у]��l�%áiOK���xi��C��I��^��KnS]��f�/l�� �=`��D�������f�<�C'M�����m�gy3�P�"0�3"���M�ߐ�mg�l)����zH����07"�w���~�6x]ɫ��$���,@��q���A$�o�.�7��{�Y���>{�kRm�/�fy���8��]�0�]`[�z��N3�IԆ�x�c;J-Ҙ��f�t��#�fQn����KQ[ KsʒN�R�hl(���q4��������h]H�s�Ѳ-�}%]���n�k�9�%v&�]�|tEm�÷)��1Q0G0'0o�K`�`�D�Nɂ���i?/~-���8��"%�k02��#���,�w�ξ��,�vX}~�f�
�Өʅe��cC:;�I~�y[�-�ֳ�ܴ~��z����p��Cš�?�婞��v̐n����"n�R�YC��w�D�\��s�+��c:5E̸���n�{��m�4?8�<�X-!���n�)�3*�Z��>R����Q9��S�j\ư:<�t7w�w�fH�a1�{�g��ٍ�ƃj���o��i�y���L���N��_���f7�L_�����ׁ�"�e��3>���ك��S������,N�ȼP��\5�y�PC�\��̓``�ݟ��j`&X��TVb�ؿ.3�(Ὕuσ�̨��4�v�P��Xf����\����ɀ�ǺCW?�1}�7�&=��L���v����5?��`�`\���}��{!��R��2����������T�%�+$��/�}M���y�Q�3����Ե��"����e�%��:�b1�v�z�>SQ���-�!o�K)b�m<b��F����E`��5!�h0V0���г;�d\��E�(�^�Y�j�`N`�8�X�U���u��ў롺柙�7������.i�`��'pݻ�`�',�����3��hu�a���[����%�X+؍��.��u$��vQk�ں��H��y�ĪV8��1�F{I+�yrg��Ywv�'=w��ʤ��㟑���6�!I�8w��`�l�&T�Ѝd',�ҽ<@WB:�M��ደ��\"��1C�{`�����
�R��=�c+��-�I�ʏ�-��K���Y<Q�YQ�!~p��R�@�����A�JoQ��ۏ3|7i�в��G���b�����k��_�˭�ԌK	���+��L�Tg�I���t �NС�CqO�����[5<������Y�!�f3�I����γ�����&��5���Pd�����D&8�#�1#�>�L�)g�V!=	�$-�7�K�L�!�A�su;#h�,��:mx��Y'>����ܶA]{�����WG�z�>��9��� �#��/Ug�w�d'r�I=:Ӫl�����H��僥f$rE�,˵���3��;��Ѱ�yE�����`�`H�To����	��5����k����[9k
���Ϛ��v���g�8��l
�+�W��`���E�}_�d�H�[F��Y�W�h�R���F��b�UV�r{�����+�����<�;`�`�8#t�w�|��y~�����)��F'���>�J����	�tG������U�z�*��EW��>���AXX�>��`���������v�<����-�E��n���1���������$���(�z�u\uLj98��X��.D%a3f��sѽ=;�=�`�I�����ߎ�.w��Qn��o�5{����DL�=`M``�`_�d�2�n4��\�(�����w����lɨu�����}�u`ۛ�ِ�&��y����\�I�w���;�3|7�Q�}(x�1K����j[\H���c�����^FLDMʅ&���6g��!�"�+Ճ�<��d��9�9]�E�\N��
&�F��dj�`�`a`!��A2�v>���HN�b̙��EdSܨ��[ÙG���%����������x,�q�<ͭ.J��ՒR�n��G�IO��&n{��Wj\N�r�߻R�LyL�3Xf�]��m�����_�]ɳ.������X6�T~���!��%�E-�t���F=:�q�O�]�{�7>ૺ4E�tƻt"��:�,v�U�Siۗ}��A.��wY �z1C:=�P��``9`���ǵE��o�~���Ԫ�r�S���cv���;�����ɼ��1U�+�GR�]�����Lg���oui������1I{;jjJ7���R�Z�C��ҥ�^�R�k8������{O%�DM�_�f\�5�,R��;�v�|1�É��T�1��#��k�������m� ӗϠ$'��#��]��D���%�mߓJ��.l�B�`���0á>�m'F�`�Y�,t[���:3x]izxծ�KL�4�]ؒ/xǘ3�3`�`�`�`����6�:a������N�zb~��s8��������čPC�w`ab~28c}Ic�s{!�:*4�e�é���R6�����!����~��PN���i�`�9�Xc�-:72�),��R��z�&�?���8̆�����
�r��2
�;zd'�2? �.|�]��[0R�r̔�P#+��u��_Q>��p�z ��c�
�L�Q;V �3B�B�Z��đ�O�31����F�idȘJ.};<�g}`H7�]l�4gA�5#���=�!�g�]�����]�`�`I`�`{���y�J�4#�E��:H��u�HN�y�9��!�3]�"�I"��C-L��ݾ�����ҡ���'��I���\�n&XlScUQRtMO(0��'��3�Mxi�Yհ/x�w�N�0;�Lll/���&�6��z+���J}���Kv��p)j/�����fqb-5S�[��~>�ͱ����f8
���d� ���5	�"#=k�X��_z�a��W&��f��'i6��G,��e�q�{$-8����ԬEtbE[�.P�-��+�#�k���p&j�`�`�����+K9��TyZ���	�[�z�OdG�Q�66�3aތ�����K��c��va�_�`��~��)8,u⻗�'��E�.J�O�(�:ȴ��^���}P�������?:���º�b�{�c�8k�J���~=Q��0������1���'2�m���g��|��f��'��7�{
V���R㕙Lq�-��
�r�.�_P�[[o圁pt]�&e쎓��8+��� �	l�خM��y�K_�֬S7yOY�P�bVӅ��X�7\�X�@�	&���ffU�[?�XKwB�L�g��O���U��h'���2�E��;��Ct��k��B�d�PC��]8s�섑�m�GSw�����f_�+-9XXX �Ƭ<5%0q��UY�c��>].�C��`���D6��G�i�.I�zyT���q�a{gyh�c�V���7��7�&E].�����}i�����'ҵ�~Ry:��&��`;�b������u�*���vٺw��e��>rEl��j����}�!�3W/�3�]Mw��.��Xu\�W�mtg`'��NC�����3�ܽ���<�!��s���ז��*V)���`�uLpF��i�y�c����}~A9�_�JR���I�!�y�r�Q�;�����wZ�}��N>�?do�������SQ� �s��ӷ�j	$_�d�v�rx��e����>-�$F�j�>�bI����8۽3�(^K�b�àQWs�Bc�5Q��:��`�`��:f\r�Emý�c%!*�T��Nf����M�)��9�#2?'�^��8�e暼&��X�����wW���`/�����bp�#Xf.�k����2�����\)���b�}{�ttߐ�DL300W0'�a�s`�X�I��{&�bB��q�ӍrR�
˚b�� �� �"�����e�浍��Ƞ����u۲G����~��e�F�\j��G�����R�� ����8���"���t;�k��,�-`�`<��z�u���zTu�ӕ��E�U00�W`{0c�@-l?�9ؕ��RыӪ�E|��G�G�ٶJ�~��y��玨��"#���j���������U��{�=���tż��I����l~'�����~F��^y�]0e��`T`<`,��O��f��O)����뻌M\���jI`�`�%S2��y9��}(�&X��K��~t��D?B�����Q�R����u����ב$ߩ��.��1����ԟ���>�8���
�������X��JL�w(���z}��f�tO����}�B��o0R�\��*b������W|}�*��\y�Q{�3|'���^Q����حV��)��I�iWE�	�<A��ʀ��������O�z�Y����P55m=��&V� &	�t;1�G�%��o�%aҊ2���������+�$������FVݻb�������=�܍k�w�D>�b��&G0[=�樁����[��ڙ�}�y5��77>�ܦ��XX>X-�(�"X�/��I��EI}/M���s'��y��	9�� �s��ҝ��e�yg^
�^W"L�S�9�D?%W[	ę��KJ��T���[�b�����dg^���)߻���b�A���X~�a&X$fHW�X)�\�߯G�5��D�Z����$P�%�1��av65z�]`�`VX��p���A5Ŋ�G�.��~� v�j�`Q`�8C:Y0��ۂ�%,~0��9�����wͺ[�wokXH��3�\I��н_L���ęgN��de*���tԛ���>� +�� �w��3�$�W[��4	����j��q댹`�4�����ގ��y=jM`���=�>Ξ��h��f�(�Wv����[܆vSkd���4t7��3P��l��p�d��]֧o�eDpT �3�B�=``����&��@f��������?��bp?�W8�%�N06�}��,��ѽ�;�Q��8w4�=�Fp3q����t:�E��8�w��P�kL��G�]���my{��e�GUCV���\�K>T��Ϟ�l �t�.0)5�����<��-<i�Wm�$#��憙h4j~`�`�`��u3���+|�&�.��!;Λ����PkKS��޾�3
�ae�dQ�����T�'X��t�]�.��g�����`J�`6��>������t�:�!�s��6�X �0a���!�UA7���E�;��(w~���c�5�P0*��Cn�D���C^^[�J�X�_5|�m`W�ƂX2X=X3��.C^�kѾp�b� ���j�?D�-�6$5�&�S��و�Ә!�0g0�I�1�¡�h��÷�����X���L��:�O`��H����ť��g�ʹ�纝Uٶ�n�.��YF�l;X;��3Y[��e���֫��J���g�*]�~׺,���D�N�����g/1qJ|2�p1��p�������R�w`�`�`.`H7���K��+����S�ђ�B�Cs��OQr'U�	-i!����i�񂕁5�\���^f�{Y���v;_�۳Ƣ`��ފ㏒}������k��)�}�:r�*��s��E�6���&��	��O�6�6�}���񋮭�<����`�`�`�k�!X���qֻ!�&g�$�����yV<�>���y���!��t��\��� ������ˈ�</����9��O8�t9�p��I�E���i��0���Y�8�P��.���m��n�r�Pk ����:�t]뭆�=��ׅJ×WM���jq`]DF�����3o��|��sM��-��w?����C�L���!��p�P�Z�ݪ>��m�θG�r�f����V���e�4���`*`��f���K����Ty�j��j��}�wn �Y��`�m���8��Њ�>���r$LYA�i)�����_͂��g]XK�b`�L1A^�!Ѕ�;��]i{�b\�D�BSh�#��c��`��&6 V�u�7�FpF��˭��On������&f�`�D��Z'���k�=}mt�����l�5ϵF�I��	�Ứ<E
�k�Ɉ�	}�������G�*O9�l"�~���wI0�J�9aF����@^�AGn���2��]"��5�H�c`���1K�D��0�I��E���DJyn2q��� �j�ȺbP������5����,Y!vsz:O��%'�	�K��ڿ���Z���ulY`K��`;=�D������#����ڼ=�l��l��?:*�O.�]f?Ŵ�HYj
|Ȳ�3 6r5s�loD�����a����G��)�����"�&�|Eը��L��ly��$�8kӉ��4�=o�0�z!��tt�g�1C:m�s`1`C`�&+E��X>�Y,s=7�s��g�o5��Fm���5�k �w�xLW�/���h3k�}}�Si�P�c��K��jݾK�"@�������K��U�%�ڔw	���T����{��g*�}Mԛ���e_�ừ�.^_�Z�F�	&�t�ij������(݊��V�5n�N���s��cZQW%��t�Ƀ}�
��x�[߮�KL�Ȳ�w��������%Xk�y��e�}�p]$�ݢW��W��\�9��سE_e�,1>�K`u`����uT5,�{E��=��Y�6��c�
6�˴3��پA���w����`j`�w>��i�u�qc��������(k�1��/�%�6��9���\��E��3]��`N`�`»Ǯ/��1��Z�l59cRu ,��^C�^�9���a�鵄U_�ږ��ҦZ���|�A������̀y����s1U^l�T0���	͘+Xw�r��	�&ҹu~�>�����c�&vڊF�?.t�+�̌�%���-�Y��V�_�ػC�M��K���9k}�e�i���l7� 2�I�L�.��h�10r��g�Rf�6L�m� �>����Q���n:K�����A����ʞ��1c�/��e�5��bf���	�#X֩�bMr�Peȣ��0,�i���4��>X X�I\w�ي�y��v���2<"1�f皮�)�l79X���9{�gI�����P�����cH���*j�r[R7~�L��DXgi�!�0ڗ�i37��S�le��Oɦ)�� ��v�8�t���$�Jƿ��>c3��ugqs�����
"{���7	�W����K��l��?��E,�_��Y�%��،�=�۝�>���G�	����ڗ��q~�)��Oy���NdR�`_��m��S���,�Tu�&�yua�����"c;�F��J�և�Ru�'�!�̹r�s	M_��m�_���)b�`�`B`���y2�(	&�����7��r�̈́ҥ��!�Ov�?�tbs��p&��}�c��{�X�@���9��?�鯯�|���j}`�`{�܉�O�>�v�6)�!R��mz+M^��-j_���Q��](��zn����pǴ�^�mS�����8���"���!��U���v`�߳=K^��c�4��&��Y!�`
`a`�j����$m���Uz��k>Xg(�$���u��,[���PJd�PK#+;��V��9?ݹ�hփL���2I���>��#�dW@��Wٿ�ש����ps@N�ְ�⋣!aE'%(m�����l	3|�2'ة��xD�g��7	";s�z���
jQC�O`��~&T଍���0�#�]���ō+;��p& ���>���,PF�VzΞ�����E�̘�{�j3�������g�!]XX9%g�I�}=���}�;Ҏ�o3[��<�s���`]�8-�@��l�����IúC�|�I)��F&�3BWҜ����z0��G㍿/N�l����ym��M���;C�W5�w�pֺ�\���^�D�ҍo���j>K?���w���s��8
�s<�H���d����S�򈉂)���Z�Y4j�`���c��$.�&qLb��5$�m�+;��fӾ�`e��.���u�1Kk3��f�po]"Y�0i���f�`����n���[�:q��[]H�F�d���{���a �Cm��(�4�3��À����ǳ�t\jO�Xݔ�s����0r�[8�w����G��c��[��a��U�h���z�Ƨ�1�!U���,g&��)��^ܛn�� +�_YvR�V� ���W`'�v���Ebv�5/��`�`�nr��[����jFt�z���ds�'�}wFm���6�l��v\:�s�����=�V���?�yFT&�5�����͵�k�痄���W��4�4����� ����/0��?*��NJgu<{{W���^}g� [�t�(���x@dțT�kh�w��E����u���=�X<��5�2�g�}Żl	vU��.��;tlC��x�Oi�U{�G����q�
�YfA`}`�`q`�`�`k-�$�'���]m�4iο�P1f6m�̀�����u2���W��n=K�5�{���O���=��3|���M�-<v�Nc���{���؉���Mf��Cɘ���Md���g_q��Y���{����R��H��Xv���;v��0�E�>Xq����kD�B��X�s�޼�;.%`a-SD&�3�8f��1���1�2��9x/�̒>�^�tHo*�|��,��6������U^�gt�^�cɽ��cK]֓��1�M�����]�{G�������z�+��_�c�����A�J�(�t�,�Pu�ռǠ��%�Ən����Ǚ��Y/vO\��I����:f7��_Q�ޫ�����֋��������0C�n�z�y���;W[s���u��V�9��q~>,��M��������N�{��_"��n�4O��cg��̇��`�`K8#tT�
�7;�VZ2�ud�)�5�S�)������J�~�!������A8�x�in�I�?�=u��5�_����8��1�$0|W����L����Z�֔�d��w�mr��F̞q��/j�`a:+���>4p��}�j�4�f��$�W�	6r!��#tU�0��ض>��5��E���2������,�	�9��V�:0O�Kxy�TL$7�������;�)�ġv,�,ץ�E(#/��c��!)L�SPP�n����%��I��v��fe������h���w<���q;��([��{S�-�leU��!)[d�=��
	�d����Pd$;��t�\�\�}������9�:�:H.���ˑ�W�]��}:k �Ib��&��e�8�� �����y��s0޿�,@�8/�E���l�9�6�b�Th�� ��{�p˴���	<���{�{r%w�MO��I�]b79�񿯐�^݃?s�"h��w�^��v䠀F���F!����&F���(�'83��<8��1��[s����n9y���ۏ��%�R�V(x��=�B�S�t���ɓ/vj��'+�H[�w����b�=+�X?����L!R�=�'�a�^(���M@�(���q�7�_N�$\-��Ε$�~�Gե�������Cc�Ч�6�v%��	��T��y)��+�)� �&Fg���T�9;1�Sƣu|�DF��	^l�}�{�a�ݐ��^-M�A��ѵK�w�`�ˎ�TP޶�z�l�YI`��f�[�����̆��x\\<�ۄ���6����P�2b�th;�럵�o~�� >o����A�[5(�6�~�k��3G�0��`���Fy��/|aϬ׋ν0p3~�gb���rH+�c��󂭆ӷ}�~�/���#���>�%�ł���[����}�Ʉ}�Q�V �3^����_n>�#X:!��"6 �ՙ�a�����¯�Y��+�D���j�m���p�6�l��7�J���Jm�x�(�d� v8$��� �s��g$���|��hs`�I�1��O0A0i��/�ML,�������)xn���O�����۶����	��.Cus`�-7zDM�<�æ<.��ˆw����捎���=txi{3���Z;M�B�n9�\gQR��Χ0�<����pL����#G���-��S���3���NQk(Xb߷A�E��3�
w�gj����3�6�-��$�5�v�R�~e��u�10ޅ�9۩���6�}9�Zb�g�݈������LSDu���YW�Ϛ=�(�G��
�-�w0i0�Z�;��/��[�\�U��r�\��Do�ML�	��CY�*��V�SG=���������ŚXe�`�`_1����y��E�2�[�ñq���h��3�x���F�]l]3+rz�<%�DՑ���3f$̏��T��^��	�h��
�&�V���8ڸ�����MY=�6���=��}�����l�m�``��pP�s��5���k׬��&�=�v|��5��DP!پ�N�xlϊ#�����|��\��ǯ�P�m�~v�	X�4���?t�,˪+�]�ɎI<�b~ʌ����͂�TUW�2��-t�miⱺ�O����	�5�Qf6	v��0�]��mKb'������D���o�r�{5�Av�g�r[ ��[���X�'�������/�ڮ�DM.��|F��070_���_'ۻ[��M��D�>}�;Fb���O`�`0�#�=,�Z��k��D��aI�7��5��8	۶����Lݖ�`�$bBL/䥓ռ�F��)�ʯu�s�ق����́�:�.ӣM�Ȫxƃ/��=��N��n��YoM��9�G�2W>��5 ƑMr����תZ�іU�N�<�y�Z϶mMy��9s/t�8�l}�9q�LjhV�4�f�u�:ze�`y`K`r`�`B`owu�t!E�%���]�|"����,54���i�`F�v�ֿ·�a	f*r�-)��77�����90�,1�,b��7b�-��W�-����{!Q1nY�G�j�|&��ߩ0�:bG�l������f�Ŗ�^�<Y��k;����,�,�>b�Ih[�� ��t�^_�H��F�LraSx����F�ms'B�"���Ʀ���SX�a}x{�bU�Y�O���OJi�E�>`�G��<eز�&�G>Vlu})a�h��|��0b��`�`+`�]?b�7������˵NQ�rU�[�^�T	=��d0*0ᳱWJw�mk�m��\ԋW_5�dvO5VА&��|cގ��5A.N��m�X���pˀN�<�����+�UK��ˌ��W՟��E�bF`�`�`8`�`�`�H'{�J(�G���@�Q�LO����h�#c�����E�6<�ڮ����|�>�IاoߗG�L�``���uUz�acj(FY�q
��Y��x�[.���̾qj�,�.7N{e�ꤿg�ű�B�,�����?�$_�Q�dP&�Q0Mv���s�N�xR��q�S�G>�,���wj��c��ӥZ�d�x����$=l�;F+Q��l%H<o!��{b��C�B�^͚�<�T\	���N*�\�+k�G�6g���/���$Z�Zg)Wm������9:��Q���\`Mt���W���,��I�SF��-�k�<rRy���8�74��
�{퀯]�<��Y�BO��?�l!�Xyʴö�L�.lf����sI0YE�%�&��t��1���b#��|4u=2������1�-X9�N���&")�ac���ˎ��������Y"��`��� &�t4`7�΁�}��Q�,Sָ|-�f�lWǩ�������}V�8�
���G���:�SLQ<�foY4���g?>�B,l���z5�70f0�f�a�l�J&
�˿�M����Eksہ�:0=0�˱�滌��.s���*�&C�Ga�/��ߞZI�����PP
&��ƶ�6)�z�M�ڿ�|�r�ز�~��|{)�	ّ]淫kkk�$I��{f��E�n�MB�~?&�J%��`�`�`�Gі�X��-{�:ixc#e~��V����6T��\�u�*�;	���P�܌}�KQ`��+n�w�B#��r�``{�ж��0N3cם�s�e����-:�r��m��q�ݢ���,1k���`9u�b�5L;%f�^S�ZG��%U��9肶�d��0,L�۳&�{qI󍺮�k9\snIW�E��GbX5X=XF��꤆o�1U�h���8;�s�e0�8@j810e� ��}"t�|��.�8k|H��$5Cy�s���|��������t��l`9��������\7�P�Ջ��br�L�40R#K�ei���/;�Nu,�D1e��G���!�����K�i�M"6Ǌ�����ȶ��޶i�3ԗD=�^~��+���c�`~`?��:w���sv����!�p��=c't�2h{	?g�C������`Q``'�����B��7}��7�i�4S��_�����m��^�u��ˈ��
��������	�ʚ�q#���^� fFF
��m��E�3�5��Y%wWyw���S%�Ì���>Z�e��:]0]ۡ�L�
��ůk_>��%E>�)� [ ;���׈���2��[�Wz�J�a(�x�5@^x�O#S���0:0E����/��'�<AI�Д�@!�i�(���_��mw�v���+92f5�/��TO�+�prڱ`��ɂy�];�WTP>?)�a �o� N��;�VA�s;��3�g��)0�3�Ok�d��������RR`�kD����	��R@u�]���4�~��ua�$����ml�!��!������f}7��v��{.�� ��ω	�� ;��b�H��2eZڹx��4q%GH������(��]�	�1󍶊���0�R��z���Z�D�ՠ��HK�6��!�!�6#j+���}��
��#:D2�y�;& F�ص~b���qhU��V���$���
�Q��AhۇX-�3+��:Ĥ�^����憎?���}��~l���k#0���^�m;�����
�͔���gq�F8�<Ж�6&�	���v��w�%e�H�:�=�$V*x���Vh��^��m�;w�g:|6,]'�YV�)��9u�!�x��	����.�/[�H��]z>�Ѫ�{���b��_��n���;�eD�L�^�K�-vC��8�"︈*Z������Bw���=S���xn���xٽ�7�p��wL鼔նy�̓჉��q_�c���mqĭ0,��m����"ձ��F��ݭ��!Ȕ�.cw�Z��%2�����N�`���i�M#���խ�Ԕ^A��I�RFj�Y��tް�)M0y��]vl1��r
͂�dY�yn�=��=}�܇�|O#4����Vv�y����2>��0�szhRʒ�����!��g�s�`�v1TG��W�k�^�U�Y���Oݴ_��>���'��u"6	�0��сe����-���+��p�so���oȐ�߱�^�̀bt/�:��<��bw�+\�&֒�xP���Gb>`d��Ճ��сM%������>��s��2{#�zs�������}`Y`T�_�Q��T0�?:�K�Q.���)��1�6��}9Ɨ���S���������;�����K�����׉n|�ͼ��3<"{ޥ�����b������=b�'�� U���5��r2wlTYG�E�H��,������}[�K;�������_������X��w}�R��E����qxP��Q�E����>ۆ�h��!uq���a5�l:a�l;�X�,����X!j[��ln�_SE�ȏ��g�W�5�ж`좋�b�^�Հa����U~ȵ3�Lqo�"���֪"�QH�������"F�f
�{�j(���]���Q�G����2ϫ��-X,/X�b�.�Չ�y��7#�5�|��K�ǒ��E,�X���it�6x���o�o��\òh�q�/�ق]�Bյr�;q�V�֍�+�������Y�s���`ʈ���;�P!�d�F��Uc��z���҉b��nE�^__5��傝D�$%�S� c{K���vזJ[�ߪf���M�{�فU�-��0:��ê�:����X��^������ o�G�X��,��%���5���>��-?o8��WU#Hw�¬c��GM0��]x�(s���tIo�~X\�2�7!����lOz�6�#$F��Fxm��
ÍI�oΣ�?�P��DH����1ܐ4՚�����N�Q���3�P|\�Ը�-��?�kL�������y/�m�~��[�$nY�p�S�N����l�|����%��```����Q��)�q���Y��7<�s�K�O�\��!�h�ќ��80i��!��"b�����d����ؽ��sZy�a�.1�֑|6|<Ce�`�`���M�� ]���� �/�#�i2�5称�DZ�d�B
&��v�&��G,��ۦ񪷆�>�؂=�����7JΠ��L,��$g�߮4<_��<yA��|lh%~�${��$X��k0c�J���٧&Q]�8�۱x/�2�ӵ���w:&��H�X�n��U����t}�}%���'~`��}�h0�b8!��վ��ޓ���R������t��s8b>[֏s*C���3���	;}]e�pW?�.X�q���d�;U0�K`9����պ�Ը�|y�n䠘����\��q�̟�6'�T����Z�g����[5�Λ-̝��Fl,����(��S�h0� �Ӯ�a)?쐖`�����E���
��G`��(+�Bw(3����}�J��]��ժ�NB���v�9�r�s~��SӲC�b\�I3C_��|"���;Y��99�B����<��"���+	��Ⱥ�VC:gO}���Ӑ������`�`4`���@[b�`�[&��q�2g����X�l�ws�Y!!^��.A�v
&��~ls�0끻����N��CbՑ���7W
�(������U0Į���~�٥�%�/��0\Q^̼��n�6V�F�m�K� B,�������	}Woh�dQ^����z��c�Lk[G��X#���%�8:Ç_�^e:�`��0[��-�m``-`4`Cu�!�N���u�u�DǧEg.���4>����B��1K0s�n����c(���*�G(���W�J_`L���ݪ�0{�`�G`S��:Ct7@X�pZ����A��n�?{ė��B��100>�KO�������o�J�Ͱ���+�(�e��K�Bl[�3�f6�q�&޹�r��EN��Bog-�d�]����s��6N�luV�bG���+V6D��9���?�ʋX�k_p�10g�t�'��ƾ��}|��|G9�q[����FF�/�z���$U"��1�?�w�3�s%�Ď?z�ԧ���|&4A�8 F&���8���W\P`UK"��tι4Q�!˷���$;�e�6���KbM� N�f�<��tF#��k&�dy0v0}0�wvhcDL�e�t�;�%�ǉg���#�լ��F��`��}@�0<�e�>�W�����Eѯ�H�ԪTHη�|u�iQ�e��hkAl?Xb�'Q�˫�&��"�ͽ�Gl��j�����}���H�����~#�V�.�Q�{�j@�(��GV��U�v�Wh�E�,19�l0N0�^�F�q�dZXq�7�#�-ؼX�P&��v�L1T�����H?Qٰ�!��H�������+�\�l�Ss�+w@YΏ
����� m�_>�i�/G������v	1TW~m��ד�]�x��v�H��n�����ڣ`�6	6F�s�	��/�z�9߃�ⅺa@A�ǲ����%�3@l�e��;��l��>��êƢoZ�_tZX�zǎ�	���>�m��:�'���~#�JW��n1k�<y�9�TH���cs���m�B��?>k�y;h�[�ޑ�f!R� 0���^�1`X�]�MlC��3��m��S8��oz�{�m�y�;�X�5؝�k�7�q1�*X;~�C�xO�زwA���L�
ʴ0�lW�	&��2T����œycf�2�3�5-�,�Q�q�5�ݩ�1>���-+���d%�y��/"X��kػ��3���v��E"�V�Z���~��l�0�{��7T��E<�_�	�R�+°���"1BF��{�s���ՖmO��Lz�H�1~�$�s`�u�Þu1�M%<d)�;5�>�G�r?L�x�>�y�Y`�'�k`����Q���^U������I����`N������s����P��Ei����G�u�]�~�B�)X;X4������+�$�;)�ɡR�O�LI��J��S9�k�'��� ���Ӆ��t��W��*o犧�w��ߴd����ì�|�t�sdQ�����
�:��Mu 7�~���'����[��Z�p[����%���2�|�$�w�������~��ē�� �|�ks
�Ê�������.���%g�-��^tz�a��S��}��ߡ;g�7`�����m�|w@�A����(��͛���n`7�&��D��d0��N�>=H8�@O�I3,��٧w���3���T��E��5����iA��r�xA�ElKgf���4{�)�C�V�3�0�]];���!�9n��	�J'2sj���V~Ƈ�Q��K�ZݱS`u`�[&�]�3������گZ�s�T��i��Ex_b�YT� ��牖��Z͛p���lL2t�}7�o<�� �[f�1T��7��LO��=P�VT���?_��}��m��&{�f���W���ڶ5|ks���d�R͹Y5"�d5�6�����O�\uB��>���ck����d�3�N�sD�-�s��"�"�!�\M<�X���Sਆ�Ky����%��nO�{�5t�����?~h�2�M>���÷[/���6���s�n�F���OVܫ�t���b�S]3����!Q�&Թ� �x���#���d��#?��4��n<u&$ѻU.��*�]^����������z��%�v���a�]9Rfm�U}�4u���ͣ��Ûw��K=O��gcjm�p��x���p� �?�ufCe����l��UE��g��qݵ��@��*�x9C�.i�ؒ���Ii��7;%f�n�u�'X�D �NR��Q�I�7���y���F�H�f��$t`�`X���w�H����s9N����[�f@٥�������΢3@"+5Q�E����2s��|�I�G�pP>�.��;�C�eM27�nD��!�E��,��6�C2EX�L����z��!\�Ww�*x����ɦ4�?y|��~`v`9��åD���n2H8�;�TƚΙ0��|�gib��˽���ۓ�F�5�]o�ُ�w�{2sY�hO�2�,�>��at{0��:���3O��EC��ﱍ����7VZ�|{�Ƶ��1���T>a��gT���C���6�5�,4�Y�}=�'��N����l+��o`������^�N��A����G߭.�O/$m�'�!g����Ǚ�D�G[�9=}7�C��n��F��Y��-{�jƦ���i����4?�Üj�j+8�I^�������2���0Y����.�3��t`�+��
�,;����o���r[��}e���s8�Ic�3��n۝6bG��g]n��X�q��-���?Bc��(s
�Z�����{6����=�z�n���H9X������M�?�D^��L����nk�9�<;:�x�M��k7��ך<�q�!�/L��zIr��7�7��`�`�Z�SC�ܶ�������s4������ח?��'����A�lb����c��J~�����EW��f��Ͷ��L�mՈ��kS��ml��ͨ�����ZX�鑧�@�<X4��b��������0��]�!]�i��i�o8���S�kU��Κ�7�U��e���W>��GW�K‚�p�_��5�����O�����0O��]��{6�5��YĤ�^J��	uD����82���������Rs-蟑~��l�oǪY�|�I4�z�����EnI�A<��	G�J�K��b�x�F�>��]I���ȫ�<�����r��~�Lj/m�}�aǖ��ן�n6cr{D��3�`#"I�h:C���]⤙`�＝P�O��/s��S\��N�[�l����	�0�΃ك��l� �����@,�s(��]N�ɨI+RQ���}A���,^��{�Ԇ�P��m�^)QοY�(�%~���?t�_HWpV5hB��;�m�^�{
��l2���Q~�,L1T�
��)�|ɉ����Уy���.,���QfI|��{���fc�^��vO.�T����6�4�O�s�ȱ�<��P�Q�PXj�V+JXK���jntW89jR�X܌������߉�-X]�X�V�X-��4冞Eq=x��K^��"�)C���؝�c.�W����~�c��J˴�k똋)>�=@:k�(�	$Q[��3g��>�]��)�O��%��H�,1Tw �ե��JX�y�t4��wiUn͢���[��A�?�����LU$�V�#�r�&����G�S���t��K������L�����'�ZJˋ0:���!m�ݑ�lL�I��]�ݱ����u<������Nb�W���������r�OY
ŭ<<�Z�veQ��S~�Q"�;Ow��|�:X)�5M��*T�y�����*Kh�W� �e�}�K,`����iHW�# ��7���͊ژ������Y�Zi���\��F&�Z-?�4Ƥk�C]���o&��,�:�[�V}"�4Z��7�${��j���QU$�s��M�:�Jesڿ�q��_Vo�c�]����}�|"����nг����)�9F00K��(�a0-��u4Dr�b�y��	��M�.33�>�z	�Ӑn�Q�Hp�ԯ��Sh�G���P�P�(j����9�v���yW��YIy�����jc����S�����a3�϶V�f�C����f��%Kw=��?�Pw`y����wJ�-���݅d[{8?)��j�f/s���V���`L`lX�r'�����!v�����?��EE���D$�L;5г$�kz����FV��H��ai�ۭ.O�o&�:���.�9on��ԡ������]^	��NV��y�{l�������]�
�>7NS��/���Ֆ�{˃�����	"��B�����<���^	�Or!����qF�eh���eX��ha���6hE��;��N�A���Ci�E����;$����������y<J�J�lD�B,0�q�$$�:9�W���}3���;�V����*[H`�p�ʺ��3A|ͺ㺰��f�c���ˮ���J.,�q�y��	���և]��%������̋^!0����T�	Z\Q�䛜�?Za8����~���;���a0q���?V}n�0�c�f������ժH"��Ԉ<���հj��$�bU������+n
��Oo�^ڽx?�+�f��m���L�.,���u.�FS\;W;�[ꖬո�vOV.����.��� ��x��}�ޙ{�/2OI�M/d���e��bl廓~�i� �5Ic$q�A���
����b|$�.l�_:fߎ$ǫ����*zΩ�����˴�UۘM��p�����L#���?ǩ���0Mx6�
�tI�{�V��L��{anV�]sa�6}�y��G�n�.��6P�"�H#e5.������[��M�,�n�T�RD��?8�*��8�����[wa�;3'A�B�ݷKOk��o��h��]8񻰖��ߺc&�r!4����;�c�ˮt1W���VaY����y(b����{~���_��v�a���GSf�O���X�Ġlm�GH;{�%M�}�,�O��o�Irn,��$�:����7�� �!�.�[y~:���z��j��+�=�)�.��o"�g�#��A�&8.����\���HL��Da�5�0�I��K�"^����ý��ir�w�b������Q��h�S�39=�1i+o%��K�xJ�M���� �/~ϯ����z֟|�F��p��g�0�8�r�Z2k���<T�1�y/���q��]i�)R���@kboD!|ӫ�x��U�H�`x<LAL�W�۲,��:�Ψ�@~p͘�2t���:Itm-M����ͭ�G\gQ$�����x�#�!�GC f��]宦��[5��Ύ��3b����m0(8|���#o����D�!���������C�8��� &j��y(��a�D�*�0t�E��b�ߟ㏄�,����8�nb�X\e-tY#;Ev�h��M�]��;�-��5����Ჲ ��8b��^O�D^
?j'������; b9����\�e6\H��	^�z��{�j]-M7�H	S�*�S"�b��⛁��?�}9�g��5�L�h�N����k�4)��� ���J�M� �ů��w�����d�Ɗ�R��u��{|�s�1�S�v�N��3�)�^gsb�2t�C�F�B�a�}7��:�b$^����ڪy�{}���o:����{扶�����yo2�l��AL�Vzވ=3�@����~j��52��I���� �e��.�0�T��w1j����?%Կ7c?-df��1��+&Ų��NPw�R�}v�� ��3�a�L��QݾquH�M��E�"������n����y��-�J�4|Y/V�E�������1�����o섟7!��1���b�1�e�`I�#H>���.�S�u��B���{f0P����M��2[�K1�gx��1�� <�b��2K�1X��$��{~�9�J�7�ޓ�y���U���kaB�A�t����r F��'����Z��� �^˹�>�M��������P������p=7�tp�L��/Ōt���JӖؑ��� F��xdmX;�n\/%��{WA��o��f��;?�O�����D2���VS:�IȌ����ѻrt'b�/U��ߢF2�CW����uNqH�~gP�9b�ǚ%L���~a��^�nm�i|�g!&�u|�����"}�-$�QD�}��E�I���uݪ�nG&�<�������LW~���֢��rx�<�����RD�H�yD��©��}���X��'pA,�.���wt�#��v��'�L<�@L��l��l`��F��x��<L[ֹO����!�r�E����������Mǲ�X�D�w�rA�XO��� �!��|�)�U/	��Zg�&,�"e�5'�e�#5_òb�����r�L��6P�e<��FA����`�<6$�:cN<���w��v��jD�f�Jw���~�e�M.�%h�m4��U�C&+����[����֝d|��l�4��Ug�;�. �=!�EUR�a��v�F�=��^bv�8�Σ��?8���G��k˪�gt��p�~��~�5��'<��ߛ0>�M�;mDM�L�LN������җ��I�?��G�6y�)��+wL�ՙ�A�m(�G�2���p��(G����l��������qU�V��[��{-=)uc^5���d�B+N�$�;�N��"}o	'�Z�JL�5K.��2�I�����ϝ?Z�����zM�]���渜�;���aPߨ���5�R	�R�������	�X�hG���J�c 2��t_'���:�9!S�V�"F�"���5�1��Pw�'%�6��Ha�1��2��wue����&�>�{�Pq�Z�2�+R�4�jJ��A��Kw�V�sC[Ҭ#��ѣv�D{H�'��Κn0�%��|�f���v�5]�@��Ԫ=܉k戗��ܯv�-�=O2��|���'�1s��i�m<��v\Ħ	E��z�-R�!���s嶈�����!�î��w0N�`P���"���J�Ɇ�
���J�gf����-u���ᬜp���Gs�ǾvM�e�"�c2�}�#$���3 ����u��E�*?Ą�"�|al�))V�H�2�?�}�R�y��?�]~��Iu�����F���N%��$��	:X	t���7T[̱�,*}3q���d~�u�
x�A|aݦ���_�g�h��D՚����RO��ǭ��3C�Z9�X;G��(��<�dH��\���Iŭ�w���jq���h$ͤsQL����\B��b�QY?�^;֭�T]�R�h���ï��#x�&�2�X/�s�&G˼b�"/���j4P ks`6���з���4Ο8]!Ԃ��~�Ԃ�m/�2a���ar�O�_1�aV	l�d�1�w<��I����|d�@i�o�L+ǐ�6���d�*������/��M��d�%!��N����O�z����E�iyP�q��z�/V;E��$�V!��*T��Dg�d���-j�|����	Z*_�_�����Ph�,��dy������}�^~����{�w�%�wh�i�������z.�6g��۳>�=*��Q��q�6�*t��	��-�G�K��C�|�F���}��GK�6̟�n7s�����0L�Yg����]>���ԃU.�Mk�ywQ���"U�΋�U�K�ه={��M�tW��D�����O����,��K�)q⑯�40��ʅtMln8_��/U�8�f���ٟ1(�j�?�\y�Д��N��G#^�u�0>p}=�xr��,��,��W��} ΰP��e�ZK(���˞�m���ב�i�pCAn%�N�G�X��X��rү�[-��~�._��>��؝,��1����y�'f
A,��Q������i�+�<�n)2���f#CY�h���4�	�]��P�����'�~���e��CyN�f����㐅JĊ�����~H��c+��S�"������%h�۳�m.�XF4��̰I�G�;��Y_�~��*�? y�y-x]kp��62�����Lq�'��!���約�ӈ� 6�����>�V���I�7���\��|�L�c���S��u��SJ����]�9R�g��r�?�Stt�Kg�B9�(vep�,�9ٌ��I���F��˼��[cKRg_�T&���Ȉ��[9���o��h�j�����* �޲�R���g���=i;�g��_��Vh<s��~�Bg�0�d���wVv��M}�ة��7��J�� ON��cE�6옢�r���!�/�ݰ�6�c2�o������t/�.�7��nRG'�*�����Q��ݱp+�\���(o��1N#��&�Ėk�	k:*=ܤP���Y���d�5�a����v�w�3�gxK�f9�!O�QC�`��1#8�������5 �����u��<^���n������:嚾xH���m���ݏ蛣n���.��&Q�d����3�slĲӣ��Xi���+E�aV��4Wd�zh�&Y>~T�4�m����{۽�0�z��9�c��^��o�	ٽ|�A���q$)/��}���.�1��#�<cƍ�	�1d�[�t�o�u��Q2�5ՑډmsA|ƉvG~4x�$���ć|A7CySw�mj��Jף�{5{>���F���2i��am9�M�<xW�⺋�c��8�֖����[�\0���"��Rҧ_2NԸ!15^;�g���tf���B~��&�b�� �9˴�][�K�t��������N��}ÿ�)bxK�~� azP��pd�z��[�ԱX�3z�#�����+[�l{��]�ڱO��զ�,GM�*�\�Xh�i��y�݆^*��P�h$�����cE�0�!��'�<�b�/;��R�����v�Sy��'�:�i`v�ک#5J3xa�>3��"�,B��i��R;���u>j��Q������|�#5sa����KȋF�ޅAJV��&W��nĹ[,W�ѣn� �\��#�3��_�Yj��V��jɰR1Jn��j����'`�)6P���E
_�q���L�ίR�Z��P'%���$�%���]�'�4H���]���~�OP���É	S=��!�>�=��!��W#(��N�$�׆\����xw����a���h��[�&���aǇQ�&~Z�zH���� >�!���gK#�p�MW#06�y��7��k��=W��}���3�ʮw%ޮ��.���?lW�o�nY�.>���KK��<���t}�������9}�
�kL���0;�W�Gaq�apu[�3=��o�Tٴ{���4�?
TN�-&{�Z�����6���z�%�4�����Ii�3I]��y臞�D�?��tU�V��4�}2��O]��5��l�[85ј�\ŧz �Ib������L%�;�D�j T������X�k�?�p%8S�a�ڢb8��M�&w����?r�O���b��9h����I^�j����ں�t��q���{[b�
%�)���2��#��/@,R ��K��ۋ��˫	�7㽕�#*����!h�.�L;�Ĵ^L�xbvo�,HypE�lK����X��C��5]ݶ����X�r� � �¨���[�'Ө�fO�� b)�!H�g�&��	���ښ�5˂ض��:ls�Ǧ�g$!{\��<�%7����Mا��e����7T<�g@LX�S��i5��?�P�Q��{��������aKM��k �1��gRtNoY�&�I����2��Ij���3�L�U����[k ���`N/��.�>�U���Mbg��5��̦��S3�EM��ؽ�p�N���<5-����Ġϊ ��[�ˢ�]d����D�8 P�|�$Twi,T�X�d��q�E 1]�R~Y��y�4)e"����� ������������t���Hٽ &��o�W����5�>;�bҡ�aT;�1��a�
�����Y vV?LC�\�
5D��(���'�lb�X�J�h2��$����#h���'T�J��$�5�n��Rh�b 6��)�����������f�g	 ���@�D�,U6�bY�ր���(�a���'澝��/����ނ`D�b&s7��
R�ë+K�k�a3��'��}܇��NK����=s�@,-I'�󥔅~�7�}�f�PK�7�~J�?#dco�'�akwĄ�d�3�Е�����KA��ݙe��ݹ^��R%w�3���b��mU"	)w`���оÀb�K칸Ꜳcu^�1�~3X �R��*�|����5*U��"{��L��I���U��^q�+��G)�$��ۗ(�V�F֒V�JՁ�Z�~}�G�d��KmF��u�4�Jr��%���l��q���>
�������f�.�����{g��Xt}L�T���Q���
�n}jN8� �$L��ߧ��p�=v" ���z~�MV�?� Axv
w}�ջ&��0�7��ň_xLdp�UӃ��O���a��^�L���BoZ��	q~��<K���,vs�J|��k�5��zY���Qx<&1��b�&r��a*#K�!I>�~8�^ F��a��,LM!����UW�bfU�֩���p\�a[���#br,&>�F��DL�SN��$�+b�3��̧}�՚[9ẅ��< �b[����ŉW�Cc*���~��ZeƐ�b��o?��?m������q�tŚh�w;GC�� [x����lc������v�d�(��?�P���P#�C6B��y; Īa��>D�<��X�-��Ng
b�]�0K�i��a��*nyX5�逘2�}�w%������~ѓBS&�$�ɌM�����D1X� �:�=�W�t|���
)A���r�L�3��ݽ݃�ٞ�P�V�Z�����&��^񥲋�U"A�~��^�@E�g!���E)�bkii��J�sO���4
*T�  F
�z@$a���7���G��I� Į���<:�,5�j���|=ѝb��0��M�k�|a�MBu�1���P�H1BE���J��V9�Q �Z�3�`����K�x0���Z�b�T�q�<C�{2�F��X/�+@L]�+�ؔ�Y����2Gkc\��a��?��.� ~�c� �D���yF��0/�`.[�X^����w#>� �Z�)���b��LU@��*�d��.�Q���+�D(~!l9);>����D &4�o������gP5͹;ڌ���>>���l밐�8�9Q]�?���W5�h���g<� `�M��Wv�E�^Y�2����"��;3ĝQȖ-�;��!B6���{�{��=���^�KMR�'�w4��s/��BQ|���j �&AI;���cm8�#��bLU�V��7�,�h������x9b��=��4��I��X�K��2" V��N����՗��Ƅ�2M;A���q4��!������;{�F�Z����P���TkA��k��y�����K�0������:ҟ9>�2�Y�5u�~-�*�'���X�?ه����>д�bX�J��;�9z[��4B�RWiăO�Fj>6־��g���{�Z*��mK,�E���K�
����O�mo�Ͱ���,�G��b��Wݮ�$��[ٞJ���.�'��a�������w��������� V�fL�t_l#E鼍��\��1��E�d��U9�GoΝ�wG� ��).d�9f�%P�}��1���N��{��ts9���~����{|i~�As;�d��H�[3�����R���k���-2����$$X�U��A��V[e��y����9E f�"V�^�[kW�TS|{��}��	b;Ů�֋	oH��N�T�Bu��j��Ҝ����{Kx]�/hb��b/�l7s��3F�Vmi�_�V��^��f�.{����N���ƒ1�q�"���n�N4[������D>����"�1m���c�_���vI!v!E7s56.'i �φ�pS����r�i^n=>2��E	��3@Lo���l��+��-uF��?Y��n8�!��������$�U�= ������N�`l�/�#�8ځ�52M ����e<�A��`iĝ���.���8*�m؍��ё��/�!�l���6�����qWp���d��;��
]�^���ߠ�1Çy��e�-��y�*P��� �Uu�1j���|�t�J���y&	b�Q��R�[��;~������c���t5��z�w#�א�`�wb��o����[�YR����Eb�O%8���x�7	��/���/�X���V{���(*ӹGO�{���A�����Y�~����7>4��b+%�����Y}��N7^ū:��������b��Ǵ�o�}��.�'���j���>�Ե������0���(n+�ͻ�X�~Mĺ}<��}!�)O��a��C�M��|�y>i%���<y |c�c�蠼=�����u��Ģ��Id$�K�����l�����a~�N���]��|���H!�8ku�Ƞ��֬�K��Cl��0i
0�]#�.F`���<�/���1�K��<��iI�<�e��i�Ћ�"������'���\gHh�MW��Je�V���
Px��_�׷{x�Ubm)�-eX�EJ]=o9xV��5� b�ȡ)��;RZ���o�xg6�����Ԇ�/SJt�)kH��Z��Z���?��o�֊^�R�n�z�3�B�rè��^P���3�#\�u����W��+�W��k�/#���@l]ѻϙ�����G�9GXN �L�"m�5S��/;S=Y٩/ӿ)]��y?�\sn3�h	sbj���"X�Ի:�_4����19�0�ҥ�W�iK��x�ۥ*���~�鳟��&R��β�H+1��������o���W�/�s��!�jS�q�1�\�%�1��/����r�w�K\dث���Y�
��qₘ�o�^���1���� �c����U����geR1ޗ_�W������R	1!�7����[��a�)�<z� W��j����A���=����<���*׏Ϝ<�h��n���䒿���]"C9���w�7� ��,�A�_��(�K$+��-KU��|���g;1�x�k�:x�LKb	?7�����{�=~P���҅?߳Ү���|C��`*@,XY.hVqY���v;�v��;�<Y�y��7����0�ѧ��5֑���$�B*�˽��a�N��R/İok�>O���9�|$�/u���b�Ju�k��{�b������]jQ��	��5U^��W��jZK9ļ�3��0���~��g����]�g���ML�
�E��(6À����i��۬��$��}ɏ�F��X^k��YoqC��$L�⾙��6->+�XÁS��_��_�[�t4hqE�m$gŦF|�$�
��l��9I�t�725o��t�1��z����(uαC?�ν��Ɉ�4�}�b���W�&ӣ3�U��
Su��j�c�x�*s�yr`����ld�?���1�7�BNU�t��e'.S*����ߺ[��*��R��%�����9�Pb�EH=����PaLӇ�Ɯ��� �Әa)�fzR熤w�(@Nϕ@�d(~��
��xt��؇}���b�
�F�"g�E�z�PNqP�������`�&G�C�tR~���}���<1�UEՁζ�L����XM�<��������G���t�70}떃�U�_1f�,�T	�z�͖�$�Umt���������ʢ�5���?��KB��`��Τ�n����D�<���Hf�Ti�Ų�v ���g!?��!ĄX��M��n�����-]��$�M��������!xs�|���1��A�*���oS8a��U}qs�כ!] �X�V���DOr.K��F�fJț���I�/���B	�A��3cT��56"[��O�����u�[�t7��>��c!�*Gj'�Ĕ7�=t�<�g�X$��Z׺C���ڊ�%����a�p�Byb��75Lr�r�2��֑k��A1� �!J�\Kz�S񇇲�t�8����0�	���^9���&�
8�i�uq^�IZ���]�o�1e�j��?/f����?o�.3�(@�L�X�E�ϰ#?c-���t����<m�oW�L�q�x�8���9��no>�Jk���u������-�{�
}����|�6�G�$� 1	;�n�,m��!D��)^��Ϸ.��m>��H���`���U���I�h�;(�<h�>Hr�����@lB���Q�>yS�z�p�����>ĸ�ݏ8(~fRBcΐф�# �i�M0:^?��V�3o����o҃���f������RUvlE-L�[]��q��~�,��b�ܗ�$~'��m*��?O7��	1��|~��t��]����р+�����J�b��F#3��R�~5@�g�Z��D����(�Ȅ��ϩ Č�g��hF���)_2�qn�9�i���EoKzq���5��>�^�q87m-���i�n���'�8�3�	���N�+��*
-\O����Ht�i��N��ُ9��>�sjQ5z2+"G�楲�n���lq�A�fb���J��!��P�.^I��x�P�C3���bg"��n���j��,��Ͽ�`<.�X3.�YQ/����]e����?j�� ��l�˔=MI%��B�k�u�����3�a�4~�r���泼v��W,�ם^[�J�e�5׏�)�XȤ�c�0�������I�A��a�q�g>�X�],��ˉ�Ƈ����r2�,uD�����9��*�t�02��72>5�� ��nxF���BC�4�2;�F�)�,�f&�:�9Uڂ��p�5$�� Ɯ�$���8Ŷ����;_�N'�F����[�ց4���G���#)v�5,幢Jm_~�Ԣ�bXS�O=��b��c~��.w@���ʐ�G��~/�E�x��;� �vd�R�	���n2�"2=ɃX���Μ����t^D�r��)�H\F����K,��V��݉N1������+�Cߘ�'��e��)(S˶�R-��ҳ�B�;�V�{�n�W/���u��T!���y+)���+g�ۃvӪBb�^=�5Xڔޥ�zRma�	�@l�R (pқOq���dGS8��%xB��.�9aD�_Mp�!&���)mD@1���Wa���fJ�X�9�.Z�\Ǹ_m�|3r��a����c��t������Uk>#�H6�s9��D_;Bl��v��z�r9?��X��)��1Ćf�M�Z�ř�������A�*9;-#_�����x:���b������1ʥ��*]����GEM!��<�@�2���Y�X�J�y߄X˟
� ���l?�����C�FМk�2��7��Y��_�Ƈ�0ͼ�b��x��'DN�k�l�i�W!&Y�˱M�g�*�YsF-:֠b�K?}<��f�����y�y?�PK���
gLN]HɃ��ܷ�6+��mP��@&q]�Dbs�H`A̦^�m2U�n��tQ��`�K����s	/94����m��O���b	�=Kw�\o&U�_�\����dn5�Di�U��<��}�j��1��Jָ�0��lu����?�1��t����ݓ��/-+�X4{��3i��W']��	�&dB�읷E�IYVM
j�hS�=2Lbf���p�GW������&�1�t1��1e'�-?154�x�q!v�^0�2���1����K�.��1�B���R��'��>�%��_&!F���ъL���-롬�L�;"�~����g��,��9�R_e� Ơ��QC[J�+��'s��^���4�UT%��ya��Ї.`��������w<{i�Λ�w+Y�@��7	ko�'M���K�������!��5T@p2���HHcĝ���:����C�K�.v���>I /�<�!in5@. �I�E�έ��p�*7�S��o����&3���I����X�T1�V	juil+��>��W�v!��E1j��Ӑ���%;�
1��g?gK	ZK��YO��A��}�Ԛō�A�\��w��ʹ�чYõ!�65��v���qA̭�������jg#��)O�Ģ�U�SJ'���j^`�ɝ]۪���zG��0���&�8rc]��bq�^���4�{�ER�0�1�c���8e
euP��X�1���ܨc%[�(VI�D �~�E�Al�������yi#Jͮ�o�#���ɔz�R�a��͸�����d��0T�E�`�1F"�u�!�b¤t%G�*�)��I�7�]L���}x��B������+K>)�{�z�H�5���W�(!��d��ߑ�P/��ؿ�~o�� b�q4�2߯��l��,�s{�U��a��'
ėm�z�ǝo
�7��AL 7l�Y�GΩڣӜ�j�A�1��3ߠ�J��j�X�C	D56	�C��" c�O^�:�W�;D�J��C,1#��E!{x���5�kga^�&=Ć�=���[�5��)�᭚@�G���S>�S�[ED���1�q��Os��"�Xyvߍ��$�b�'x�w�E�)!��T�gv�[!G9��W�z2�|�:�Ȓ֝��^x��������lF�=�<�!&��a*���ʘrs��~K�x9�D�6�.	LqL1�Y׿�"3�
����XtY�]B�T������sV���a0͉�[e��ˆB��ms��u��Pc��JOd��c��O[<�XV��$뮲)ފte����p���F��ݲC����[X3���e�q�i}���a��E1��x;�{�b�O��	-�d��W fm��>N�k&����DzBLk�xU�ǔM+��(77��%�^;��&���Q	�ԡ�:�g���ؿ���-h���UTl��a�AR:$	�n	�PBRBBAJJ��FZ	)��FؠHwww����ì��0������7*b���E�	��<�}���ZQ ���S�U�9p�&��վ_���-�S 6
��<k=N�g@�Wcx	b���n�U˓g
%w=|^��ݲ1b��]��J=�Y[�|�l*'�Mwn��V�u�ͤ�?��-���V@�q��N��V:��m���� V7Hhq{w��a�����JFk����-@yP�d�b�	E�֋1������z�B'ܿ�Ph\?c�-y"B<���P芐�߼)���O��D� &[��Zh���;�H5u�e{b1��U�x(^�vXU
l��*�|�y�W>U&IP
������E��=+#UJ8/��w�
Jo��b�!���_�mB�6҇$�nY����dq]����{��.�}K�6�����%+�ϟ�.$��p�1A+���AH	�D*��2^oc�*SyA>ڕ8'�켔}|�b�k����89���a�J;����،�C��v�ť����oA,����ө1���J�T����(�:��9�2]Y}��:ͅDPbM�ӱ��^��݂��������UŲ�(l\Mb�2޿k3'h�b^��K�#��Y��?�Q����b֧gp������;H�pe�R��2�+�:c�3�����ÃD��A���cީ�[�U�1*����AL��٨��d#?3�k(T��o��9�e��±m	IY� ���kkH�& ֪+Vř�}��c|w��ށJ	'��Q'�qRE�RQ������i���X��=���>#�G���D�͟��ؐ�,~.��tNeIvC�oD�3�}��\����Ը<凭��^���e&c�"���6H�OTfΜ�fQ^���l����DY7��d�N��Qcx#ě�aN�����钱�^�N�/��_&a�lE؄�hQ6r5�(v��dV^	���Df��a�3<c�� �=���ɇ��Ȥ
�
�g�mX v":��t�zW"��?���� �N����eh�G~ӣ)��5����n�o�|*��o��!|`u��SĜ>0��>�sg�j]�:8��c�P��WQ�R�^�I�נ5&_A�N�כ�^�iZq�d�9�-�����9v,�����l��7�X�x��V}�N,�`���-��u��UD�4���ijOQ5m�mg:/@C�I�@� �n��{�S�KRa�FϠȘ[ Fj~��d�C~��2:�kw�i{��y#`��e�����M_2�7��o��em�`��a�D�6ً�\�1� �7�''�_ve����@L���-��N0��X̒6�bFYF�5�w�]G�a���c�1�4K�DdTIK��|^� 7��hm�D�Z�!;�tUՄ���d2L$�!���4�࿰�_V�%��I�f����(a��J�Sp���z�fW�Y�2)���ɰJ@Al�ee疾;�a��AW<�N�مK�OV�}��}�&��x��X�O�M���U�^��&l��;�����%A�t.�D2H�s�e�07×7gm� ��\����)$pW�'j��y�ߌ�Y\���~)#����L��~�)]�&bx*�Oz�V����Ej�Ⱦ�#��-���<;��TT�G��c���L�o���4��ǹ��~Rtݚ!���'�J�M��>
���s!Q��3#/��)n&{4�R���3��"�&m$˘,��J�?ƹ��b^��'����q��?iy��b#�7폱0C!|yw�1������{��5�c:+�w����p80S�c���W�Uf,� �������b�v���{K�����;fc�32�Te�JS�@��]ď�M�ay*3}]ּ���/a���������~8��4��3��R_cL[��#��L��������ҝ�9�<?H���&P�~��g�h�D���6��
�ᠴ�t�m]1�E��>/߽�a�e�W�v�~bN?��Y���a
z=�<]�G�G ��"�u~��ӗ���k�DA^��b�.��d[nx)�eL4�2����֓��z�8�H�`��r�1��h���i	�n�ݓUS*7@L���G����d����w�!�����e��>QCԆt��TŇ
d���f�/��|���i�a��b�S�?������&�x��`3����k���fm��!�)Gs+83�+�?��x��-�wR{bl�ќ}JU� �l5�*��oZ #�^g�t"��7s�_ꡢpM_%g������A� ��%c�0��sUG�|���0-�iJ����W��D;5#�x��i�&����J�b��*?f���3��.^Q�95j! �M��t�|q>�4et�E�X���:�a�e9O�>+E��;u~*�30�{�u�2�˝Q�@�K�������d�m f�Ca��՞�ҭ�,Ñ�����X����1Ca8�������NA��*:��<�����:^�_�Ȭ/)��T�l���P^���ޜ1I���
N8N*Bd_��m�Y���ū:.tͼ�ri�[X�e:��] l�]���?ߐsyk��(A�C��મw+Ct�d�ã^A�d7���&��vF�D+���o+�S[?@�bR�~e�,��E;Q���2�Ps� ��M�j�d����0�|�������L�����Ȟ]���9�0��J�a��~�l4`����X��P��FP.&���$���7?e�Al,fI����]>A�u�1�7W	b�j�A&���i���a���<� F�]Z!��"��%�}Z�� �<�Ĕ1��gQ;u���xygj(ҭMĮq?�����Z��Q"H��>_��H����w��Bz�� 6�:�5?��=� �I��/�X"��^2���3	Tvw������Н��;d�@l��YT�]־�mJ�\[�S����	��{ň^�����Xr���(;��HKO_H�����k �g<g��͢Q��n����!����5��Ni�����>D1hWN�X�d��d��Vo�gT�?��]��d^W��w�>/?���+�H@!=P�ׯ����\��%�{�$����5=#�"����;Qb8���h�߮�P�n�A�r@�3X�EcZ/N����Ĩ�a1H�=韏��_�������,BRn�Y$:��F�sP����l��}�"��b��jҕ>K]X"��n�����BM\�-`��Wim����9�竌���'H�"��� �m�͐������e}T_Ґb��	��O�\� ���5�액 O9��T�t�|6Yr(��|����0��ܺ�e9���x�8�s�x�V�02u����aSД&T���� bO��--VO�GY�=+&�{�f�ĸ���:�n�0RY0s�A��A,�{r&��YEZ�kҥ�6��^%�vR�����g'��Q�B5�%��F�/��s�zU���-��rS�n��1I��Kkgk�FJ�Xys�k�1r��K�L�V�S��lv}E���o;�Y}�4�D�ӷ���s���Gb'�U�ԟ�e7�芖���D 1��I��]�=Y3SJ4�#>K_St�{6�
��@
�Ѩ�cf��\骬�p�="�\��B�H�/�o�u!|��5,�/Z��R�X�Y�C�O��q_cSYu�o�p]a�2�cG�����>�RR�������_��7��N�g�\җP��y����-���wN��b�	ߔ����:V�E����k�����?��5�3�n�c ��[����d�Meb6�-'��.��
��kM�ܠ�b���pc�/v�T���u���U��y�o�/���J�%�@,x1�E#T`�'�NRC��٣�byLC:�݃�q��::Z�ƾ��� &����ȘlL�j���?I��b�����G�C�nz��:My!�U-�����ω_�w:�rÌ���H��%^X���䧒�vٖܝp��3��
*j�U�WᬜZ�G�^�� �4�U�_��[��J_Ò�q[J��������^� �k8Io$m��R�%Y�<SNA��D���ND2���
�h�/Ds K4tv�F�)?��9e]�r�¦��Y�z�y�|�J<�P@�-�v���/wn��eY��l<Knl_�.	�f����w�,�����1��C@,#Յ�}ŕ3�V
�
��0�5�j��r��,�q������N�E ��z�v=#�0���g�~@�i&���R�Ao�����h����	O�+�Γ.�p��%gk�X����8��,�������.��� [�Ԏ��1����g����P��
� 2G�o�r��7���jA�z�fpƒՀ�APe,�^�`K�0��7�w"��CS�ݮӣ�1�E�|�)�[=��,�'�Ut�b ���5�yJ<��Pe�%<X2��v����	m�M�:lКȺǧ�bK1nu�~�J�K�u��K���A�D&�I���b�t��kbZQ�[ �=�em�lRds-��ٸ����hi�e���	�J�@B��.� �8��`6	��-L�Ñ��kJ�s����a)G����B̺�"�]��,���.waos��a�+7"uW˕�}T=�Ai�r�wd`��U�שMb�Ĩ7zzZ=�ϘMTSy8�i�}Ae��x�9ߜ:Qe�-̙eM���"c0:=�1����/ls���0ĬV���V���*�hKɒy;��(YQҍ�m��[6��J����������s��s��OG�c[R@�'���b�p=�`����y32���'�B?͵��)�W�~1ӷ��)]7������bb�<�*/�X��s���p��ث�X�פ���om���'qC̙�� &�@.�߭�H�����"ҕ�d��d����7�)+��U0<�v�bA��<��|�Y�h�u^4O��;� �iJ[�D�v�rl3����G�KG1Sy��CQ����ʩ�Q&�(��w���b��owS>������.b�ل!.K�K��ӝ������®�B�Qȼn�K�e�`�$l�{pa&W�U�̼Ʃ]vR;�'����G��}��� V{�Ut}�Tm��x���@�3�y�/��ߖ���)��O���yL1��uE��څ�\aWu�k	�
s+*>��)%��}�5�@�ޙgm���%��m�����<�b�{7糨v8>�(B���[�A�8u��h���B*I�\N�!�V(녭�����=�k%��9�<�B����ks����r���1~bB�@�nn�Md��.�o�CG�n��f��s�[j��i*��Q:!m"�h��F�8%$�)��n%n-ay�y��q��(M#��Q/�CLE,u@�7�˦D�H{$ӹ:-sS���Q;
��"�a�-���.� f�����ZW��I�U�,� <؅�^aWu�A_8zI|��� ��N[n)1��b�,G�zy�*�ǁL�y� 6&Ӝ�_�&:�4�b����jT+���<~�ξ�E*���-��p8ޑ�VT����p7���x����Ő9X��G�O[@�< �<6N��`8e���05�J�%y�a��.�H�/v�����\�!�m����+�:�w+�3?��l�d��H���b1U~�"�*&�*���U:4��./Iy�b���Q���b�z�<b/����6	[��o2���tn���ߘ�6%��b����&��7BQ:A,G-��:v�ɹ�z����T�?L�wK{���eȸ�)���t{N$Ć��XD��g�X�~U>�䛂X�ާ�[�x��|������˃����s�h���eW袀a�[B�KJ^��i$��A�����x������>k�Z��8�|����<����&�X��S����Sͦ�7�?��Ѯ�1��x���~���J�`&F��|��ish�;W;L�	b�U�	U"×�GS��
��ŗ� ��D��DZP	-_ur>#,�Q�Q�Ć�٬�ܱQ���ء?�^����Q'��"��J(���t���?C@�M���w֦�?W�Z��ʯ^���.VI#i�d�=փ�^�)o-!�1x"ҁ��0xVC�f;,�"���1��\��7�m<�9�Q_ʠ�ؚ׳a�ؤ��A�蠲�t��6�o�ɂ�����>E&2Z��<�l�-c"Dl�d
������f�#}j;b-�gxkw���!�\c�2���Ҏ�c��^+C�P�x�j	m�Tە���Lzd���s����`"b��ϋ8�E����
7ܒw��f���_uE��|JDh�k�'�צ��#�)@��*獕�?^DZ�����0$���˴ߣ;��y�u�ocY� 1�9�x�g˸�[}C����ҙ� 6J���x����,�TV|cW����תz|�q\i#cúj�&��@�:��ı��rhp��Z�v�k��m���:I�Q߀�7�mt��)�1�/�`ؿ���v� >�/x+60����� ���q�M�7멍d�W
���@�e�V�K���GU�{,��'�DJ
�`��n!cʦ��N�/�8�kE���ԉ +��U��s6K��M���݂l�%�)䵬y��29�(�����3���jN�g��%���\Y@������!�����+���G�JG���wb�V:���>�<@�1v\]w�L�L]�V������k�_�_����	�!�-'��o�>�*� G���8��S9߃~뉴j�8,�}���ϱ�{MK����7F��U'�.�W�3�]�?��=�|}��MJ�z|'e#�h����.f�p
�d��W��h)��܏��ق�ke �Kg�x�����y��������t&F�%��Q�C�<G鸿����¼go�t�4^��b���1\��SH�j�S����3��+� F���+�=͒��Ub��d�ŷ_��_Y {���B�,_4q�\���Ȩ!��W{�htx�2���f�K�"	�b���g����|ؕ8'^�ܣ
�6IG���u�GX��8�)x�@L�o���7�ř��>��hT��D�J����h�����G\9|���q����q���*�06��?�A�g����](w ��Vl̛I�bL��aG���y�1Ep|m�{+F��B@��O��gڢ9zlS���l�fR��X�Q����b
qR��AFP��Cʩ1A��1�[RQ�*xC��z�e]�q���I����b)�F��n�`��'V*��q�@�ĕ�y�)��j�#!���g��#s�WD_�2/����� GU>߆������>�F1��"���+[ v�9��jDx>b�T���B@ ����\9�9J���R�-h����Ũ*�K�y�3��M[6����Fi�:�k:QQ�h�q�d"�M�d��Ą�.���[zCN��A,�D�ҙW"o�ٻ�VL�u]S! ��9��H���U��*��b��ߘ�����l�00dʏ1�iJڎi��Ω��bPZ��cF��D�R�41��]@,	������P-AHy0n�JF��o��Ϧ�Ҝ�Z����G��8�&���";�}/��!�3�%�k�G���n�~�N/��,i���*�ia�b��8��(}jO�L��:��@,�!E�w3r�mXcf�!hGl�v����񸀈E9�>�vXφ��=Q�Ĭ*'�6j�c�ج���a��#�@�__H���ϥ��w'y�
bf�%��7��vK����/g0���@��"����I�k�,`~&�M�F��t�U3؅����W͹�"0 Ɗ1�Z&�
%ωP�ߜ��m�1�ب�=�����)����i�n��T�����m��J�J�b}���w�bs5i�Ee��6# &�ƶ��U�~e����*���tĔ�s�/
W��%R~�eM��[��̲���zl�~�5�+p�#5K9U�`�4X'1c5���GLS"CUT�DC�%�1V< tN�1\�鉑�P	bO�������]�g}c�|] bV�c�7���o��E�4�b�@�L!��嚜�M��{��Nzz>�d�@�\��tT�M�Z#?+b��l���%��ǅ99Ɨ���d��/���J����9k��MV�hX�0�2,ǗHl��Z�ĥb�l�bj�@�
���1�@�������s[�I��|	Ra��?��i$�m1
�S~�t'��D���ʲS{	��|5�а��cG����]�����u�aX���{���	��!� �){��z��m%��W�bV�.��g�Ϧ�\������β�p��9/%=�B��t\�#)ɉ	�� ���"���B|��ł�_�)W�Y��Mw��"e?P,nj�N��F1	��������4�7��?��AL2]�,^�Y*��Y:����@l��>����
��z56q�&��	Ķ��t�]�HNyu��(����-A���n��3��ae�Y�G:�h�� �}e��0���\0�� ���A!�u�`Cj���iD����l�bAlx��Z�Ͷ�����eւ.�;�A_c"WmX�B�Á�տ���1�Ov�u�b�r��0+xm-P:C�b�$��q���и�3��@b�V��Q����%�ޮ��y��h ��eg�j�<�.�h`�\@�Z��v>��v|F��`}��mq{��F b� &HJ:_����G~�,U�b�F6~�����ʁM��C��I�0���n:H��[%�1��k�:_��]��)�\��p �X�����dM�h��iz���b:�٤x,����$R�
D��2����ms��{\M���S�@�5����:K����'Z*� vaAX�gd"�c�.?-�z(����� ȩ�K��%:�x[�� ��u��hʒ��'��S�h�T{'�fUw��.XY�ܗb�zFb�]x<|0��
���!��� 6L��v%�#:GԭC������m�n�վ�V>��MN3�b�����w��Q��]q��-L�M@Lٱ�H�3w�ų�hW#�ćK
 v����܀��{KXu���Ó6�$3�P��
	�]��I-Y���yb�	�_3Ռ�&�-���e`��К����*���x㮃��zk�V:��^m�f���$�:iYYb��tU�G�]f�1h���N�I &/eP�|ڐf�A�*�w��5��d�Ld�:!7�����mq��v f���G���V�敋2~j���9�	}K�L(�Њ�6-aaT������C*k�ޭ"O�cG��ـ��� /F"\Z����X�E��~^І�&�ƙ�6�T�bE�f�́���3���3�c�� ��,�G��,ͮܮ����+������TK�K�Q�����G<2��;�f#�����$���.�=�� &�$8��\~�Xӫq}+u�b:�s�7��	q�3��U��x@lM�jVd�2���H�^��m�=���������J�A}b}hPߐ�R�a'��!Ƀ���wK�!]Z��!y�����y[��`��!�f8�repJ��5�Gο0ſ���9�l�V�2��z�&�`(&��Q�����Fa/ū{��CfL�0�E�y�7X ��Dw�
��xci��T�(j�=xC��q1����u��F/I��b�x�f&�%��r�r���%J��˛-�؉O�4�=�/-�	���h��?���Y2���8jd��jq�/�A3�L.5�zW04mdU�.��=k�b��Fތ
u׳�	���!�
$2���˅����b� /M>�$Y~�-��}o��dG2	6E�C�����'��;�ֺLZ��<��?��^C�gt1,1�3���	s����
O�vg3@�QH��O�a�G�$�)n��?��A̖]�B�����c� >�1Ĕ߱��0V�8���	xq�b�g'�؃t5�gU>��ap
�Wi;�ۚ�1�k��{����9�S>}�Og�s����c�`��U�cؤ�j�ƒ�U9����*DΈ�i(0�9�n;@��,[J��Xh�V۹��4�6��I�rg����qOjjH\�X�7l��i��������� f��B��3��R��>ŉ��<bWX�.��hz(�}i�T�����ا�ů�]Vb#<A{��^u0�|����5�"��ak)9�J_��l�X��:�E<����M���R �p�ܓyo�9V��]�[b��y8��8a�f_�|1%��wA,pT�M��4+?oh��w��<�
��y���%h�a*�0�&՟oz�bO��hٴP1����f�){5������`�7�Ϫ�hP+��|8�߭��!9\T�[<�K>5�M��uOK1���R��^��L���A��bl|n�՚����G�5]"�b &<sӻ\'���Zť,=֙$bUE��\	;fÇ�$L��jt� ֠�p�{�$���S����ӗ�6�H	(Z#�c:��D���!�ػ�YcO�̦��������� �Y�|��w_H����2x���M�1���Ebp�|������������,�Qq���Y8���<�H�ܟL����ԛw.���Xn�]6M��p������Grr�B���Lo���@L��A�^���c9i�/�xnS@�SWuV��8��	�tN����s��MT�MEI�3W�=�>qb����<,qz;
���P�B��A,`[��1���w�95�ҋ��2(+΃M��Kz�t^����X���܄���5Cbq8�ю���2��	&�BM��cʘ[�oxO�Als��dݿJż3'�`TR��U<�������a�T1�;kf�`�?%��鳷o�bu�����e$�`�*$J�Q�7S@�~A����R2�u�B6�NP��2.����<"�@Lj����(QqNށr�O0�]#bS�¦«q�3�8��B̕� &^���&,�v��ؼn�{�] b/R�	#̮�/mLdM+:`�L;#$�S�'nB���r�D���o���U��1W{�� �8~�Ѳ�i�%Z�D�ǪP��(��W�tG��?�c�Y�t�z9;����D��[�崖��GN�j�*r�r����Q��κ��F�U�z���I��o�E�[�����殊������ϸ�ͨT��٢ۍ*�@�fe�ߺ����xB*m�p��~�x��Ў?�!doۻ�%�RNW�w��L9���vw�GI�B�0x �f≅�B��m��r�l֦�%,�a�8�X�g5�h�t�&ixB
�As�������G\����a�.����CX�ק����9���A�"4~^+��
A�M��*E��^�)��Z�&q�k/ܳs̓'�$bph��ti�ܸ�SX�slR� ��f�k�vh��O�cv#�bD���'\j�O���`�Ve��|Al�u5,���͒�������
���ϑ����2@�ĸ������͞���۹�}����Ĥ��Z�/<-�'��E(�>�ՀX?Y�̖3�l�e[2��}����q�Ρh���uT肀qBRD���Ci����N�IiD�>Z�C�;E��ݻ���Ό3w��9π�����G�L�m���� {'&�_M�"�N ��îڎY@
���W���=)��GK�a��b�VS��Ibk���]�6�[�/�O]��^�;f[�jQ��$�d���yc_M�#�6�}�J-G�������x�[�3X�,q�� VdZHl�u}�� �\���;obA�x�]�c��s�(?�Z�gU@̺'ҍ|]�t�xz�+�px����\�A�q|��I����\ F��LN�#��U�~�YD)
�
bc��r�O$yϠm�B�Ɣ� fy�|Y�Ӟ�}vރL�!�<Ӻ�\l�����HTL�
1�N���E>Y)�Ni�"��7��ȓ V��X�`;#�%"��R�5���S�;쨭�
r�(x�	�˦�@eY�S3?��أ���o*�8�1�QҶԻO��jaBs'�h���~e�n�ԥc6y��x��]���&�)�{m�d5�I�AJ�T����@,���Ed~$2�a�Z��^{�Z1)q�qۼ`��0#�o�l��<Li���7�L�Ċ�&��g1��u���S�,W,�h	=>�m	�D�=��#�{�}�I�C�c�\�_tAԸ�H4��TI�G
�T-` ���Y�8�CO�ds���Ӵ[R;XI,}#ɺf�-"��uL��
bփ	�<G��8-w蛊U �8�ƛF ��<����B�z,�	Ql�{���hv'��ڭ���}q?J�,*N����'�;��L�z��)���l�&��h�.�*�ĒH���եlyaW+�T�ё@���HT�v"�(-�KBn(�(�t��ge�4A��OHDp��@,��]�(�z4�G{PXU(,�GC&�%�8�(�IO��!���y���v�c��yv;�������A�ꠎ2�j��_?�⧎&��j+�}�4��Z��p�P߈E��r��1�j�gV�wdϢl��"����m���v��� S��B��*tKN;�|�d�]�Њn?Wuݯl���wX�؋���9���c�����Ħ��: v�U�L�
�r�epI��$��:�i�'��,(i)����w�ZD�ʔ�LS�c�vEX>�
�N=����1`PvHPia�/��?��{��~
�<��U�pw�aUTJ��b��=B��ZM%
�O:��GMA��K'J���IQ���U�����m�d��޻Ϻ��ʵ٤�V��1A�P/��jT�xD��5a�~2�%��q�k8�Tq y|��	b�1xdF5O�\�ҭ�5-�~��X�Իԓr��3y�����2UɈ &�(��:����W(�U���yb�1&�x~��сqJ(5�Z:� F�"��K��,4�~ڧ�jew�_�I���,h/9𕕎P�<�����e���^IV�ߑ���߁���1�~R���;#Ud����y�[�^ac6�;�U����xU(�Ĳ�[�.D�	���g4���A�A,I/�l(�\�]��v�ޚ� &�ڭ��\�%V>��U^�4Cp;�m@L^F(U2����]1IAb�J���Z�by���Ux��\㸼��b#�L���O!#��|x��X �1�.a��"�-d���I<'лbV<|6p�)���$�p�����@Le�m��p�i�B�Mz<�TU���MO��e�ƒ+��( '�н1��f�Zc�%l�|7�a��Bk�A��k�/�\W�^v]�����k6~+�6�T�7S�gN ��6���(��Z�rȘ���B^�Z�60isTk�D��ӺRс�i�ju���}Z����Ĭ *1�9ƻ��L\�ɝF��V"�H�$� �u�����	�wD��ї)��� F-��6�+��s�}��T��`Ė�����s5KΧ�Jq6X�N@�BA/ND]J�[��	+��4b�|]J=F|.��%!���Oqؚ@LLͷ�������v-�m���W��4Oă^��Y1��{~�
F�~��3j��x(���*"YS��1� !�t�&B(��W�4;���>������/,�P#���ŜSM�X�]@Z~;)v�Q�94������vtI�KE�mγi�w�(���VA�LU���
����\��{��\C��b�x�]۲Q�"f��ꆐ\ �vft��
 1�l���e�� ���t�j��Q-4H0���S�]-���ZT�O�5�a1��X�f1��l*��!ˈ����y5wk���>�c9�1�6�j�V���\,җcihI^!l܃݌� v��~?���6����b�î��sRV����|���4Յb�^=f���N{�O��s<C�+ؑA,����xΙ���B��F�Q_$�n�=Y�0h���
�?0� �Gڳ�S'#�|/b.��Τ]@�4�N/R�ӝ�39]�N0Q�����>/�y�)̄MD���o���2M�=�Cc�|ú��q��b��|�x�%*[�>@���$;~�b��L9}*)|3��#Y1���,�A��U�S9�95�Lb0�¤���|�+��,$�I%�����b��!����.���O�W��@�LU�|����"�Ͽ\9 ���|�6r��b����J�6�t���ps��i@��Oƌpxz� v	u����׺-��B�������`�,���{˚+
7��e#8�J�È��y�꿸=���[s�r1��P�(A�:*�7��c� FZO��K�S����-�.��%y�|nZ��#��I��&�񜘟��_�h�؏�݇�d�Lg�i_���l��ZE����R��4m�q����?�V�FU��ϑѣ��X���%�7v�Q#y֠��E����-Z"�0�A�q{d(	tA�4��.1N��j?_��|,eu���4/_uQ�*M��<����^���W�	c�M�[�M�3���$U� ��N��.^-u$.d�J�����a��Rm�8#Ϊ�����֫K�ش�T���n"��Tā�6L �îsp��dP_�z@e�����	��%啱i�H���fxo���؜ނ�ѕW�a�
���a������ ��-���Y���G|2S�>�F^��$�g4Zn��Ü2�����TI;S�ZR�aJw������I�a%t�Sn0h9��W���}^w���)�.{4\�i�<Y�91�����[����m�N����bc�"��e�n�DZr,�R� v�=�IE#Ӟ��AN�~lb���z}�!*��E3f/D�4@,N nV棇��""�v���ba�Z�����~l%�~���	1	��Q�Я��=�|^�<�#g~ F��w�,�R�.Cb������bG6�E���[��y��@�"�~U�d�uF��Wc;�Qc{bzv��� ��ѫ*�Ǹ1[bK)��<�_#F�^���d ��؜qzvDW�ZA��7��!�tc`շ�86>�>����ڟ9]b�W|I�E����m0e1O%�A���������X#����'c�cB?���#wy�g���Xh�WX�W�H�����eȂ�i�mn��*S�,1q`�X0j$�9���\z��u�=@��m@�����*�B��ŕ�%��~w��J!c��%ӑM�\���[���h���.�U���t}\�kYn�9���W\�ǌ�D�qL�'F����v93���8O=��5����y��!�`��H����
��Yf���!D��^MCY%��ٝ�վ�B޽����6���u���\m� F{aje�塋Q�^X�O���b��A�YF�s^yiG�a����Y����٤~��b8?�]O�}: V����SV�l�[��]��M�Е0X�&�S�ʪ���1�1�*��.��>3�=8�7 �\L2�$��Q��ؕ$y�4��T)��i�ꡕ,@3R�����u@,��x�t=�c�����+���T f�Y������`��e�$��)lu�Ѹ-f�Gx����ut<A,�D��w8�8����ҷ'�k�r7���n�we������a@��)�=tK�{�َ���=U1�X���)k�_�[ly�<�6b1�p��G��p�2b�|*r��1|��,Ka)Q8��.��!X�bc_ن̣}��^e�Mt��l��b���#D�%y<O��/Ī��@l�a	b�و}J�F���A6<��]�����vd�3)��=��`�ߢ������\��P#�c���Xw[-5��@��(+"/ά��.����u��h��ɦy���N��Ĳ�c�.p蝋2e��=,�>��1��c�,XW�p�^X)��^�����n��3�$�����r�1l��CwJF���X��^��U
��I�$߯���)G����՛��=4���S?��q"<��@�fl8�Ɵ�(!��k�� z:��=�a��<F�v�Kc��3��c�f��<����9`��:E���q_^1>���Ew���9��U�U0���-�l��Ĥ|�pz^{'X�81��<����5��~�eGP�$:�}G��^������,p����_'f�o�$�S���;�G[ե�L?+0�8ѷ	�v|JјH1r��;�iȾ
�K�	��1�/gi=���ɲ���b���L[��+Ys 6�	9��$te9��{l���{���C7��g��33�-&'�adlsb*�C���C2>>ݼO��rA�@>j��¶`��{�c.5�� �8o���P���J =���R�B����eqς5:2��ԅ
uR��^�6'�/��w���Tr�)�6�Q&%j��^3����Ά��vu1���3G���`��Y����g�K�5�~�S[1lC3�B1
� `8�B��q���Z#��v��l��6�b��mwy����Ѥ����fxc�A�x��뇵�5�n%�aQEN�MAl~�m@�:�n%�7Țr�7s��ƒ��sY�����y��3iv��mT2�����8���>�Ϥ��E�/�`/��$ÿc���dҞQ��R�lY5����a��|LˑB�.8�s����u1<���a���!�H��L<�e�j@�md���Ƨ�a%{�l�������3��Vܦ�8N��ƫ}̽B�����sF>��Qk,/q2�Ij����o�]JpO5���zb�l���˵�Ή�?+���A�;F�!:�*��WgE>�fx�L ֛[Sh��J1�� Q��!'��)qST��xN^��� '5aX�cѤ4U��O*�S�\�,9�@���Õ7*�ͧ��jY[&P���o��mh���j�~Jij͑�FZ�{Ĭ�����/l`��ҷ1��^n�������}v4}j�%����4���3��2�}'	�/��]LF�0��. ���y���y�WP���dH{@ݮ�*���
b���^��	���qs��� �rk�&4w����I/����9!�>��-_0�{2�V��ઓ��'?V�ύ`����`A8���Rz"=ǣH�wF�;����}��^j%Y8.8m5/�E��3����z��Ɓ#n�;��d�O�h�[��W��g���d>w���q��3��.^�a����� �����������x<�N���4�fL0�1P^M�f��4��Z���Z���$�;�%�+��s��@s�}�%�������-$�;ɚŅ�$������ ���h���g<z�q�̌$�̬����W���^�eF����{d�d��^����9�������w��6iE���>�A"�.�p��"����A�c��1ov��ۣ|�r"y$�d�!�K�][�]�l������zml���������]��Tg{ҠEW��uP��Q3���J8Ref!o�:��Q��Ic���QR�k˗	F�>��:J5���`(򛶟O���7�Ygc:Aa��֘��f�
b"|8i
���?�'�;�$��x~�m�̹(��5Hq��a�b�ŁX�z���t��ʻ��NK�Yb�7������f�;�]&�V�Ո�L?�[��� �@tL��zBR�#_�An�hwC�w�-�HnX������0P���Ԫ��$��y��۟U5��5:�X���'�DA�����F���_X�����6��^�ן4�4g�d)Ac�ҟ���Ù�s��ۺ�S�q��`_u��ݚ�#Ԣ�Qŷ"�zI��A�
]3�lVH-:>Եu�bHT>fw�=ӷ�첡��c6���F����"���$^<{��yy����ĤYJ=T8��Uk����%G�A�I��<��0)~�9�Ք^�eÚ6��e��mz,�%�������~��WY��`�|8z��/_�����b�R|g��&����;�F%� ve]E�D�6�1��e�	;l7�ё�H��.�?{���	qS���D*�NE�X_�'�g�6���b�r/Y�>�{��߯��Ě[pM��n>���0o�z�f��삽��}�=���"Ի���Hy��Q�~��O�1+ 7���	��}�7 �����;�$5�w9���e���Ă�	���1iH!�pl,��c ���D�Zu���̨�WǷf���e���������D����#����o�]ӕ�qm4M5���	�3p._��X���?f�s3���č�?٭���L�� �>{x rN�dޘ��`�g	b7�g^/;yW��z:�N��PɃ�4V�=?���e��&>-2k@d�nn�.t@�/<��?~�
b�K��D����	i��=W٭�A윷h��SK�m�ug�����2��sk6E�Rhd�:[Km�c+B�w� �c�����5(�_Ɂ'l��sV�����8+wp9:V[�-�u������3=�AL�6���������3$#�͖�0��>�7�iZ�ؓ��u=Ժ]�C���PJ������Yl�d��4ǧ�"����߈�5�;�D;��)��� ��G<J���_Y��`y� ���g�-t᧺��ֳ���ط�����	�>�:�&������������nj��@m�0Fi��YctB�֬����LG�c�"�
�s�O�}e��ۖ�;�6蔥]Ë�4j�)�$�A=�xh�͒��qi@�y��w � �f(%�H|{��Q����rZb����OK�4'���Qt.�X�~��(4h\�w�Dg9���N��!�//��(ɣH�%���-�i�g*k���ٓ4�5� ��o}m����6�Tyң=ݏ��|@@q�?ykB��a��J�tkV�tHmq�ث`��>w��	��vF�~r�, �]#:��8��&��ai��b��v�>�2���=ƞ��)nA�����~�Ɉ��O%�O5�8���X#q�ݎ)X�>9�nl�	�S*�d�V|�W����IZ�T.m9"[�蓺#W�T��z�e�����b��*�z�Q��i'cMZ�}^�\��Hx&@J�0�b*h�DK�.d�E:r�.��m����(6]� &j�Ks�@�L�#�8�:j�|4��D3?*�s�3cܗ3}a��ĸ�ē<,sd�2g�?۽��u4�����jը{�J�*o��DA�����Aό�{=:���$��9Fc}�o��=�gMt�g��i$̉����taaqR�s!u�{!�������Pjrܩ��0�!mͼ{, Vs��;rt���x��OY�G�ʕ;���o{S1�Wl#�����ds�v���"���⪂�I=�\@m��E[��ԉ֝:w�؟��i?9�n��߸��H��k=��t�q�"�	�ܦ�Al���S���9;�|�@^y��n��?9v8kWF��.�"GW�,���K��1n	�����zL��4��5a1"�Ѳe�y�-;�7,�s�~���z"�|�5=��}��r �΄x�t=����K�ָ�Ŋ�{��s_�&<s�l ;���N��O�N�5q($I�)OO7ALn+
N8zyL��o��t�jk�^�w_Ni���4�8x���"�b#�]�tu���ς*��?�����bGc��3O�Ы��9��� �v���׆��?:�RWH����Mh6���V�Z��5�l����+�:��C&��o�
���&�s+op�8A�L����z�x��eĒ4�����g��aww���A�pη�¹t3^�-����h� ���5��,L�z��xS�WA,��wDp� �`�.�&��W�L_����1�ך���7���{�5��d��Ao}�JB��@c�M��$��Ď�����d}������ͭ�1D�'W�ԃ�M؍w���9�@�#����h���Lk����s�@l��&Y�z3��������W��X�%�;V�R�'����}��&�r ���Dm�*
�7Y��q�� �=Cܜ��e/�-$���g�b 6[f�7i���1�P�A�z����3��؇Z��'�zj^�>�Z�NH��S���+A&�� ����N&Fan�v#�lz��{��Jl��j3K�̠^���%���b�eM����mQ�N�rZ6��A�ʂ߈�U���!�]z�}�K v����Vڱ�R�q1��Դ��9����a�i+iY�(����r晀��8�h��|z@���]vA��s�cUeC���s�D���b��o���{e�x�����$1��uy�~�������)[w�B�ЧA,ѯ���=�V�,
n?2ZD�!"�-U�uNz+�����m�����<|��L6�x?�q��N����	����e
b^�=U)�R#3�s�{�1�:��U邓�b�<�ڬ���t/?'�q�q��Z\;��\����#2�IQ�k� f����S/��9Rw��ܹ��v�ۙ�!GJ��Ɩ����5�VAl���V�|��-�2�l]9[��MV����_S��<�,c�1M��:���I�*�"���h� ��X��v �Y���bO��'b
�㎇��8�\Sﶔ�} V�ǻ�c%��*�vi���Y�r*��N+0
�G2���I���ɱ��N=�����O�b���� �a��й?0"��/-�<��bA�����n�5�G��m`^����V�����1�^5��t� ��#��i���\e������Z�y3+mlu8 �\�GNQ��-�(11x'���h����Z��� �A.�S������Y�F+y�9�Q�g;<Gқ����-�|a��I����;�T:�����yX*bB��T�q��V��J�[�Y�u���9y���~,F+����W�ը\ �@-�.��Y��j�f�~�[9�/�g��_�;o��o�>���I��90A9�E���Go�]�b�+(�{����fK\�Ă;�u �Cf3�Ѯ�V��Δ+�������h��v�!��kdu�J%+@�I���pF5�4h�V���&�J<��Rt20�;_9ߨ^�<�k�1��S���z4��|��Uֱ ���g��ا������6��W�ݓ�E"�):��Bɀ��m���b���iU�����0o�1�-�ou�؈������lӨKx�y�� V�@�w&� ���2/�Hg��8bV�iG��}��e"q�X���~70�˜��%��DP���
;jWr}zz�&�����3˂�<ۙ�M�%g�]N�	�����y�󧶱\u_ُ�3E�������i�[F�O�qxe/��9��r6�S��RF�����3�?L)�cҖjV��/�ZW4�dr�������`�BïmE���H�L3ng,F'����
��k�m^��m�>�� �|�����k%RL���:���m,k_�tx�M�.X����:b������ID�A�N�O�xlȮ��m%���rս�"\�ֵ�1����7a4H!� �弇8_La`�N���l��PS1�*.�%I�t�n%����&��6�'��"���E���>�;3!:TM��)�:�3*�v9[nt,��hW� ����Ra��]v�z��(��v�%���T�IO�bد)6���hփ�]wn�Bj	� �+�ܘ�w�I�L��(dɂDQ��	�W�o��m7^}�5tW�Y�c4ww#�6vr��^�.�k�����K�˩��|��q����nj�3`Hƌ���\D>�K��Z�ҍ��;�Ҍ�����v�Ί`M�<��Ȯg�v).b٢��mբ�4��%��P������Z��G=��|m�.ݭ�z5�"N�s�*Hb�/���q�<Y�a���'��n�gd�ӝtQ����-"�hRɶYD�̓dY�����X��*E@��:ց�D��]������%]r���k����m�[A3y�D��+0xǷs�Զ,��),��(��,��8�G��_2p�J�M�k9�q�Ǚoo�/�wh��`��㫮��Q�zД��,UN�C#�����jڲ��t�*�v���"�aV�e��Ej���8�W�f[��Pn�J�ԗ��6�$��5{Gg�������>��=rݽ]�Ŏ�������΁����U��jf��������'��~��_��lO���v���tb�	mG|ܚ�J��ӼoAk�v]���먾�i촡�l?<v`ס9��_US�JcE2����_Y�r� U���I�M��?�s֓p�Wh�	:'˰�o��y`s］w�v�x���"ϐ�/vC�te�IK�]��9��l�/Z�ؐ���듫�y)����g���'�G���u-Y��Ӥ~��X0�ߧ������
'9�����pN�O.��:t�� WF��1�h0�%!�p�z��N�j�U��8����:��?�$0�Q��7J,�C���Q�� f���,*~�O>�K�hv�9!�-*Y�UTkP)�]J
ʒ���M�&��Է��R|��E����m�DA�PC��_��xa�h M�s���K|n���Tڎ����ѭ$�� ���(+K>��ݎb	����@�]����'�����^g�f
���fd�-��Ij({�Nx�a������#$�0M��TR3�jg�v��w����{+1��iM7�����gC|D "�EM�w�[�.��Wh���
�Qm�.ﻞ��z릚��U̡$�O_ �:Z����fls}�w ��O;��m�?��P�_>>`�����P���a���뒫� �nc�A�7|��֚�4��Q�gي�	d�>�NY���U�㕬�3��hL�xc���m
�.�ߩ���{��Ȥ��<����M���4mG��'�Z�����C+��xex�^�|�����?�`XC8�_D�r��w���ף1�� �W=��
-�5d�v�}���қ�rv���
J�_�c��.o��½B[�*�7��vJ�Y}5��][=p�GR�q�.ڠ�}���,�qS�H������0	���gl���N|cU�w4Fb���O����G.vz�xla��9!����ۨo�
A̅����N�3�r���b��W�&��m�_�[��U�4�|�u�\vp��n��e4�uM8aC�ǯ@e:3����|��_�h����i<M��	܂������셺�p7%�	�Ie�k�&�M#��ߢ��}��cH���i�ɈaT�B���W,�gf>�Ɩ��v6W%Q����r������;��N�����E����\�y֣���%�Irm��Ĥ3��#�Jc���EOKCw0�A�ˊߢ$����A�y��}�E����P(x�yA}�-���
2�A�D2q2r`|Uߺ�uTT����K�,<6�taW|��B����(���ҭ'�0L!ej���p�7�J�\���S/�A{|j��Gu������16C8~�g�&���K1�[&��g�����ڈ�d-��s�&���6?�k=�~S�zf�7i�bt3a��b\���/y�ē��Y>��B%�`�B�oܿ`v��v#��x�$�{6[E��M�A^��m��;��A�^+�8���:3Ȥ[�Ñ���1�=��{�g��I�[�kY���������]��H%�s�/1�o�E1�Mf�x�6b�6Y�pҥ�y��>���WD!w�+ڍ<쎄5h�e�=&H�v� ����r� �g�~g�GK���F��!kyJ�&��10[�I�+� �TKj�鼳1em�]f���3�mݤW+3&4�[��囱w����a_���Kp��#��Ǭ����^���49�w�y�X��s8�����Ԫ��@��ח�3��7��#A���Ŝ����Փ�:%b3oXp�.���c��s��5����7��h���eXh��a�C����K@��A��Ni�.�FZ@AB�n���R�AJ��x�Ywb���}=�ź�x�}�� JCB	�Ƞ=�q�&?WqS�j'[_��7���	ĸ��Rzqq*�ph����W2��X0�$c�b���ٗ��w?/��@�ӱ0I#OK�/�"���w1 �$�c���\�V�������/���m�N���cu�ξޔ��1�J��fb��	u��rf�i�0�U5/?�ST���0v���v��W&��;��6����t��XJ�<OywR�ґ��ES���]��F�;# �,c������X}��;��ECWv�J	���o �q�O.���[��("",�'�u
ĈHF�F���m�P��I�Kz"xA��}Y.�'05EVg��k��PM� ��FU�4�g9g~���p�S�b��O7�*�dy\_���G����Jb��O��#�S{�����M �M���p5D!ir�,;�5� ��L�_?C;��������5ĸ����`�_�ߓ�VU��ָg	bJ���*��w���_����}��ܛLq�V[Y�$�� fR�zx45�,��@���H�B{6 �洴^�w���g\1�,����1��{?�9�{
X�<���nZ �]�J�qU�3�tv�l)œ��bW�O�\0*�6�>i�	<k#��[>�=����ϖߌŠ�Y��	��8�J�&j��(G�&6.���#���E�a�Q!��521h�tJw��͑цwՃ^Lw8�h@��W�ڴ��%옾��^SWf8rK-�b����0 نjJt	'�A��3��d��o����}ԏN�1@�3� c!��Ό�<3�m+��1�i�J�b��dU�'�2���9����Z�M�1�a\���dӉ���7���֯�u$rb�C��,h:�Z��N��ut��ءghc�L���OJ�J�/� ���F���p��� ԫ"�3��~��L��:�Ob�K��.�%
��i�6Nz��0ݍ�f����w9 �,rm�r�ݱ�ѭA��b�8
���#�����H�fYI�'D�`�(�z��.[_ڝ�
��x
(�A,bK5xK0��\�K��z��F�5�dҥ��u�	�Kk�筼z|��U%����x�tf4�hn��禂�b�	'L>�[$�Sl!�8+�a�&�ٓ�I5�
��MǍ1�m��<����ύ��9]��]A�U�9.Ӥ`���M���rrV?��ί�C�D#�j����1�&+C�`�k't|�)S��u�6���x�9��`b�Zt���9%���i`���A�$�a&��:U�������D�[c��+��ly$J-��hA9e��b0#Cq���7b�Y�$RYa �w�0� 5�]�E�ܙ�JvD�bb\LºM�-��ƅ �ƌ,礍A��쎗�a���{L���U3��%�]���?�ؾM�uCø�p�-b��?�2E���%���ј���h�n=
��"��VtC�AlޢtW8ҁ��F������4�q層k��ӻ�T�9Z�\3��1S���0��Ay�љ���~;#�El�/�_h��{��
w�����95R�<r���ZG1
�1z�9�4��u�s�B>oTGD� Ff��T�����:+�v���"�j��@,���a��,X�tlm��	b+���LQvIHW�%��� �ʦ����"[�]�.;����Ve�!���P>��Sav��	b:M���Lެ���f��'�,oAlW1C���#��T��@�Z}�+��¿W�nf!ͨN���֑�e��OL%!m���'�Y˃��_H��@��ћ7EX:�N!3Ö�����d�L�s}��i
b8���{�����X1���cR_ҒG&x�ċ Ɯ�.��Vj�B�mƎfX�'�
�
������m�%�&�.)�'A왷a]c\��,o�;�ٮ�*{zST-�I=������|�A�	ĊI�"�S�b{��e`���߁�rKe�j��z"Ӫ'�F��W{%��ԝ��D��(�y?��i� ���1�z!�W��WW�3]���1|�Z�D���W��\}ӛ����$ �#|��5YvX.��eϾb9	y��{����{�x�ѕW�7�@��pP%�ʡ���uEb��
ĸ���"�mY��"�%m��Re	��Jl��%�ƺ1�D�X�I��>C��q�~ D-k�V�v�~b(s�V���mU���SV8dSJs� ��)nh��w�����������{)�b�x��`��%Ԑ��5�I]7y�p45����k1R�"���bWې�ZA�o2�7�L·{. v�~%�Bs���ģ;�@�qV�b�&W7�g����/�lX|k���Lj�VP>�i^��hϚ�8���N��`W��\�;0�=���1��
+�D�����3��1*�& v�G�����^a�l<�sgP.�_ā�ž]�tv��tG�؉}��X!����h�����v��{��ա2��`���R������K��$[0�^;4�jv>���~�b����_(���_atMx<��4����G&!tPSv}�B��6J��� ������ɱ�HOBO�ܾ��)����\�)�U�B��qDL��r@�t𘜷�C�0ږ�nAg�Li.�ޛb�y����~O���t�75��φ����%�'�P�f�&��&�9�[��,%c�{%�0��ZG���X'*���-����"1��M�e���D�f�x�܉�t��Q����d���m��1��ٲ����4�#�Sp{�;��2��a��}��]�_��,�����t�E�a�����C�,��V=���o|��;�f���/�����a��Y\��Es`p�nq�����`��y'���!`��С��ҹ-�4c��|���N̙Q(��om����~(�!Z)OV��:���P�tY�<�LN��X��f�#��#��ļ�O�#-�C��/[�@)F�KF�z0��ݖt�Y�>�GN���ul�O�����6�GKy�gP�Ҥ{���6�k��}��Kp��~�`\����]��
�ߩ�8/��@r0q�n��%����Gy���ܻYn=	������hٚ���y�8�\������<J;���#��� �����qT����F&o���j��T2�i��H��xI�ԑ�6'w��J�����G������׊y��|Wi9�������w;������[��/�<�����a�Q��Y�	6�p�d6PO�4�����^�U|N<���n��K�aއ�u����0z?w뱧+k�P�du�QO�����<�ĕ�Crr�jY��旍�y	j^�Ή{���!zYE���,�S!ZN�֩{���JMe���y����'��m���/E�Ps�]D\?6>��jfÅ�_��v2�A8���*e_aҾ��G��E�ܽ��V����"�}�?�e�=�PA�����z����j}��<��`F��n�~�ӈZ]yRR�)�w�n��%��:�Ւ3_��%�aN�]��Y��2�T�P�k�Փ��X�����E�uy���q�����uz�P�>ω��l|8S[\̚�@�I�]:YO���|�W��X.n�L�R���?�S>�_��|D4��� O�)}
�o�� ���\ꡦ�$&(xo��s#�k8�oOkB�c$�/˂I�{�e�I
�٠&v�J'��/�ў���I#՛�%M]�G���U<�#�Ną:(5r�|U.P���Đ���\�p���hΉM�	P#�nު�>�n��B��~�_�-Li3��w�)�4��y�*'���Ē��5���E��_s�T�(�ت����9�՛�V�[��h�W�0F�[6RbJ9�*H�e~z���Eq�u�����F��jo��F�%]9o��a�1���@�#�ɣ뾀�e�bj����[�?����{D�w��������y�2���%�5V40B/�X����Ԓ"�����ѴEB\�sQ���'��C�����u�:��A����c��M��`�R[8�zUA���� z�N©�R<����US"$��^!���Q'z���9�^�#�Ļ��?�sS�c�t�%��Pu1��{-�)���;Q�[��.>`��Q���FEQ����t1�/�YLi���ر���Gh�?w���3��;c���B���m�0􀄵�^4JK�|i;r�q�t���Et�7���v8�f��n�#�j��r5O��B��£V)AL�2�U�+�0���%w> �����o��R���ߖ?�Na����밖 6S�)	Z���z27�J�F�b����i9���� �_��6��7/��o�z��j=��[&�d7��
�J��#��-�uϕ��J�A���3�f%p�E�8T>�����h]Ĥ͌|��pt�xT:<ļwW��~��!�~����_:檻Dm�l�27���´��4@lt|��	���T|��ʄ�c�l���?,�Oc��)�;������w�7�q�iC?�`(Z���y7cQ����#G��Ǔ.1y�;?X�8R2�[@�E�5����z��c�f3�7s<�?��]��g�i9�bg�ߝ�7�0a�Cn.���O���bA�%k��� C��P�AY^���_��X湺�`��O�玖n4�0f��J�Ad��O*���i]ږ����8u��S��.�������LN�	��]1�<���$թ�[����儤��Аҥ�$Sg�Xy�.Td'�j@(� m��͑�' &;}&�h�)Q5e�܍L�C�f��CDV�����xO�PL_����{���g��ݤ��U^[&n )3���#��m<��'��R� b�[	=G��P�Bs7��{3b���p��E�@�mVk������?AL���<p�"T)t*�Ψ1Z_d�ܪ���0�.���E f��z��3�q� f�TX�x�`^�5��)<Oy��0��L.�	�4��v�0}��9b4�Fv�b��,�>#9��K!����Z �V��_�
��7���!�hb�F��W+����LǶ��X�Z V�6���HlTe$���كgp� bGt�h�I�,���!�,�2�Nb Fno{�M����z�RI��v���'�-]�K	���^�N��*��b�+J9�Ĥ��lq�f��� 9�F�WN���g�?r�G�b�&�Q�F�:�c�!���� 6!�v���j+?7���6���İ��JCĤ��vg(3a��"j?��Ӄ�h.YC���H�2\=�� 6�k|��u顊��P�N�	( �9���`QZ�� ?�TM����r�*Ea,}jV>�Tf��]1J7���F���h�6>z�|� ����/��jL� �h�ML��	b��i��!w��l�Al��K_�_���� {h*!Z`���b�/���sƔ��Qu<���bg�T�����Ԫ5�V"���@�4Q����j$r��a@[7
Dn	�(�1��5�{�>��4�����m����>�q�d�SE�I��ϳAlX����`�?����;=Ě����[QuJb��el�@LL����i�Ó[�1V�b��/4_��CW�Й�oa��,����L:��N��J�
{��\A)���y��J7,�������� ���P@�#���I�����ޓB��r�f=�_�Y���[l�U0�����pA�"	�[�+�OG���A�z��:6�������������Xgk�����p�v�S z8j�`�dbd|��w��,��ⶊ�w��
��L6X�f��)I�]A
�
֨R���5������kǗ�g/&S,�A��q{ F�KNi��8G7\<�@&T�1���4@��D/�9�?��N�\u��y��v?y�7��A�].��f5Q;P�u��M�+�Өeץ\Y�c��5�e�M�s_��v�lʔ8}�Ң�7W��Zi�L
�j=��m�AL��F2����T��p�
�\6>.���c0��{Ilv�~�H��Es �<xhȃ�Df�W_�肍��D��hC؞��aS>#��LI����ZcRT���W,	��
�i���jۢ.���C��C�Cj��'+R
}� �v:��h����gb����L���&�I�ᥓ�ae:]��&����+�9�zU���o�gK� _ٔ{�j"�-���B���!m���/���O�����}�%3��$^����WLh�=����7{��[�&��SW�O��g� ��`J�c��t����aD�aq8l�����O�Տ�� m���8���?}I���"�ir�����9e����K���'I�M��C��ѡ-��Z�g�D���;�{�E��ٱ��E�B��o�	��.<|�g����k�DL�;{�=8x�o������V'�:�Rw�P�#�����h�u\l8����1��}q���-磾�Rg{�cm̃�5	��bZs���7ow�=YX��**�7�q�kc��:�X�;��遚S�/I�����.�oz��:9Tw��5�D�u�����0�	QV���ʋM��J}��}Q��T�q�3(��0�+_�����,�t~?���E����t=`b�{������惪˔��Q�v��*��;�����vq�tO�����@���y��_��q���Ҋ5�Ժ)�qVEYgX�k�[;Ơs�&�G�M\f_v�e�?\�����Z��Fi�g�	\s�����<�ټn��;�u��3����*�]�E�:9�O�ɥ;���흳2�����)�oͥ�{�?j휱2�������fl����ھ����?��l>�-���t�IK����ݿ��p��S2#�W���hSFϓ��vϜQ0'��b߲�	
--L�sc�٧��$���"EL��uj���E���z/>��k�M���J�M ����ƽV�h��'#�:5�W����̪S"[��f��ᄨ؟���z�4ڱl�4Ol��v��5�s���O���[eH9�ǁ�WadditionalMissiles
game
hero
perml00
perml01
W?MzUx�G�I�@����Ka``����ʣ��]}�#<�����v�5S2�t( [��q�S�x��<+c����D�y�:�ɡ��j��EWn�9r�}^)L��G��}�r��g����]7"��t�����@�"�����w��}�B+���<��+��)�� =;�/�����!�*�<^HET   -   ��<�'�g0��`M<��|`��8a�h�y�^j:;�K��dL����0�����8�?�H���BET   �   =gH=0�� �5���5h���2R�6xexd6�oG�����3�\��)+W�U����<̚W������J��W-W�F��[���ZvBVt���"<m&j��Cn+pQ�<����.	��yPΒ�����` LZh���d�tm���G�f�����"*6_�b��y��^��D����U�UL� �h�-���QH,�O8��:̓Ė`dEn|�-�d�M�O�;@7������#�j� �ѿ�Jl:��gH_Dނ3�Q��?�`�l�Q�ͣ�<����(�ry�ysy!͹�FaQ�6Kݵ�R�H�R3-�[gH=`����5�g6�X��z�$�y�#�W�B^��X�#t�_*�	u���
�Cɗ�Y��sm̲�����^ـ(�3�r?�bK`>�'-��d���݌���b| �