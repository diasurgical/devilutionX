MPQ    ξ    h�  h                                                                                 �TI=H���!_�V��m�`��w�!��69,�i������A�O{]�d܄c	N�+r:a��U4QO��L���ܤ�^2�<AB�0�Đ��������,�;p&D@,BR3e$����밼FA.����a���/��-�W	�&�5dN����ڨ>q�=q��΍����/�2�hQt�-�g���CɆ'��h�Pd+4(���*������:y�͋�����nƞ}��`��>��/6p���H<�#���`�=�I?��eEȬ���*�p�
4�ALo��?@��ex�jύ (V� ��tz[����Q�j�`f҉���Mv�}A85����VҮ��%n2��l��� �!ed=�(�̕N���̥�Ù$=�K�t��1CB�Z� Pd���G��I�L�lD�)��8G����u�Nc�
�@ՃPZR�}ǔ� ��k�DR;��TQ��Ԅ<�BĤz�1�h��!_���Y� ˴H3h��Q8�1:u�!,�e?�0I?0���!&�Z|��b�[�ǂ���҆+��5W;�����5mѫ���B��|g^�z��n��������uF�hW�CM|�[���v&����=�e�~0� I�f�t�h�1�B��3��N���^^0������9"v!㩊L�� �T\)"R� �j/jK��[2���R{$���z�I�m�`ä5b��c����o�R6>�@������b'��g%	n6�6tY�$�,��N��&�q$ѝ���,Y�l*�B�	����w<��S�����`��8M�:ٛ�����@��I���r8pp���|�?m:
ܐ6L�W����&�l�Y`Ju�Ã^=����]�\�܉O�|�+�=�z ��8�H7u�Z�Q+�ڔjaPS�p#�#�*6&�-U'H���������|�&� $�g�|洌�o��1W�MZb?�j��_/���t4���'�����RO2��'���{�Т����9��[H4a��V3�^��� ���Ej��֙�y���J|wTO_����F	V��%4JE��Ӳu�ʪp�1��fr��c�A*�7c��S�F2	��&�u�
��� M�Q���6�����k
��tp|�ԇ�� .j,�G���\d���~J���#�]�����/�'�G3��>���rz��uBM�;f�i�$�mQ�v�*�:�8�50�C�?i��]�n7"y��'9D�y>�k����T.d���b�a'z�M���� ���3���k��jp8��r (%�04��r�Ж��N
U���ON�����]�wL6iF�u��ȟܹ2�^�5�������<�>:O8�Rۛ������+zc'ʶ��upʾ�H��J ���[�M�¨��&V�)��⛀q�󈽣Ođ�I\R��Be6S�
i��6��#*e�*��Ql%X_�e";#@f�QMH� J`"H;�3�rq�� ����ɖ�-DX�C�m��'D����4(���5����A�$�]����_����\y�*DSr�7���'�b�JK vP>�޸B�w��^�XIQ�bXA����Aneȱ0̀d�Z����1��t��dl<g�u��4�5��)Ĥ�M��^��S�9�����o�2yc:W����^6�{�<ү�H���3!�b�0���idPFDK��_�{OY�[�}��z��y�<ھnޕ�-�&	~���Gi����6���ƕ��W��FlH��:�Af$� ���7�]�>r�t;�۲��չ�+N��H�RSL����l~0�����Kq�2n�l=w�"VtF��r��!�!?���[�����b��|��������.��7��5D���*�3m^IF��i��8+QC?���V��ݔ�%�f�n�����e��D?�L�0iJ��b_q�Z�����s�����x�-� X�sZ��PZ5=��۸�� 6š��4I��a�^��_;�6.n��l����S�F�by�L�n��$�V"���:{�|��o��K���¾`X�B0?�2��嬪�f#ې��$IdA�G�h��*�ruZ7�F�-�D�{ݜ�O���*QY�^m��4�t����[+VT9�G�c#��4rq�09�?�
?���<�Y��hn���%U~:4@�(5��E�����wW��t���J)��aEڈ����ҽ�_��,t�3�m{�!M�J(����7�Нo�ݕj�R1�љ@���h~eV%�O������Q�b�~���<��zfLz3p�}N�'�.��f�����>�/�W�8��	^b�eB�"�2�d@���1�'�m��	���h�J�*.< ��{��c�K�*�2�IYu�.�$SJ*�q@�ٍWj�el�����ꈚJ���W�n�:���vk��U���3���䒎��EH�k�m����J/n�T�[C'�uZ�;�����f �:���3��~m�X��=ͷ��\x[LZvarm�ʴլ��sPA��b�|˗���hg�j�n�y�Cջȁ�FTށ��w"�SzXo��^>�� |h���� Vq�������4��2M,4J��[�����[a��S�&hbg�@T�	B���E��!�u�������x����<�G����QiT�5�C�.}P@a
i}s��d^
���"˯�d�TsW���3�}	�2?@�oIN�&ç��0uinx�7E���u��kP��V�������,�,�"�T9��U�?��ND���y���<8c/NQ�1��Zmy޻0�E���eN�c&�A��Pd�S·5Yf&@�(��{�9����ƏS�"q$\��ެ{0�h-Oc���P�A��H���H�<���2�z�Z�J��]�}�����(��SO&>m�* Ϭ�s�O�ρe���o�4Bo��/���2�ɯI���d�\����XQ������� D
����ytˠW]t��yU�=���$ κ�~'���_����K��%��L�v}���@�!�ю��u+��J�klmo�j�`��x��pA��pxᓤ�����Sr�xl�z���-L��؎"6V ��zB�*h#hvM�f�N�@E�#�v�9ڐf0�%�$|���#;D2��B9�ZA�D�&	U��6�k06)�5x5Q_P�уRm�w��B��G��WP�.�L�q=�d�h�܌PW�KY&��gd�d�ZOq>l�qۼ��f{U���|��2��#t�gZ�'C�Y��P��(�&�*-��ݹ��y���(��l�� (`�ǡ�Yů/�����w<�㔃����I���e \������*7
�VL�Ϭ?��`��j*A(y ۭ���|�|Q0o`^^��ɳvG\g8�̫޷3�ָ֡��m��l������!an�=�]ḬZ�c'�E$x�^d��ƅBI�# $��=�Čw�G.>)V�8�mC���:N���B�F�k��������T���2D�r��O|H�/-LƤ�*n��(������M*���|�˯>Kp��w%�L����^e��Jˣ����`&=;��N�[ +4�(���|��p��.t���o� =��#�|��=zk�|�OT�+�WǍY*�c�l���a��_Њ|�U=���ٹ�8軗0f�:������r3�۩�`r�^9�O��Y��v�WvЩ�ئŷyTw8�R��1j
����y�.�{����Y܈(@�`ޞSbd&A��:�������>��o�R���g�oB�6g��6t�9t�H��Ǵ�N{�p��1e�y�,tf9*���B�L&���iw�pS��i�8�`B�983�:T�K����=鐘�����չp�>n��"?�f�) L2�� ��&��Y���uCyή3I8ɕ\���O�#�+���z[�H8d-��3ILQ�ŵ��a��p����%{}��9gHSȻ��8A��q$�<�|�1�j�1��1M]a܅r���<�ڹ4�'A�i��R�l���������K�՝��Z9�ΰHϳ��Q�/^/]e ծ��`���_�T<$��r5T���e[	�,�%��9���[���Zʅ���2�����^�*������a0�S�u��e?� �E�����6�ض�^�k%�T��|▯#�;E�,[Fh�z���u��O���R��BU��8W���	��3�BЙ`����^��1p�c�M�-����&Kv��9�D�����C��͟WK�n����LR�Eֆ���6պ2adܒlb��z�3ּ^��*��.������;tpSUYr{��%�#�����1��N��S8ƨ���ȹw��F}���!��T��^�ɜ����&c<	�:�Q�R����:'�tc")��5V0p���H�2�J�9��u���Vz�b0�&Q�y�L�,{����O?A�q�\�[r��&�6N�vi��!���H>AF��*��l`��_U��; ����H�M� eb="�Zc���qa���C���>��JX��ˈ�'��'�j��4c���n8����A#:�]����z�x�qzT"(D��7>3>"��b+�X 1����{���J�9�tI�x�Xܒ�� �Mn�3;0�W�uQ[�F����6A^�d��,�Rˬ5�X=Ŀw��Q�.��p�/���-��:�i*��KЖe�*���l��!550%���d�fF�7wB��{jȧ�����x|�&W�<���i�:��nĀ?���9�2�о�~�'G7�AOA@����7�;�p�j ]�6]��.�vF��g�����؉Sgᙯn1�~hX��Q�-������ݱta�fr)nϊ����G�b�(꒛]R��צ��n-��4���}5�<��M���ί�^DU�tW����+l4z��V����
0U��5n��`�H���OL�%J!PPbﭔ����1�s��u�v5��^X��jZfA5/C��8��/`�6���k����lyY�_���.I+Vl@�ĺ��F͝�y]`]�)� $#}�"!�p:���|���oBZ�K�ŉ���Xj�!0Zz�2Zq[凥���yj����D5��j7 hyРۍ�7f����D��{�f���Q�m[k\�����(}4�{�TI�GG[W#�e3r�*�0�/��t
�7��7;YWW�h	K���W\~q�!@[�г�y�҄ަ�tD����)+lE�������8����X ,�#�|����J��������a�!Q�E~�1j�@����c)V���E3��Ϥ���ay�a���1iL>��x�(zD��r��ڶ�P��
���i���{�`k�"B�����q�U�m��	�I�a���.����6�Bc�n��d%�$��O� $�y�l�%����� ����p���%��ܒ��Ղݫ� ��
���א�}�	�pE#�aᨎ���l�n��7�7g�0��;1)��ur�f���u����{~h��_�m�r�\��Z��rH�`����H�� m�����k|�h�c�j�o�y4�~к���FO�����2C�n��oM#>C|��?Է�yVl*$�ހ~�̿E4(��2Ȳ�Jse�����O�[\H��\�h�@o��B�9� �I�\�p���j�G��yx<�.�5�G-R��xT�\"��Q�.x2,ae��}.�o�HT
 g"��d$�]W�t�3�*I���S@רNd^�u�ͫ2�iB��xV7��R��BiPN8��J?����,u[��q�Q9�kU�-��i�>�?¥��c�<��/��,�]Zt:��4��`!��8���>)|A0t�P��΂�f�8�(h���T������js]�\\�2ާ��U-
��<Ӻ�j��#�Xe�Bj�d�2c�b�_�e_�����}���&��(��]�N��>�p �Q�s��*��$s�]ͼܪ$�4���4{�)׶�߈��؉�םN�n�\���lߢ4׻�
Zx7�4/��ro�	xU|BN�#� ib�~"[_�س�K糧��'vX�
� �������(Q��PK���l�W#j/����Pī���X���n�X7/�Οx���z0��-'���)]�)3V��m���N#�4s��N[�Ҍ^Ⱥ��-Nf+���"����DMP�B�<Z��a�R�|��k+���_�x�M�P�e`R���ڋ��7*��y�.�c ��9g�����W��&fy�d�Q����>g�q6�^�!�2[i�i2&t�_g��4C�LŒn�SP�F[(�{�*��Gݔ�yM���F����3~�`a���t�/,�u�x�<2 X����/�I�-�e�����f�j
�?�L���?v�[ �j��(�P� ��^pWţQk�`�	k���Uv�ZM8�Zr����L��֓m���lO�����}!��=]����J�ދ�\a�$�8f�W��zDB�� �_�*�y�?G.�"8�)�_J8}Z{��UpNg���ۃ��/�s���	��%�D��|�JǏ���]���r�^yW��������?@˪T?�����v�gJ��Ce��P��]f������&�;l�VZm[������1�ī�ɨ��m��a+1�M|��z���Z���fg��(]F�^%	����������*��y�=��?��/�V�f�|��p��3�m��9^~��9���v
9�@�1�rPYT�ghRv�j��Lv՟�HY{�y�01����`��b߃���2B��O��>�f֭�x�"�]��g:c6O��t��)�bϣNvg��'_Y�4g|,�V�*�BBx�ׄ:JGwr�S���o��`�I�8N�u:���� �x���P
6����DY�p�-��	�?c-���Lm���G�&���YQ�u��L����-�\0{�O#�+�Qz���82�ϟ�pŐ�Va� pY	� �P��=�H���p���7��*$2�|�A�e=�1�qM�w�ܠz{�Uzt�>4.�{'���~�UR��IS��@�ƃ���"9�YHj&z�L�H^�� ���{�]�
M�/�����gT������k	ݿ%����������`\4TY���X�Yzl*\���zE��|NG��ɪu��z�� �����w69߬�r�k@���j������v|t,�d>�u��������ی�F6��̈����A,��e���=���=n���������)M�?:��Uy���v�6��3Ы�&C�ڟ�X(n�{�4��o� �	���!�c�u0�d�G�b}�zΛ��W���6�H�)�^�!����pn��r�N�%�6L�M/���!�N #�@��E �S�wB�vFXd:�����S^^�}��8;ǭgť<${C:E�<R�M�u���#�c������p@�H�dJ�p�Ɖ]�������&L2&�u�&��/{�5�O�t�0�\��ʴxd6I�^iW5�a�Yx�/(*\khl���_�޴;�G��(H�� ��">�7���qA��6B=��4o�D"�X�ˣ�':I[�Ey�4�Mb�	[��g+A~om]c���G��u�/��D���7�����b��� �-�_�m퍭� I�I,Xw�����un�d0CNv����4���՛|:�d�������m5m���0������	K��W��`��(�:K}�MX�б��ҥ�&�G��!U'�0��_�F�CW�n�{�W��Qk>�S���aT�<C:��d.|������'h��L���<��<�z��V��<R����з���V2���(�]�N���A�����5�Hb�%S�1���~�*/�O3�����(���"���uEt|1�r������̂���:��X���2��)|H�[��-gW5�Uш1;�ik�^?����eȸ��N+�E����V�S%�EoY윱�n��q�i�x���L�IJ���b����a%�̤�s|ar�љ����X���Z}0�IY�.�y��\�6��%��2�Z7�+p_1�l.$��lC���U F���y����h$>:`"�-�:�:Q|&?�o�,K���xiNX%D�0u"�2��b�����m�3�?&���Gh4�ۨ{�7�tϘ�DI^؜��OhQMGm(��]������VT�1�G�jI#��mr'�0�a�:�r
5�J��SxY��yh�ɜ�ʩ�~�<�@�P���5���ށ�WAGt��i��-)n�vEP�J��ҳ����w,������OJި4ApS���✾� ��1P"G@u�^ĨV۩� ����X@�<n(�l�L�h��s*=Ձ��ߞ���_������l�X���?i��[�1"�HM�����\����m�.�	#������,.�&���fc�� �C��ʨ̊�K$��gޚ�C����_9�!dJ�� � km��v��pY������c5�|�_��)���QE��G��3�&��n�IL���y
;L�.����fʓ����<�i(~c�L����-x\�?_Z��r#]'�K����_���w��2��&2hh�Шj�<y�����ȷk�FJ�G�7�s��c�
�o�~�>�`�|�,�Ru�Vg˲�9A᥇� 4C�2CYaJN�ƌ���o[W�H�	HDh��V@��oB�����������P_����f��x�fG��N	G�K*x�XT���C��.s4ta���}�f��L�
{��"�}rd_�;W3�3������@��1�H͆TYi}{x� ����n����P	���% ���Zf~,R�Ԅ<����9ONlUS;�䄮y�*9��ۘ<��-/���'�Z�'�T�E�{�9��LxAk�xP�H|�}�f�P�(#n�o%����E���c)\=0�ޢ��`�-Š�1�}���������{�4����2�oq�)ȀЅ�S��}��a9�(Kn�I�~>#�� E�s���w��8�u��β4FG��Y�鄛�?/̔�7�RȤ�I,x�8a��=�����
�g���	������~"UWgG�^u+ *~�r3��nM�K1
�w�Av3e\�;�rW�����+�g��~Ql�_fj�����Nv��͹���ȓ�+�⳧���Ix�ܾz�-�l�d>���HV�7��Ȑ���U�#����N6������o�Cf&{1���5�J'�DhB
� Z��y���$�Ԕk&z&����x�j�P��Rc����֡r,����.��p�'Vǈ��+��yW�0�&AKQd�^����>bV�q�+W���35�r772ZXtZ�g���C�_.��_�P�U(��/*#���o�sy���^��ɨK���`9�ӏe�/�:8�S�$<mNA��u����IP�]ev��	[u��g�
Ž1L "�?oVt�j��(��� ��爵2�zQ���`7կ޼'4v�x�8fDܫ�9�?l�nA���l��(��!�$='�����Yn�7�k$�a��h��OB�WN ���E�=ں!q��aj)�ĭ8gK���ANt����������e����`\KD#B��E2�����#��ˤ?��齺�~��� ��*"�˥�&��؂�,�������e���6g����&�[����[6Q���������3da㞡9�Ѽv��sqk|���zak�51ԡ%�À��Y���TP���R��1͊r�=��d�/����f�ޓ�yJ�s�3Ӄ��V!�^�T��t�=���+vH��Q��-�=T���R�7Xj�����3E�d��{}�ʋ(b���0`�bZ �5ձm
s��`�>�)o�����K�xоg��6*^ut
Ϫ��	?Nq��������_Z,�f�*��BS2��u(�w@�S�d��$`��.8i�B:JW�xI���������#�����pO<��$�R?�֣m�L���V��&�ًYq�u�0W�P")���\kz�O���+��z��8�V�Ƌ^B���k��aDp�Z��e��>b�H�UM���.6g�3$NG|�� �`��1hB�M��ܻ-��OX򐣜4i��'w��y	�R`At��*���A�o�f599WWH��G�=^�( K0���B���
�I���T ����x	g�b%e}���2���8��;�Uo���7L��T�+*�ɏ�5������I�mui=��{ ���{�6�c��c=k[������e��Ա�7,��l�p�z�m���F)���ZH�8dݢ�D��|��� gm�8j�#�o�$���Y��Mtq���A�>/_v���Ks��f��C(���M�zn�X��oE
%#�r�|��0N�d�b�j�z�#׼�D5��߲�$��|������p���rq�%�i������gwN���	i6� 6}���w�F3B��54'܊H^�Qđ��#�"��<?:���Rl�Ĕ�Oه�N�cGٲ�2�p�;WHyJ�b�������e��=�&G�.��~<��F�١�O5 G�\��
H6D��i�	��c�tϠ�iD*7�l�G_�Kb;ࢊb��HM� �ƅ"�E����q|�M������[��LXL�Y˾`'�[� Y�4�(�������DA�Ĺ]������g�f
sD�O7tn`�b�k� ����/bw��Sݭ��\I;�X����ѹnvj.0�du����<��Σ���6rd=g����X�5(|���	��G�����:_�eO�#_�:hL���C���� %8�"�!�9C0[t��Z�FUp7�&�{�Y���p�.�u�q�<��߾_�Y�>[_:�A�B�c�/*d���#�w��]���7u��$��ro+�q�Ӫ`Q�]]�#�%u��"߆�#M<�+�yi$S����d�Q~�v��q���)�#9��}f�SYt��Sr�N���b̽J-�^���S:ꍍ�����W��p�5��H�ÅQ�Gg^:���*�N�CŚ+�vȇn�V\7����1�7��n�ޡ���um�L�$�Job����̚�gV�swF��,9�^��X���Z����ig�ey,6�QE�!�)�����_���.�ԭl~ ����pF�s�y�>���$Y�"�=:��-|a�`oxOK�1*��nUX��0��e2P��=�����Q{:7o� x�h�'��.7\*p�~ZD��3��I��+1Qj�+m�ؗ���w� �}_T���G���#ד�r�\0j�hUz�
�pb����Yͥ.h?h���~'�@�^���A���\�-�qtz����j�)�ÁE`��:j��.]��\�,%�d�k��rJ9���b�!>�L{��׹1���@�TP�Y��V6ܱ�g�����ҶV���jLK���n�-0߻M�.����F�����������Vr"�К���~��g����mfl�	Q9�ז�AW.M�y��.c2�ݿ����ڳJ���*$$���b�Kٞ����	&�<Êf�ޚ�������Pk��t���@�7�ː�����[�E��������n���l��Ȧ9Q;gwM�k��f�}I������~^A1�v.��[�\��dZ�Ɗr�����U�D�����ҍ
���uh�]Pj��T�b��&��R?FE��ޒf5���[���oC�T>xK�|f���SVb�=��!ĥBw?4^h2�
J)q��B���[R@��dSCh�k7@�7_Bؿ��Ꮡ�?���B��Kb��$�x�h$�臆G#�NS�TO����.nVa-�}����px
�;"\Rd�KW�Ǭ3��<�C��@M��j�:'�a��i��Mx�E����Վ�R�P�]��5�)��5S.,�e���p	�7�9�0�UiJ䟓|�5����s�<0��/�"(�Z*5�f�q�.����A��mP5��x $f7��(�[����-���� ����\� ޝ�?A�-�o��LhP�}���&έ#xpn㕢32����l�ța���@}�ca���(�	�D]�>~_�  ��s�cu����� �y4����C�������l����$ƣ�s6���2��j
w�Ȫ栨��vyU2�p�U} �~�8�m��)�8KLA(��'vU��v�R�J��T������{�Zl���j%+L�w��!��AQ0���1�8J���x��z&�i-� qɟ?��_<uV�s��#L��[|#�7�JN�����^�
5qf!��5����D��B��QZ�(̜��ʏ���k!L���}xf��P��QR�T	����N�(-�.�}=Ƃ�'�����-j�W
�&=�d:�/�+m[>]�Bq�o��YP�`�$�25�t�N�g+*wC��S�$�PP�(��)*����J.'y���{lĦ����t`ס�Ӫ�/"���.��<����T�����I�ހe1ד�$���\6�
�[�L[{\?���Q�j;|(B.� ,P�f��7Q�;@`��,޷�NvX�Y8!N
�/)B�C�I5���l�'����W!rJ%=ӻ��?b���3��$)Q5�G��D6BZ�� <#��`��5@�ث)J%8�������N���s+s�����iY�l�a��%D���@�R�@n}Yd��ԢTz�:������$�ˠ����=YF���K��@e�$15�L��͎��&N�\���i[Qy���������!\Y�9���% ����.H-|�V�z�ܯ����ܿ�^�&�Ts��橰Ghp��ʷ���*=�9Z�j���C�f�`���g�.��3�,��(�^�K��pa�G��v ���=G��&T�%�Rl�=j�1)��ɟ�1�{����?U�Y�`/M�b՞�i�걨�1��PU>���c嘘����g�6V�tE�̘d�Nl�x��b��x�,Ŗ*�B.Պ��&_w�S��0�%�1`sq�8��:�Ր�S�����K��g׮���p
kP�?�2?Y��H��L��=��^5&��ZY��ut�%�A��&Z�T�\��}OY�+��zl��8��W�g����Fa<<\p����
l���'H�%����/��"��c$�|m|RgW�[��1ñRMF��־��KE��kH+4�'?�tDR��/����E0����A��9�P�H�k��B�^@M �ݓ��f� D7����6(T�e��x�	�% y0��$��C�H���A���U�O�*����2E���%���\uD���y� ����v��6�K���u|kv0��`bݖ@�n��J�,,�k����i@��D���������כ0ʳ3gqV��*Ѝ�'/��ԿAMO�N�UP��c�v���:��!;CC����xn�Ux�����݆��׭��닒d-�bsuz��O���¯l��[���Ǚ�ln\p��$r��0%b�$��k���N�8M�d�.���~�$w80�F@@�p���%�I^�E�� ��b<Z��:;^�RG1��ۇE�c]�F��p���H)��J'�|��9d��3��&B&��+H2�]����-iO���-\>�X��+�6?M�i�����F��*��l--_&ا; ���
�H* �(�"4��՟ZWq��9�lY�������X"���k�'0
'��X�4$"�? ��:A4:f]٣$��'��������D?�R7<��b<� b?,�J���c�8��/)I=LFX�����n�5�0��������~�w�R�d�
=�XcN/5�=����'ڿ�Cu�- ^��A:�m���Ѻ��cOқ����(<!�k�0��UX�F��s��{��}�G�/�	�
�׮�<y㼾Z�����H��]p��'��v�������՚�2��R�h�-]��\��ۙV]8���`��G���1u��U�4�S�1Y�ߋv~�-���X""�����^�]Et��r�� ��6p�����;ܛN�Z�谛��y��9E�#�_5{�'�����B�^5B��┸�ު+��ۇ�KV7;���M���^�n�䧡�y�0�La�J�.b�Z��FV�(dsrK��΀�0X���Zs%\�ܵ���h� �`6�!�|�_�Ќ��/�_'LS.�١l��fċ1yF�yn��Z $t�"�NV:{zZ|�u#o2gK��D�.��X���0��+2���V�R<ѐi��5h!�{Ȉh����a7�`x��iD��#�L2��'Q�#�m���������~.T���G,�a#�Z�rݽg0%%�p#H
+=ƽs�bY}�h�&�����~��*@�[����\����7Ӫ��t���}��)$��E���U�}ҩ����,`��M �-0J���u��<�(�����4�1���@STH�T��V�.�v�'� D��N�1��]T���iL���i���\ #��:j��@;��α�u���Q��"Syh�PO��e���mAʚ	�5���6��.����g�cM�ѿ������ ��$�8��]�8���-�Q�քWF���蚶�:�C�
Ϧf6��^��;+��I���ߒz�UE�C��Y�c�\��n�h���'�a�;�N���Auf���&#����~Y���p��ͣƔ\�Z	��r٦D��-S����B�贅����h�
�j�;/9r�/����ХF@����;W�ce���o���>SVL|T�`Ԉ��V]mĉ�!'���4y�729�J'ڌG�� %�[M����~�hN�@��vB�	���B;�����F���I�{�xm����KG�$�.��T��*�y=�.i�av� }_���
q"7�!d���Wi�E3�����0�@��J�M��<�}i�"4x'����z؎S*"P ��P9����`,�d�r  }ڝ93.Uɶ�亘G�[��q+�<kEI/��F�Z�b��^�𱑑�s=����A�N�P�3��sY�f��(��p���]�uS���{�~\s�ޘˋ�G�-;^�g.K���:Ҵ��	��D�q�2t�h��ȶ?�I�}j����"(��b�?�G>�8� ��!s 7�m#��[�44|H���b�:�w�._�*�H}�����+I�s�C��
k���e7��eU���{U���U :S~�?(�w��x�Kg��m��v�d𴱭�����������6��l�Ϥj�vȂR��\ڿ��.���-��i��?��x�"�z�)�-�f��`�����V�ϔ�~'i��#�.�u,rN�Ü�����f�-��շ����D��B +�Z���&E�M�k>��p
x!�P��fRY̼k`+�萎�öE.�:���Pv��HI�W��#&�N{du�n��a�>XF�qG��R��kY�h2m2�MtЦ�gƉ�C��4���P�(;�*J��%�*y�}t��F��ě�D�N`�*��ŅY/�a��	��<�
p�������I�#e���?Qz��$N
{ML��i?G�}L�&j�N�(��� G���:���9Q�d`m��޲�v��8�w��J|`�(g�$I1Y�l ����O!��=�p�����O�e��=S$d�4М���YiB��y �b7�{^ڰ6����)B�8N೶���N*�&.�t��������G���֜4DY��;h���xp8�v��1��*�h��9Wd�`G�˛VD�2���9İ�҅��չe���p��7,��9&����=�[l�J���r��\-�2���1��rm���>�|�$�zWnn��v�����'�OJG�
���R����h��=a�٥t�'_f���/�e���3	�'�LP^�b���by���v�]�QJ�ţ�T�NR���jv�Ȭ�a���W{�I�Awh�`J�\bP\oD�/���$� `�>�_־c{�S�a�zgg��M6�m�t�ը�3��Ngq3�8�v�e�B,��}*n�B	����D�wC�S�vk��Y�`.548�4�:@t�.��)ΰ�!����,�U� pŹ��Z�:?ԉ�#ͧL+���&�fY'�u/ĸ�R�[
��\��O��|+��z��t8P ��c8��!Aaw�hp*^^�ϳ��
hH?��$�j�m�$���|�cF�V��1A�M�R����Z$�F�4�a�'��&o��R�+z(�`�b�7E:��W9ͻMH;>��=��^�2l �1l��r��{מּ��/�q��TVS���i�	�(%۔5�9Ͳv�����w��m}��JN�*m �����h��?.xu�R+� T�Ϟq
T6J��J�k��I���s����'�:,ǀѮfE{�#�����ό#㤊.�ʢ��c��S�6��.�y������Bn��O�M*5����t��v�r�"����C^��CA#n~rp��m@�P���ڹ2�զ��dH'xb�z_���������2�'W�p��8rg��%=/9��9VН�N�����v�3�Xw�~fF�]������c^�Y\�I����aF<u��:��tR"HN�&�����c�����pq/�HDwzJ�C�W�y�tS���ʰ&=�S��1����^O+?1\->\y���Imx6:��ihͅ��f���>!*�h�lL2j_���;
@-�J�H�8� Ѫn"����z�Hq��Y�){���i�U�X�׼���,'����x�4O? �ڂB�A��r]�����%�](_��~Dz��7�)��yb�̎ ��e�m�ހ�����Ix}1XH5F�쉖n,!�0t�_��I3�2���Y��-�2dsξ�H�d05�4�+��=M�ښNN�͑����C�:���~>�h���؟V!�!0��>�P%�F)�.�v{��*�z����6<�1�U����i���ԜxJS�%EF�}CI��^��E,�-�����j/��!W�V�]V*��;l�؆�_y����zOS���Z?�~w3T� Nd�g(���3we�ɀt͢`r���h�3=H���$�I���C�ҨZ(��T�Z���%5V`��9���:^�^0ц��P���+�87��vV_����^�m�vn�>͡z$J��օL*�%Jgb[)��� b��wsmpQ��d��X	C�Z�O}�V���M~��-6�Y�נ���g��a%_���.���l��&�9F���y�	!�f9$�1K";:VJ�|�@:o�dWK�;��كXV��0���2Fߎ���?��1�m80�Ϧ�8he������7R��`�D�����:��CQ ��mG�c�����C~Y��T5�G�eB#�A�r8�30�-��
�)v�NgYCthu��_~ݰ�@Gx(��
����t�B��xDz)ܗE����p���$B|�c�>,������u�J��r��W��ǖ���D1�@�s��O��V��1j,�;����]�ͅ���L����dd�����Y{��˪<���v�	�����LO�"�A��#�,�F�}O�mH�	�n[oP���	.�}�"m�ch������;C$Z�X;b�T�~��K�rg��\?���Y�~�A�Y��h��t�����P�	�ZzE��7���2n�=f"Ih��;�E#�a�f[�ˤa���:�v~Taα˔o�^QY\��hZ��r�{������zf��X��C��W[h���ju�l
�ѹj��Ȉ��F;��H1٠y��no9Q@>.�/|�R��#�VXnG�JB
���I4��d2��J�����D���2[H����!h	��@�3�B�Z���Ö�HXf�!j�Ym�w�Rx(�*�ZYG�{	��T�9����.d�ta�O�}m
1=
��i"��d��W�V3�!���)@�G�Й����z(i.�.x�����rw��!�P:�ks���,�y���x�F9`U�U�$��ս��+$��L{<�U/U6�$kZ௴�W��̡��$�G��tA-�Pk���n�Bf�Y�(TC�������C����I�\:ޓ����F-�l��n�sP�ҏ�>Dv��GS�`�2�z�N������	~}EKה(��:�6>42G v$�s�`��bo���@ܖ��4������镨bpޮ�7�o����Y+��@�g�l�
���� Z����q�l�*U�S�v� �@Q~�B�؟>�K����WvĔ2���(P$�� (�<&����l�7�j�0�-�ė�w,蓋���ĸe��|�x�u�z�8-��)��^ؕ�V�K���"ð�)�#�l��- N���J9��@�tf������{�/D�4B{w�Z���M}���/�kPպ�[dx܀yP��R�c�F�=�#��^`.�K�8k�~o�cH4W x�&Ҁ(d�F¼avE>S�mq�� ��C��_�2�t�ga	�C�XҒ�vP���(5u*�� ~y99�/1>������`M���E/%����<�������IaGe� �Z��R3�
V�2Lэ?�PRG��j��(��� b\\���(!QWd=`��ޭ�7v�f8����e��8����|����l�4���w�!(}�=IE��7��ʉ���$�ak�m��Bu �ؖr��+q�����)}�P8�LL���_N����������_D�"��mwD�h��63�����$ͤ�V�J���C�3�t2%����˖�7��س:���꧲�ea����ǂ��me&}M�B�v[��$��n��MIėa5K���]"��C�U�|	-z�Y��s��R�ǔ��JA��esA�����]e�㫊=<1���{R�� �f������C��43$p��Ǘ�^���%u��}snv�����v]�^oT�cVRb��jQ�x�8+�5��{%rʜΛ��M�`ea�b�9�|��#L����>�2���Q�U���g�6���t�&��y!Nb_ʁ�T� 
M,�V�*���B�z��&�Gw��S�/���1�`��8���:�2��	�A�dk����O�����p�(q�uAk?O���LYq̤'��&�f�Y�J/u� �����\8pO�DL+���z"508����.���pa��hp�l��w�O��H�$4�*͍��>�HR�$�FJ|����Q=�1y�M�")��2�A��!��4�p'H.bj�Rqpg5*��{����Q���_9GGH�0�8�D^�7 |�^��:�����"���!�T���z�	x�K%�о�!�}������ {�F��E**�{]�f�����º��u���f�O �+�l�6�8��Fk�"��V�V���b�z,b�a���~��w_>�>W�c���-u��#�)�g'�D��l�]�6��$�Mǣ����-rv�zA\)�З �Cy����ynY��� F8�c{���a���g�ag]dc\�bi�dz:{1�C�گ�_�w$ڍb���_.pڵ4r�E%½�9(m�88�N��g����1�N��w.�#Fě�����[�^��ґ�H��S�<��.:1��R�0�a���{�/c	���mp,��H_XgJ��2#��b}�i�&8�p��:���B��*��O��H7l?\�������65W�i�F��MB�Ŕ���*�RWl�W�_\Q�;�\�s��H~� �L�"*�B�Udjq-���`U�� ����)X}���f?'&K#���q4�z2�u%���A��]OE�����أ��x�D�7�7E71	COb� ��;��+��YG��;rI�ΰX㭯��/n�,L0/iK�������7�4h� d�x攟��5Y!�FU�¸���u:)�4�6���e�:y��9�U��Iґ��6a!A00,AJ�KFf���i{��_�=uQ��%e�M��<�?�PN��O!�knԜ�DG�����X0$�(�#�.�u�(�'l У����Ūъ�]�����Z}�����YM���3{S���~Rv�;��X͛�$�Ɏ�H��Ut�]�r���C�;�n�3�/���D�4�W���~�o3��M51���tB��ՙZ^+�7�;�a�tr+��ڇu++V�u�1����cn�N�������MLE9�J��b6W��ʳ�8+sh�>�=k���~�X$�;Zi�*|�R�#��6��6�!M�2�+�Fb �\_W�.�Cl/a����F���y$Dr���$�n�"���:1:�|,�oI�K����>�Xǜ0�p2�
���k ����*�+*z�1��h ���7�-�;�7D5����c��4Q{z�m������4�Tp�QGb�Z#�H�r�j�0�h6��=
!6r�)�Y~�Eh��1�~8��@�8�1^$�G���@uC
�tK���s�)��E<W�ԋG�ҟ��>��,��J��x�݀JJ��-�;�r��∴&��N�1<C@��`�J� VG3U�Gu�VN��D<T�����X.dLS$�_b(A�	~�7���'B�Qx�D.j�����G"	*�����GI0���m���	�_
�=�杁.^�����_c�p2��w�k.Q�v� $��O�S��ٯ���Ƅ�����e�lzHܹs����ԫ��j���hSi�$Βp
EjaA�ϱd���n�2h}ݨ��8>;�\ڗ�f6��������~O!��&T@��A\�fZ�6�r�p"�7.�����Ҟi��I4h	��j�j�X������#��F6&�ޣF���Ɲ��+o�,�>	̂|��eԾk_VS�Ɖ��m�s�4�Q�2/3MJ��-���eV��[C�'�u5hď�@��Bx�S�gd���格���Ͷ҇�x�-T�9�G�}��8�T ���z$._|-a,�}�Y�L�;
g�8"협dKb>W���3�k͂T�_@~����ғ���ii�=x]s������	9>P�Æ�4|�����^,>�Ä��us��9���U?����6���'��<��/�+ҔZ;@p!��щ�=���AW+P�n�i+�fH�(烛����k0�ƱFR��$\�2�ގ3xR�S-��������f�j�c�SI��o�2*i`�	:�����?�} �%M��(���5��>�K� 1is8���c�<����ѷ�4����-���M+��R|=�>�v��S��$v�ߩC/��
!e��۴E���6�甅U�:�J�� p�~	B����Z$K��3�c�v��Ĵ'$�����D���ݬ��l��j�m��zm��f��J8���8��3��x2x�z���-n���P��0v�V����4>�����#
ˉkO�N�E錅���ۯJfW�FB:�6�yD�}�B��Zc���������Ik�r�&ͧx�+P+*�ROh!�@�^uI��)].��ƓI�ƥ��~g-W{z�&���d��)����>N��q��y��ˡ�M�^�S2ƲtF��g��?C��+�5i�P�;�(P�*[!���!yt�Q��;k�`\���"`����%�/�{��#�<YGo�%����]I�W�ebr,�uǟ��a"
1��LGA?}1?B�jL�(sj^ }f����ѸQ�(�`�C�ިcvi28R+-�����������ϗ�lV�z��R!�Fg=:G�R��E���$�;������CBki� mB�ر�ڦ���iI�)��8��|����N�����iW�ڭ;��q��L]�D�`��1��Q���g�7D���P�����-:��Tˑ�����n[��"��~,pe<�J揚m�ю��&_���t�[��
��(���/CЃ㞍���(�W�_�K|$!�zM�o��t�ԍ�0�/O�EX���i-�xMd�3V(�^Ȭ=���m�]f��r����__�3?TW�B�8^[�=�`����tv�;�����G�T3�R�A6j,�8�sh͟�O{�6��E�a`��bF7��(K�Yk��V�y>�u?�t�h��B��0g�d<6���t�[��i4N]m=��!��ۂ�,�*uu�B�}��a�iwy{S�բ6*[`�J8�
�:6C��@z�����W����+���p;��㐧�?ʼ/�^L��!���&��0Yݘ u��*�j$OZ n\W��O*�s+�3�z}��8�)�2�j.�;�׼�a�z]p`�������3�H�T��E����#�W$:��|#���L�1Կ�Mw�#�'��ڼ�����4U�p'��Ue�R�j��o���b�-f5��4�9C�HqC�3]�^Q]0 7���#A�q�\�v}����/T�.e�Ы�	�.�%Q,̴<�6�lR�ʧ��[����.��@&C*#���!���Š�53u�@j�~� �[��gx6 ߼��j�k�����g���jԝp�,�ݖ�\I���}J�2\��Y롊$i�Z���hW��lM��$�����[�xL]�E��M�xf��,����v��J�P��R}C����9||n4�[>�vc^��}���D	�)d~�.b䌎z���~�d�=�ˋ5<��ߧ���-p��r]`�%�t��t6����N�s��uJ��D�i��w�{�F����!�J��V�^��d��֭��<���:���R�9��� �=cQ�WlVp碭HzY�J}4��͜��-���&3��<dT���Z�E��O!���0\��ӴP�60-i���"�k�|�.*�\;l _�=	;  (��(H9� �"��s�0�qhb6�=����kh�6�X8�0�*'��S���4�ո��ܕDAEZ�]
�.����S?v�JD�7�d}$!bM�* �
������-��[��I�?�X~F1����n�W�0��ڣ�(��z��g�d��j�;t�r5C��a���3&��PF�&���I����:ԑ=��wy�8��������[!|��0�ήFF�a��E_{׸�����*�&<JQ�K&����&1���^��ز3=/�c���Ʉw�#A_cn,�^�C����L3�]ɥq����2�����eS	�A�Pm~-��v���R�]k����?($t9�rߊ �̩���ʭ��?�����!���怊�����65��ѯ��p�^&O$����/�s+{Ƈ���V��l���R�n�R,�0���a��L`�J-{b'������\sc�o��J(X?1dZ�dW���U��+�6�Q�΍���}w&<_��.k��lja��\��F���y����n$��%"�h:J�|M7do�)�K����?�2X��0�J�2<V1�&1�M�:�&� ��yrh�V;�/;{7H��V�Dp�k����mQ�U�m�3��1���
�cT��<G���#�or�p0V:�ޤ
�b����Y��Jh�"��#~��@�-�LR� �%�ȧ�~L�t�5�n�%)5u�E�>tԦ&������,~���dJ�e�m�������b�g�1w��@$��E#-V���E�q 翔��5����_L���Z�����9KX�#�F�2˧�,�����F5o�BM"d2���*��b�!�s�mңl	=A��q��Q.��𘊸c�枿��r�F��̱+�$���Ni�
La������	��R�ϚG���s�wj���ܬ�*w-�#f�?fa���EE ��
L��-�!n�G�ؑ�Ȓx�;ӓ�W1Cfe��ײ��pg�~Jܱ�31���N\5�Zz�+rj�ٴrރ���ԃ�b��s��͞Qh$ҿjk�3����S�Ⱦ��F1����{����&��o/(�>�6F|���Y��VN�A� �P�.fd4�4�2�y&J�0��ƪ��[>�����h�"@��B�]��B%^����W=��h�->�x��A�T�LGZ����T;觬JI�.ZBa��Z}�f�gA�
�t"ȯ1d�T�W:��3�������@9W����D���ݭi��`x�]���dp�P�(áG^�^�F�,y�A�C�n��9�1U�_h�hY�!�M<i/�b��Z�������"b� �`��A�I�P����d�Qf���(ʪӛ�����ƌ�����\D��މ��� -l�	��@,�i>�E�8����ぞ#2�w|�����qʺR(}���5�(R0�(>�s ��]sS����Av��#�4M�����KQ9�Z�mc���|���m��_���D@	��k(
|�Ȗ/�|��b��U����� �u~��9���*�K�ur��O�vzT��b�^�ǎ�,<��Ж�ghl*hOjƂ���ݯ���������z���p�Bx)|�z�8-IX#ɋ����V��yW�GW�#%I�搠N}����1�v�Xf�ꙡ���߇D��hBqpZ>�7�Ë��k�k��^�xR��PF~R��_�T3�����.�1I��é���[����W��z&�D�d&������>I�	qXp���W�w0��2��&t�ozg�h�C��A��{ZP<�3(k�*�~ݶ�y�g��efp���U`Ä8�&/���� <����!z�8I�e����>�H��
�LG ?2D=��j���(.i� ���R�V�y� Q�`>�QޣBv��s8�k��_�.v�ֵD�
� l��k�ث]!�/�=�N��m/t��ȃ�~:7$6��t��X�B�}; (�4�̀�!F��Ds)��8�E���N;�_S�(��Us߮���m�D*x�,)���W�ipF�R���@�����m��H��1o�ˌx풺�)���	{�����e�3!�������&��>�@�[�`񷅛���a�k����у���|?O?z�Ⲓ|�I��������@����ٰ3/��No3��=�P�V�\��=�f��P�@���3ZX�����^6g����y����v�ީb/t��>�T4"�RXLj���š�k��{�4��R�b�E3H`���b�T!�� ���6��N�>��I��J���P"�iAg��e6qut1���NX���I����,1�6*�(�B��2��_ w\�S���Bi`_@8�:���C��	���M߷ծf�p�e"�-D?E����L�y+�]�&�d�Y8�u`
6F1���5$�\�V�O�1�+��Pz�GG8��M2���Ų��a(%Fp�����s��)Hp��`;�ʊ��%�$u�w|���G��1/��M2�B�B�~�7[���G4�B�'~�`p,R'�������&坭_9~�6Hv��.��^��� �p�+Z�챖�Q�Q�"�T'̪���}	.�%�]�W����wʂ����>7q�;B�*~�\�܍x���°��u���j� %ω�b_M6[�3�{�!k�6�LT ������gv,��}�W���4oc��xȌt����9ڢ5�[�YN���������[�����	M�J9�A�Y�Evwv����'�F�C��I+n�y��V4���됣�C�����8d�&6b_��z�S���B��Tn�0�C}�XѐpV�r��	%�G��d��n�N�s������6%w$*�Fzw�\Fܑ�B^�U�ZS���<��:'�:R�bŔ�d뇱-c�AŲ��Rp��-H�zJ�x����%ᱨ��&.�����ʀI��`��O����I\*3���6+��iy���!h�bQ�m*~�/l��_�J�;����)�lH�x� "�" �P��=q����/2����f wX���E�'P�g�64 Q����7�˪A�O�]�f��7H,���>Q�XD+$�7{���$�b�͸ N.\��Q�O4 �6��I)�kX���ݍ�n=��0���2����=���p�dDٔ抭��g�5τ8�|'.®�|�+rOac�l�x�
	�:/3���D��S4�҇j�i�F!�t0bʮAL�F.�_�Y{'Rb�3���u	 ���<�!�F�����@�ɘ'��]��jj��W1�dT1�S����T4��0�����]�}��LU4������9�� �S$����B~\j���?��j�
�C�D�����vt41r�c��-H��ǿe���:�~�T~9����ߋ���5犆��
O�q^!>M��[/�ꅔ+)L��k�:V��~�����>9En�f������L{��J~l�b�UϤ2�3�n��s^����&���XZ�Z_�)2�0��-8�l�"6��	��.x����6��_�1.F-Sl��B���F���y�ՕFWo$�H?"~�:�y.|�bwo�8K�oG��iX�H�0�T2��d�ҁ>U	��!læ�Ikh�2N�J��7�z��FD����g�W�Q1Qmx�d�L������1�T��G��4#���rI�0,��T
�N�ߚ�Y�$hFa��5�~�D#@x��gf�{Vޣ. ���t�߿�i{5)��E�F���%�ҕ�����,L����8��BJ �h� 	�nc�~�J�B�}1�2@��Y�@�V��bcӋ���:��^�m���LR��U����s��ܬ>{`������e�*���Q�=
z"�Z��<^5�}��m��}	x�$@2���%�.;��SI�c�|3�7��! ����$+'ȦI�F�e���=:C�Ê��͎
�"�/���ԫ�FK�� ����F�Z�\�f�pE �^�E6����n�|�3f*�M��;�����k�f�x��8~Eͱ�2B͏�\P�ZZ�!BrE�����Q�K�\��Y��T�u���h?�Oj����й/��Y�F,2�Yџ�O�+�]o�C>��y|@�;����VI1��[c����74�72%�Jp>3�����[9ܿ�+l�h:�7@,�eBn��ʑ����$��@���xYQ��o�2G�Vz�0�Tv�y��7�.U�a���}K�Y�q
]a"���d�fxW�GZ3�e��
"�@��!GV�֘ͨ��i�חx��w�������Pkk�ü�/r<#�|�o,�����i��9q|�U�-�&�D�=l��J.<WRq/&�p	�|Z�W�����"��;��A͇P<�8�_}�f��}(����hn�a�2�gBi�:\��ބ��M-'Y��ӆǺ�B� ���z��|�2�X���"�5��}֖�Ô�(�5;�+�+>E�� �R�sn�N�Y��Z}�Gl�4�N��״��$�����jq�4g(�k�o�@���\{���
ף��Q��/n����?Uy����$ �w�~���q���OZK�Ry�YКvU�ٴ����ݎ�r�M���"�elE0j���ω�Hs=�H���|�����O�+��xD/�z���-$>���%��f��V�g��ԑ�F#@��a�NXG����H���f����.���1ZD
p�B��Z���Bw���4kF����x�:Pa��RE���;���԰/U.�n��I�
�<U����Wq߯&c֐daN5�2t>D��q�wˍ>�1��HT��2|zt�G5g2H�C�q��fP��(�O�*�ݑuYy�J� �M�|���kw`~���1F�/�/%�u)�<�?�[�Y�nIrH�e�y�������'
�PEL�i?�Ra8̂j\�(�v �ށ�`7�T��Q `�:�ޞAXvϚ8�^n��@�z�֐آE��l�����u�!99I=z�g̈�<�;f�Yyc$PPL<c����B!�� 㡑��7 ڜ����q).Ĩ8�R���U�N�ba�C�f��X/��{��xDů��'T��$Fi�mw��,����%�`��Fˇn�HH������$�~�t�e�z�\���W��P�&�w�s,�[��� bS�ު��H��Ut���x���a��Y�|Z�zC�!�W֚�Mo�e�-�;���v�E��0��i���Ta�=͔VّQ 蓌f�ʊ��y��Xg3u|'�8.^����kb�N@�v�������ŏV�TO1�R��j�:��B����{��ʭ��� �R`���b<�_��&��[����*>�[�*-V�?~�OgxU[6L�tlb�̟	�NS鷁���Q��,LgD*k�ZBu����
w��?S�/��z�`�p8a�:,.��������Nڛ���pIp�4�����?�o~�p1L
.��HI&��Y��Cuk�Q�?m�h�\��O`��+�z3�8<ӌh�a$�ōz�ac�"p��e��"��`�jH+@�{��ٿJ$�f,|Y���B�1���M��]!ڲ���`�4�"'�e[KR���f[���!��#a���V9��,H�Ȧ�)�	^u ����8S[�gݼ�,�=�]�yT���ms	�/�%�Cs�r���bc�]eѼ���_t�6~�*�M�藴��9��+t�u�Bwy �b��]f�6��j�6�5k�}���`ǖ����2,3���R��Ꮐ\���㌏s?�������{�ע ��88Dg��v٘��B�;�M�<�|���J�v�R1m���Ș�Cʺ��/7�n�%2�ю ��L���^��IՒ��d��b��Fz��\���t�s�� ڞ:�:Xp+֙rSGN%�:���j�	�N����+���bC��yw���FU)��k��,8�^��ݑ�"p���k<�5�:���R�����q�L�c��u��p]�qH���Js�/�Ô �`P
�:e9&)���!����{�FO=���\e�괵�z6&�Jiԣz�~A�zsrhl*Y�3l8�'_-w�;������H�#� =�!"������q�b�s�4�|aW���}X���`�''���B84;���F�9�!�A�df]�'*�R T�I�a,��Df�/7 ��E�b� 	z2�����Z����Id��X��|��y�n�0`��MB���,�ś��$d���dT*��5��lė���)P����*l�����:��D�j1m�n�M�r~�D�!!�FP0�->�<��Fw{X{B�/׮�P�����$<�:��A6X�`4������������?��C����D���h�v��B�']u���HNb톨W#^����WS?��FM~��Q��)�Ɩ/ɟ��OMt9O�r���{&��o� �8�5�M�A�F#����A��I�5��%��G^M��LJ6��?y+D=v��5V~.��⩪��?:n������M��)�L�m�J��?bǤs�m�a�	 tsYD��Nؼ����Xu�MZ�9{~���b���O6���C�N�w�Qj�_��W.!�7l���ĒWnF���y5��=�$�� "�P�:���|í�oo�K�u���.bXB�102;�22M��_��y�9�p#T=b�B:�hQ.��e`7>QW́&D�f��S����4Q�l�m3!��gP6� 	�łT!�/G3t�#��r���0�=��PK
�/����Y/��h���g�~I�@3+³����g�~�-�0rt���dx�)��Emnn��D!�����g,��T�|���J[|�^����x���<ߕ�1�@Z2�;)�VX�9�苧��絥�9e<�	�RL���P�R����ŬY[b�(r7��`����| ,�83�"�����L��J�iI@m�	����}���.o��(Vc�2�}���Ȉ�'�+$�rئDw`��hD���Ȅ�+HS�����j�2ϭ�W���E���丙��u^����EE�������c�n{�V�Zk�XP;	b0�M�3fǘ��M]N��`T~@!Z�7Rs�J��\kNQZp�r ش�S�愜��D$ү葐C�XhZL�ja�+v�p�V*���}QF'�
޴F��
�dF��o%(>�l|{�Tԏt$VD�,�������4 [h2�f�JK��n��' �[4(���7`h���@G�EB��t���4	���8D��T��
.xi�~`Gsgu�:T� ��F].P�a=M}����
��."~=Bd��Wp�K3���en@���<Qy��̓�si�x.�*����?�P&�z�כ��9��W�@,�6ڄyn[d�B9�uUp�A��������_<���/�`W�:ZL%sqza�8"������A�Pׯ��ZVQfY{�(@���,����k��B��5��\z�����c�:-�爼�슺_6r��[�0��v��w\�2;���:'�=h�ʰ}��;��(��M�&ي>�W  b��s���Ԡ-�5��܂�(4� ����?�z\����ג�qS�F������z�����/
2s���J�u�X5�UT�Z��6� A{~��h�k�؋�`K�OH��pIv0�\���x��ˎ��������ݓ�l`�j���*�ă)?��b��w��0:���+�x_z�h-�C]�����~V�{��EPl��p#[�E�s�N3��6�-�JfL@�W��g��D%�Bg�Z�oΜ9�Tj�k�r�7�xȳ�P|��R���B����F.��7Ƥ�k���X�τIW�Aq&>�~d�;ټ�;>?�q�����/�+	�U�2Wi�t�?$g�G�C�d��F �P���(��m*���l}�y%N����:��1`9���L��/s\�P��<
U���1���I���e�-j����>��
®kL�2[?N��3 `j]/I(��� ��KH:D�/��QC5�`t�ޙ`�vź8�(5��A�$���k�G���l'�U��_�!�b�=5��̣�mʶ���4�$�����Z�֢�B|h ����}������)i	�8U?����N��e�˛�^O��K^+��0|���D`D�"�>�b���;Ф����6}޺�}��`�q�gԂ˂���J؟}�?�A���eͅU�b�>����1�&p�0�.8�[�F޷{H���`Lă#b����~Mx�9W��.|u�z�%��27��>ɜ� �
�6]a��r��R=��"����=��,��ط�.��f�!���|���3��+����^�ޜ�>��Yv���h��J��Tj`�RNj��٬$�����7{��,�l�����`�	�b��I��\�
��'�>���օ/-���L5T�g��6'št�d�:$!NNW���I��_,gW:*��BPF'���wJG�S�SV�G�`��I8&<�:�lb�u
��P|�(�՟}��kpl#d�ᙽ?;�gj)LLE[����&��#Y�Cuu��l���A���S\�FO���+��Ez���8��C�0����h��a���p1T���`���H棡��)���y�$�[�|�2��==�1���M����x�k�-�f��u4#�'���VF�R��!e��~?���c�9��vHB;2�$O^b�� h��S�D��(ϾN����LT]g���d	���%�������ݵZ�8�����t���1�{*4)��R���T��¦U�uf6R�� [ɞX�u6�a��k���B�ږb>�N��,��S�M�H��5�c㌪g*����t\��d�=�ѳ������^[�ɉ��n�MqN�?��{?�v��Ȇ$Ѓ/C�埪D�n���� G"X��ֹ��m�M�$d�p�bU6�z�Z��/[���;�/�����pFv6r��~%�M1�%!RФN{N��n��� ]�,�w�F0�Ԅ������O^}�đV-�?;�<���:ךRi0�MM����
c�b�h'�p�yH��J�a����ꙛ�6����&$}�M�W��U��EO�����\�G�P��6!�i/Xf�9�(1��]*4:Hls,�_���;�_3��f�Hj� X3"l����q���wi���XiD��{�Z'M���;4v�D���͗AV�S];��md���pd�D���7��2��b^nU �����c�E�\����I�SwXO�F�Ӆ�n�50�b�h���@�Π\�T��dz���;;��w5EheĲy�¤[p��)����Ul� -�:�՘�%>=Љ\�}�����!-9~0�g*�7F�&\լZ{]P��)&�+m��9��<�d�<nz�>�W9<��l����?��#q�H�S���nt51Џ��.�M���]Z����[^����%t�33��VSZ2S����~����'�kģ� �������p�tT��r|�
����Z˫��?��0V9�
%I�r��� �3�5����`S��AȰ^|S��X��`"+_N:�a={VY�ǔ�O�tf�n���A���VL�iJtKDb���3�����sT	�©<S�{}DX��ZUY�N�����6��6Ξ-E�2�dl<�_	�).��Ll"i�-��F�P9y�m8��B=$��"t��:�9�|��o�A�K���P
X�I�0M��2����:d��!ސa�.�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��{ ��UWPCHh1D3�f��l�V����g'���P��,�!��Cy~�Ȥ�ו�%�T2�m�y�^�1P�8~u�=�Z��A�?� ���u#�_��H�! (��؝��/x�l��s��E��>$	[|��C��%��(�c�o��`IP8��$���ܒ�Y������HI�����uR��^�43�J-�ѻM9bu����"�W��#!���M^��7C�'pK����L�]Y�p�� 90sQ���E��{�]���.��"���|eJt;��c~q��x���vkJĩ�W��V:�$_�_�ழ����w)S�$��pÞ�l��)��n_M
qd����������9:�F�cn(l��a�N���F`�P��Ƨ��'���9��~+�^�~�>2�K����ƫO�'���x����� t֪��L���њ(e`$�[��r��.�� 2UmEyX����"�z���[i[��?Բn�T�������1�HM<z="�<b���o+1
�ԑv����0Ǧ�p̂��8;�X�vw�q<b�����A\yA��f��=E�sp.�U�+����� ��)s�s+�ڼ{t~�|橕.�]v�t:@2O_DI����)_�E{]90 �/�k*�KL)U��(���P��K���y�!cy@5=�����U���"�'�{&s�d/�а[����QGJ�z��ϔ�3��<�]�G�/p�M4y�����x��0	Eq�����<�FC�e���}����Ӗ�4!�C#P	��N`�x��MVZ�ڕ�^'�|�b��{���#�H��h�����S�1��/�h���5����3x��D�����A�XZ�`�k��WTJ�x�+��l���6��
��b0�7���d �ډGJ6<d� �\�F.���l��L�ŗ=��g��߹k�.�(rvBq�jg2#&]��a-I���6�x��`���]_̖qq瘶�2�CU�:�c,KߡL���er��(|���/)��X��\����K�7��܎؝Ґ�\�8%S�f���X )a}�~�9�I�)�������`V%F�M���&b�k��%n�ȏ����@+[Y���Jc���Ϧ-�&��Rt��[ Q��ѐ����9����1����0��}�f51�ĥY�vչU��T2O*PQ����봉0hfٸ�K	1�x�x���^��q]� FLx�e@T������{1k���].dK�%	�Q��w���r뾲�/��61�\?v�N#�SS��3��}�u>�.�8�	�DЙI��9Q�����т)��M�][Z-z6���&ka��=�F�R�	J�r
�SS;P���G��:�ϝ@�,,ʿ���@�4�r�B��K�[�"�#��Y�8�h�4m��늇�fEq�`Pc ٙ3�Z���⇧q?�^�/s=�N&���e�/�-�%�k=���P�s�Q�t��y&"��js8iWT���m�!Mm�s
��[���6^B�u�MaNY�mw��8�%�K����q�K��k%M�IQ��rޕQs�'�����ڥ �?d�7�G����f4X�UA&�'�e�,-s*y.�>�c��¸�K4����3t��
!]��w�90�M:;%��Fȼ��,|R-������Pa���s:�ʠ����n8��p���[�;`��-�ϔ�-���&@�ߡ���T��P@zU��j5�B	�#�_���{z��뇮30��}���`��fB�Km�� T�d����[�瘬��H���u�cp*�1�> �݈i��z*��ڜa!dA���.�#��w��$�[W�\�i�h��ֳ;����y�C쳓DW��XЏ�z8�2n�'��P9J*�E�{C.%��NÕ=N�TV��\[^�#�P'JuՄ����AA2���ˋH��u��'��>����#�b�wx��q�Ld��Jݼ��L[�^\�X�%�ґ����	��I��%��Pр�'�}�-I��l$��]��uv�^���n���_�]Σ[:U"6Zr�5Ǔ��
^���C+�p�W��C*2��MY�	�NW0'o0�hz��	�@����ƶ"ݠ�qJ�u��^��U��iՅT�J��hWM�NV^]�_d/z��x�H
wM�\$X��¿JlV�x��_�=id Y����z��D9�/�����l�����.ޓ�tx��K�
'��h9���~O���A��bIy�x�v��O�N�K��;��s� �����D����
e�.$�H����.׭ ���E�7���Q�>Z�z;��[�,��Q5S��<��D���Br4����HqX�z�ݓ�%��=<�+U���5����L4�J^�̦��?�X����.�ba��g�yebfp��E�Wz.�z��O(�Z���1sJ����+%{Ҡ|
r�.s*]���@��_h����)�I�{�N 4n%�[��o�:U��b�	�ǈU.�	V0�=ydŞ�.�M���U��S�$�'��P&���/�C�c�~�Gn�����W�;<���]G�/�V4��"��I��!�	������<�Uy�f��!^���P�2�E�g�	�|�N�i��i�rZ�@�	+�М���S{�����m��"�d�ڑw�3�?�h�5�O*�W꽑���h�DB���V����?�J�e�+�t����^�7T'��؎[N����U�JڌB�&��\XP���/äDO�Ż��M�O�j<��Џ(���q���2GH��F��I.�6CC��M�p_�Ðq�Զ�8dC�w�KVK���L���	�8�L-OE��/Mz�X.��ی{Kt�� �$�vq�\�t%�0qf���X���}2����Y�Ij)�e�,��9�%����1k���������ɝπ�˲��mOčHDc�.Ct*-��l��3�c�Qvߐ��5ٳü��]^�;�"Y��ԣ�}��f�rB��*����y?"��T0*tȰ�4���� �f}��K-�=x2�����a�Ü�հ`8�(o�`�xO܍�d<�@[��s:(���'R'��w��x����c���R�	�_�c�^4��g��P�J�s�q�@,3
��$^t���d�gnl ���W}�&�AA�7LM=t�m��X֠/�����Ե�/Q��A��%���h�%�иZ���y��`)��}����(����(mW���A������m��,�ET�"�63�(�^CM�����_^LՂ\�Tc�&���wͺv�tǩ���HN�Ϝ=�PN��\�����5�H5�3��v�"1#�`��ϙu��օZ!gq`�>�mj�
3��࿁{Y�nG�M�l16@&5�)K�u'W�-s4{G������wv̄J�c6�b>hH]1gldǐ4�1�{Ճ�g������'4�Y�.]�䞕~m�b�H��1Z"
�f��D��M�_��]r��"�\%/A�.�W�7�wѸW��g�MOhv���i���w�D��te͍7��M<���� ԁ�w(2�]M�pDD�Z��n��(o���(��dc�qD��IV0���b�s��@L�@מw��ne���9��VA��k����<��M�p�]�=�?I�q��츝h3]��/�d
��#�zl7R"�3`�g�d��{Q�H����dK�/#� �ZR��P7?d�G��묑�#ͩܥ��茤�e"�c>50H�Ry��:�+�'�Q�g�>z��(dpgSg*Y�y�����KV�1ʅ~�Szu�T��\�-�@Hh�7�E�`"fb�2S�d��(Y{����d��-��nn�Q`쬅@�B�YbQ�c#� f��_.-��%�M���(��%#!�[�$A����Ӈ�(oHk�(��c'5�>֔����Y7FҘ����8�����c:t����;�6��|n"���R)L����&������$2�|1�#77�}x&nN� SF9�e0(�{��*g�if���LM�@�S4+���򰙕����\m��8�,NZ&�ԹW��"�;T�	�궐Z@�g�?df�bo�Ny�{�"*iF�q�4�O�*T�|��5��T�ob�ty�z�_ 9��I��v
 �Z|��!m��m��t���M.�7�T�Iki���%�ߚ.H#=�$Ğ'�a�F����1��D�0���ڔ	#N�g��Tu&׸4[�I���Q>^�0��	U��6�*�!n@��mtLk_��G�z�J�������>��S�X�5���b��ƜCP;7���@�߽������h�).��[OQ5�/���yL�BI�GO���Nݾ-W�����5<
k�o�(��_���2adN�]���W�i�\��ީ��跈�1��E���ds	 2��|�AՁ ��6!�rP1/D�v'��0��I2��J9د�sV֣���^~xp(�]�>.�E��!�]��/�7G&��6��2=t"��W��	�VXrOS9S l�C����m��Y﶑`P��2@^�r?Y|�0������#��p���e�6!���s����!PH�˙�� Z#r=̧-q�?�^�Zc=��D&���J�
�����J�Mk ���s���t_D�&gGO�t8���Wy�ހ���!���s#D� ���{H��Z,�M�ݝ���a��`̥��P!�2q����NлPm�M��[����WC�%$'��<�g���?I�������Ь�4m�U�m�'��u,�'!ysH�H+��F��j&4�=٘P�����n��~���2���^�F�k��ԣR�G��`����g��5�sL�i�����趾W�v�W�`��`!�-�w��E���_� I輗�]�zZ���>QBF&O#�K<�.A�z��sk�J���֝����B�}���1Tb�7�����Ŗ�"�w��S��#a�v�K ��6i��*kĜ&C}A�.ˤ����i
W�aUi
-����;Q�a�ޭC�D��������_R�ą'�/�P�U�r#C"?��m�]����T;��f�^��P��uy���lA�8��{<�V�L���ғ��4-�N�I�g
SxI�����~ʣM�gC�[ńF�C�%��O����I�i���{����G���;�b��u>/^�'�S}������� �"�ǚ�:�ɬre^�CD�pt잏hO�bYOg�SWu0̞�����H�����9���uc���J+�,c|����+Ņ��J�PWS0VÉ�_i��wR��sw2��$ݓe���l� �k�9_�+�d�\��&����}9c����le�U��3E��ZƐ��'���9*��~t�`�=��4n��
Y�qƔ1׫0��ء4�B�+ ݄t�c}��蘚�eI�^$�s��t.�%� �\EM�#�\�z�=[rl���qB��	��	gp������,H0�z���
F/��-�+z���/'�7��O���K1<!��X�y�0ճb'�6�,T=y�6�fu6�E���.�0ۏ4�I�������s��c��{h�|��8.�U}�i @?��_���t\)�G�{� ٙ��T�>�T:�U!��.l/�iH�n�M�=�y	�n�s��Ҹ�UDJ~��?'q&���/�xP�$�g���GS������|�L<J޷]t�/
h4B�a��]��	v	nk�6�<doU����&�8�fvΖwis�L��	3N�3��.�Zp�����u�U�K�?{��*�L�L�GZ�{�s����H�h��5Эy�<<%���Љ�	;EK��	IJ�>	J�8+����!<��\��H�����u�k�)7J�G��:\ݽ[��MI�	2I� �w�RK���?���({%Oq�	2l�Q���I��@6H�&�r{���_�>�q����� �C�D*���K���L��{�N�$�1��ʉm/r��X���@��Ky�WХM����\��%|rVf�-Xir�}����լI�f���a@���T%o��V2����@������N����вڮ4����c�J�9�-=�S����
Q�����l��8$X�6e#�1���Z�پu}sn�fc���#�ٟ����߭*٫߳9M��RQf���K�Ix��D��T��c�a<��5*84Ni;Y�]r��Q��e���8�$�S�R,�ױ�=�����"э,� R��6_G��^�J&g ���6��SE,���#?�t�I���g��l�1��ΐ���AƆfq�?t��b�S�����	��d�/6D�AB�����-@ܒ5�#��i�lΥL1�b>S�1��((2Q��YԪ��0�2	Dm�U�,��k��߾6X/�(x�4M�����hE���|c���Y�캛���n�ƭnrϡj�P�l��
�Իt��\�3�ʓ��M���gUϞ�-�{(�!R^�`��ͩ��cjx�ܡ��unLF�M@�n6��!�@\����R5�{�����|B̄��\6�C&# �H�J�g�{0��1����h*��o�~2�>�]Lў����'�b�;�"ſ�Y;.�����D�M]��1"�Z/d.2�Y7��n���S���OM�#�R�a��Dgwe2�P7�^�<���E���\�w1x>�5�D	���47��-DٵN�w�`�A�V�{PVU���[��b>���E��d���x؃S�߰���{V��0L��2/�람�p}?=�S��V��q�����Fƥ)�V�����a�RX�3Es��S]�� �KȖ&�G�4� ���R(�5�dH�r�(F�Vf������8���0-��yG�:��V��RQ���>�������VgJ>y3��KB���Y�S�iTLʩ����E��*�7�X`ؙ#�1�S����vť�v:d�'�-J�n��`�X����7��QVVo�[G0���A-�����
w������e&���3�����̭P�k�:���15[nq۰�?)Y|w�m;	�[����(�7�-� �@����0�ngnH�7�^�J]&�<��J��2���(�+�"��n�OS�*��0J��"�i˗��Q{@�o�p�(��I���nցiL��푈�Z+�V����"�@��b�o!�Ze��gl_}f_!�o�sY�WA�"o�ÇV�84���Od|����o$��t�����zA ��I��
%1�|��!��3r�r�I=֒��7�AWI��j����ꓽ����#B�x$i�֦�ໄ��wp��S�0w���?�#S�����uk%�4@������>��J0E��U�Xu!/���72k抁��^��o����i�Σv��XqCXV���:�$�_���w�;BEG��D���݈ܛC)s[ih>�
�F�4r�q��)ȉ��v�@U���>.���b�9����J���g�(ԋ�`/��#>*2�#u�Pu��o����nCx9$���I�Yߗ���Y��eg	��6���$q����*npr��R6���Ӧ��e�U�*�e7�Io6XO�?�`n���B�u`�W7��~y,��}1LtX7m��*?��D��}�������� ��IzfL�:a�j��$d�&8j�9c�Q'|��,^����x�:j�>��D��E:���ы՚	��ןl� �&@�x^M�$xg��E���a�qͼFz9{� tYf%��)�7�,��7Zɝ;׳��ץd�Խ��|KY�K�X(�g}Z!�U�O�l�D�w����K��1ħ��u��+�)5T8ϮP��<B�ڴ��cY_3�F�Ŝ%�N��O�o9�]���=Ɠ�Shn��Ȥ[.
\ܬ���~�O ���?*�Eh�?�	=��[�P��������ld5��v��h3�a��*��p�BY�'��L��wI�5���.=�j	S*m�A��]|�<�3'�W��8y/s�t�#2�=i�'��M�	�a-nd�?h�n6?�.a.�%��ޮ�h���v�i�ב������.��}��x�:%f\�Q���αvT"[���-3�$���-�qqI�ø��H�"r��|�A��:ލ��b�0��c@b���*�y��
:��Ҧb��yo�)pn.�w�'��S*�@��ж�<>�e�ks��"��UH�w#��|�kfɠ� m�Q\7��#��)�M��&�����P�?Z�#Q��Ȗ(D�#���+Q��,Y@�ޗ¡Ör������9:8��W�$R+�°28�}�d�<��m]��F���8s�]L0��3`�);����[s��0��32����։T���`��ђ�{:�8Q�����C�I\쑡��08��i�ܙ1���pp}���Q�z��<�[��_�~ʁr]��8Fǥ ���=� � ��-���
[�
���?�FK@�+���X�� wi����
�A*�ɓ�~-���sQ���mrڂ�������H012�_��+?�6�����\m-�2��N? 
�>n�Gq��|��.��_��τ� ��Tq��u~,�Gf3+L2����ɏ�0��!�%��M3�T#����i��n��c��a;e�!��f}WK�m|r���3nT����n;h�Gh���.߳|�k9ɩ������<�?!�M�o�[5���B���-�N�������b*0�CY�T՚T��DU�g
Ħ�+��R��0�q�b
�Y�Mt���#�����3ݺ۰�/���(m��8�@a ���RJ8��Z��a��N��x-���YwSj���+=�O�[��ڶ�c��Gd\�OTq�G1�(���Gnifpr�	��IcT���4q��]tC�=���~wתp�=1��JQ �@a���ʍ���)A=x�2��?@*������	��U��/�Tܳ��{��$�Q�Eg�fi"n��*i΄J���qy���$��I+��޺Ε�~�to��jf�p=_6�H?�4��B3|4��(�̒��~*c��� �C��]6��6�yq��	P��1ܛ�ݥR�c�����˓�ݤj�f�Ɍ2a�<j;ץ��j}u&w�K�v���e�� ��$2n�:��D�ZM�w�n��A������e���qN^�Y�92]ȁ�K�1N�p�o�����T��G�+YvX��DĚ+4s���]3P��49�$�x]�˘i���G3��@�EK��\�3qos���مM4�Dd�3(|N@�_�e����B,r1�-��ϴ{!W��f��6�=���_(��ZxhV
��<�8�ҰJ���fK����N�^��+�����9�5_x����3	���7���a��q�ep�NP�Q�<ތ��TgГ�*�|S4�9锜Om:N\��3�`k��=�g�(�9I ,s�B' �l��&u����um�]�����`��l:�������X��:�9u�P�:��yGebxFt��O8!�$|L�wg����񎳌��\^r}/O��=Tb����S���D)��A&�\�eR�u���PLͦAL�����)�*n����G�zH����֊��\���O{�8k�緦��9��~v��q�>�UT%�E���"Sa
�x5chs�%��@��j{��K�.��M*��r������A=�I��8c�8j���S��|)��4	����x�̷�����$8	��H�/ԑ�R0R\ C����i�?�V�eE5��g�o<]�ґ&"V���c�i1�x�k\�9l��wsh����0vu�O��,x'3����k5;��Δ����|]�EH�w�3>{x�{�oP�
��fi��8!�˖PE[�
�/dO��0˧����^7�7<�n���aF,�8�MU���$��q_����d���!�,�լѿ�?���3#��-�	��뢘>n]�ˑ1J18sӕd��2Tņ�Q�kz���#y���q��׉��.��Vw�X4�e%����#ӭ���u���Le��kr���<ݪ:��<jz��(�r�P{�*~Qi�����0N�:J�՟�QL��/�sϚ�,�ʵ��/��T�%���2xj�R/a���"�*���9��&�#F"s���dO>a!MڦPN3�>l�M�i;?{}<	@5�I�ӊ A�ǲ�H�1��˵;贚��鍦��L���'V(�'HLtRm�Z��A܊9�8\��{��I���Eڋ���b�%��}hp�}�����]�)�Y�#S�o���O^�J�:4����AvRp��u��oPՊK���՛���s���m��bV�����n������6�`1'�1��X���O[�V]<1;%Qh��;�[/�m��Ql��c�(!>���(�F|}X`ԾJ�h��H��4�NB+�����
iI>�l�}#�5B��O�rNNj��Wؼ,W
q;ho�h��.��Ǆd;�󅊯yW��\�s6�)
���#�1�¼�%s]d�N7	����'�N�dA ��1ܝUve�p���֫I�LUF��}�����˜��
�e�]��[$��]�|��=K�&�4���=3
���	��cr���S-����E1�aR���d��o�0�;@+��r����=*��T�`#Kw�����&�ǿ]���]OM?PU���:�TZp��̔� q1^��=�_/&pw�W�(�a�lޗm�k�Fi�B�s�G�t,��&��\J89�RW�a!���#!?7�s<�V�ͺ!��:�gl|M����n�����=\VN
�qv(_�]�]jnM.-g�/E�U�C�Q'�/d�	���W!o?V�K�y����4
6U3f�'��,�wy��Y�U�H�*ٖ4�u��%�D�<q��;m��:C�?��W=F:���ީ�R���D$���	��7�s,=��	��P ��0��hۍY�`L�-4���G�X}�Q��試p��}z���܁XB��>#��#���zU&��`K���#��tXvBs�֧�#�T�0�_\������>����>��`��� Ʋ�i�1*U�?�)dA���..��Z����+�W�*i�핮LL;>r��k�VC��D�"��
���l��d:'K��P�u��7��CO��:5F���TH5���^4�nP��xuI��0��A�j��V祋/k������w���1����lxc��<�9����[ҵ�:F%���9���{��IWK���"Ѳ�R��\��qk�^Җ� �u��^2�b�`��ё����@�"(<�g��?�=^NjC`p![(������0�Yܡ ��T@0�AC��q����3UKƆX��x�ݒLIJJ9����j��r_��;yJZ	�W�Z�VP�_��	�D�E�N/w?�$�	�4�l,���	J_#��d�!��:z1����9{��9wlR���W��`r���5���'�2�9���~��2M�W�T��!B&�(��p�=���N�f��ȱ � ���v�"�C�g��e��1$�k��H�.IU �u�E��B��Y�j�z��[!���j�6���	�4�����H�*ze����W�o�+��&�����<�|L��9'���X��ڡ��bt���DVyW$f���EU^r.9O��A�&��r$�#!�s�k����{J��||��.%�p�{@쒣_�ċ�a��)u�3{3� �p��S9�a��U���{�f�0c�����s�y��]��"����xU�ο
�'^t�&��]/���e��@� G``�Ē^�ɿ�<7�T]#�/F�H4�`�Q�:��		��^J�<Q'�{�S��3阖�5��YO	���N�D��
nZ�!����B����`{��h���Mǔ(z�ha��i�I�ϲhT#5=�o�Iܽ�?4��������т6���l(DJD\�+�A����&��%��5h�M�ݗ:�sp��J�O�$*\��4�;SD���ŭ\I�i��u����*(�0�q�g�2�����I�h6u�G�ӻ��i_��qGZ�8 �C�-��y�SK�̠Ly����-G�>B%w��/��X�1H���VK��[�rmǝ(B{\�[Y%)�Zf0�XV�0}$�;�huIs>��3v���D%��(��|c���������^�8�G�A�kĿ1�c>�&( -ʉ�(:�L�)Q(�+�����E����������}@��f��;��Y��L�����v�*f O�fS	�<f/8�K�Jxd%d�Y�^�Ǘ	a��D�8������j"�����β���%�#���RYDα�[Gw���h����R�]_4;�^&v�g-a\���s�8�}K,e_��p #t�T]�VJgBEl��޹;J��fbAsO���7t�iV��Qa�nFΆ: /C�A�g8��=������P��6���@ӳo�3���m�c �(3������Ƞ�?�mOfl,�o�C�%6��(e�Mz��a���9ic����'ۺ�d8�[(�:���5}P�L,�U���S�z�T33�i��s�R>�����H�w!��8`	Rǩp��jhD�܎H��m��ny�YM	6��R,�����{��a������ʄ��'6f�E0��H��g�At���1�}/��Jn�Պ<_�K��]�'����r���"<ᎁ&���1���Q0]��\"3��/��.��#7��y�ɴ��şOZŐ���o�eK�DT޷e��7�4h<o*g����iI�ޜ;҂��D��������Z���מ����c7E��V�W�Hr4bˏ8�r� ��>�)�I�`*{�̜���
���Ǚ�*����pL�I=6�A�c���.��N��3���$����s���eR�4�3R*Iű뙊�ϗ������a� x�7R��Z�Br�d����Q�C{b͛@��.�-����u�0:��y��O:.K��f�Q��a>�t[��?�g8Uy²'�hK���w�QS�{XTNp]��� �Nz7�7#��`Ņ�T�^S�|]ؚw�Q�zd�B-��jn��`��%�2w��ރ�Q#�U��~�´�-/������q�����S���������Zttk�x�}i5莡����Y���z�@�P2����E����m�!��%�n��.�D���� &��7�7��2�pl�U�м�0�n ��S�Ѐ�k�����6CiXo��~�+@Y^��O0�����B�������Ge��ZXg���&#"<&^�J+��Z�6�gY3�f�rdo����$*�"�� �c�540�Ӝ�|r������oQ�t���,�| +��I�_
r�f|��h!_�|�����+���΢7�I��юI/
�>� �S#oا$6C��!?����$�U(҆0d=7��F'#��;���u؛I4M���.{&>�=�02s�U{6�A,�!�� ���k���y�F¼ϰ��06
ׅ"'X#���K��ۜu�;���2'���
��hU�)�(�hKe��h�rL����[�s��v@�U���>��ӟ�Z��r��&������������$Z>�9�#��	P" 	o����[9�9����n&�q�Cm�%��e����՘��G��*�r܉f���r�ӳeG��*7�7xy�6�|4?�?�������hWD�x+'^����La%�mm.�?4s)D�6P�5�۩9�Eږ��L��������Q���������^�8�U^>T�e]j�#s���vm���G���5�����ƭ ��<�������x4OE\n���ih���� a��%�C֒d�d�\�uZ6�;䐅̈́$c�!���|��	��x�(p�Z��տ\.�lP ���ϴ����y
n���Z��G���^8����BQ8Z����Y�H\Fӌ�%���"��oF��-���YASU�2�e [[��\���">��� m�?w�)h��;	�!�[$ҥ�sX�j-l&�D5/]�v�_�h �č0�W��Y�K3�i�r����52��{�W������y����©Mg'�_I��;s�![.=���p�wO[h�f�Ϝ����W;hvi�[�'��bA��B`Љ�>q�yÍ%�HI4��� ��1����ނ�����P���hb�=N�AЋ*���=2d���b�l�o1 nJ(�w�W��$��*�
l����<�Zd�`�e���륊�nw�o|
lIɵ=�^UQ�_���˄��m)��q������?�%Q����#,F����+&	�,Ί%ެ[�K.F�����8A���J��+�r���'�}�B�<�vh�nMFա8�S�]�#���)�����s�s�+�(�?םD־�#��jo`S"e���4��ɤ`�C�5)�&&�����!� �51�E�p%͑���z�����F����~��^]��FܗʧG�%�Up����k w
C�̓�P?���1F`w�+l�]XM��w^RРhİA_�ѓ`�2vz���~����mǯ������/��}�(2����>�O�K�ۭrSm�?�2ӌ�?�M>��$GF�����O�C�u_Ə+�c�aOT�u�GOG;�cL��ҙ����h!܉O�B"IT����u���T"�c�����L!mfrk�� qr������
����ޓ�}���cnߨ�� ����X�qA����%M������L�4ʠ�&1�-���67�dܓb?��Cԟ���Ś��w���6��?��'e�0 g�b����EtC���:�UMe��T�j-����!�@,���J-����aꌯN�Pg-B7��E�w[�03��D�j[:���`c��$dѕ����(��Gc�op�5�p�c���b�f��t��=B��~l�p���W��v�a�)ʢ�����=�s:xJ�Կp���y���~x��j��/�I��B{��$��E���>�E�i����\��Ѳ���$���~gy��}l��r~�@�ߐ����b6����O�BhJ˫�c�c�~;bcm���u����R�~��y<w����+P��C�P���+#�~���t$��Yj�8A�'�2v-y9��Թjr��wiIv�`�:�N m�+2&N̗�oND>���l�D$߭�	��x���цsPǸ�Y��ARQ�����1���E|0�Nٵ�i)GG��4Y˛��9r�+��֪T�(3%~4����l�M���b�k(�R@fw����3FZ=� �b(�D	"}R9N�k@DVe�{��1xs����{�|W؍r�ܥ��҇ޔV~�kOh˙�QJp���q��HvK�9���2E�� �w� b9��ixG��qт�Z��5#����ΆF�qe}I%Ne�����@�@~�\���85�����픜��:Nq��3��7`���2����Y$IU0� ���-���Q�$u����5��-��::����^��m����K^uAS:���G���F��O+WЙ�D�g�n��f����\�H}AcO��T���;��7s�)o ��6kU\-I.����m�����BH��X)&��n�K�� z}ǔh�K燶�G��^��ȍo��5��L�	��Y�Ո|?�UiU�����w�,V��3J5����Z�z)j��.K�Fݢ�
��T�����-,����8�8�j�����|~�s�2[�r�������ǀ���	ۚH�l��j�RQ#ZĔ�i0�V��'5*��������{����Dcg��⹑wk1�?lA2F��7�.0˗�O�e�x�>P.s`k
P��Z�ܽ�8|w�E��(��xRL��3�
��Si{uC�#K����E�
������"L������'��s��7��X�s_:�V"�,b�VM�\1�d�$�_�qtx��h[d���ź�"�,l�;������$ٝ��s������-W�@^h>c�l�&�Jf���j��ԧl膻x!k/�H�x�,��9�c�G��
@�+�lX�| %08���2�K�jo���Ӟ!�qr�wmѱ?�:'\��=ĭ-swr�5^�~�ć�&�U�:_���I
�L�y��h����{�����ƃ%��Y��G�_���a, "�	.���9)�j&�����K�}�O��av&p�ERm3V�ݲ��;�Y<~6��^}��?�[ �t���VH{y�� ;�5L�gJˍ���L�I�8��VF�H�Xm�`�bF9Xy����m��z/LJڀ,������ZJ��cp3c̢�@����}aS���+������6��A�+Yq}����@xB�j����AT�ݡ�m��lV�ٷ�O������Q�e��--���/cVr��;��h#id��ag��)Q;k���(�����Ќ����}�a
�?�^�P�h�i�B .=�n�X
~6G�!c6}x>.B�j�OO�N� 4W�:��1��
�mCoJ{��
���=�d����v W��Z\�۫�>���y}1�RY��d�H9	�Z�~�w����y���	�11��vZvBhW�=���{���~+����� 7���m�	��K0��4d`]"3�	�jB&��0��=6���Y{p	���r�?�S���Eꑪ�Ƿ��Sn�_P@��dr��#�������v#@���Y4�[�ǿ�(��M��bThP
�虏|�Zek��)Ofqf�(^�� =K�&��҇_5���ތ�k����w��s�at�0�&�^�.8�~�W�$-�a�!t��sqi�B����T��MM�\ގ�V���(�r6#�q�ڔ�(��AM���<N(x��'�4�~��l��?�5��A��P4�x�Uh�L'��,��y�Dy�
�����0�41���Zn(�`���6�� 3����	�esF/x��s��RT����7x��L�s���k���E�'�8��8T8�bRn`��0-I��Է_���,�FK��>+�z\��Q: BȪ�#�`��0�RzJ���`��T3���s���B�ġ����Td+��TlJ�.n��:�����Jc����& {&{i�*J������A��.���a|����WM\�i]֮A\�;�
���9�C��D>o��Δ�!�&���'@�P��v�l�YC$%�ȯ&֕#aT�W��}<^)��Pn�u;�����A(S�kL���6�N�M����v��W�i�x������&b�im[��.�4%�)���J��Il�7�[����7��o:�㳩��(�d+u]l ^G�D���=��WD��v�"]��<1Ԭ��b^c��CҬypvmu���7,�Y;�U��0��/Yڼ�S������{�a������J??�n���C�[��WJO�EW���V��s_k���'�3w�՞$ߺ?�)�l�v �-�7_�Xd�P�O3��	9e���*5l���Y��5�O�[����1'NGw9,��~�
�����Xg��(��B��˫��>أ����� _�K�%C��ۘ�Z7e���$�Jz�ę.>�� �\EĴﲨs�%��z��[4�w���������@v�i&���HX��zzt|��`�Ġ5+��_�|k'��7�Q��̍����^Xl6��2*�biʹԮ�yy���fw<�Eʟ�.N�N��/��;;��s����%��{P<|��.:F��j�@A��_��ֈ���)�٨{�� ����M��ݒU#�Ėp�a��,ƭ0����yK� ��a�Ô��UF'm�'�5�&��/�2�f;{�UGg��pݓ�G<�e ]6|/z�4���f�����i	pr�S��<�Xf��)�(O*����C� 2	��N��۰6Z2Eo�.䷥����8{��K�N!�ǉ���6ۑ�sJ�^�hɌH5RL �����1k�����J;���A��6�JY9�+e�L�#e��f��`���N
�E*�C{J�7�͈�\�ȅ�0����"��k�T���N�R"(=z�q�2�H����IE�6J�w�����_�5�q�_M�-��C@��®8K�t�L�is����U��:Y/�h�Xu�����K{H���ٝ=x�\WT%~\f%�X�Ͳ}Y���hI�*�,�ܓ��z%q\ �G�aS��W5��t���k��\]f�e*�K=c�\���-��(���g�_Q=��M�o�:]7�xa+�ñIY�ۨm}���f�ՁǏ��١/���+�?�a*���;洔��fD�K�"x��)�NY��\��a�18���i8v���q<�y@�S�%Χ����V���FR.ޱ^np`��U��.�R��_��}^[��g6U�1S�0����,����eB�tZ�ٕ��g�[lѹP���k+A�o��Xt,���Ѫ�/�����Λ"]/��	A�o�)]�oȒ�9L%������'mͳ$os�z��X�(��t����w�tCjmd�x,X�	��
6�� (��CMB�����E�҂#��cvQ��[�8��?P��a�ot`ϣ(EP ��#Qq�ғ��K�3(���i���Ϡw�Խ�!�:`���œ�j]i��#с���nN�M��]6��К��k��H){���Ç��~�E�1�6{����H��@gӰҐ{��1�}������՟Lr� �1]N{>��A���	��jA"�4��cH�F�*��]��"(��/��.���7�세>�*�._�O���T
��Z)(D�ze�4{7�J<�����}T�Z3�q�w��D�k��L��/w��,Ϟ�����RV���ݘb ���GϘ�'��>1I��g�!�$ϽW.��uϙ����p�O=Kn��3�s�j�����Q-��ϊ���aUjR�'�3����3��U���8ܖ�ٟ6"� ��?R��c����dJr��{�ص����B��Ǥz<��*�0��y��:�bfEQ���>��2�.�jg�<�yN��	n�K�Uʬ�oS��AT�F�r�����WA7&�`Z��W�S¿��n�f��d�^H-	Y*n�}`X0d�g�����Q���$�wh�-���}����L5(i��냺��,P��̯#6knp8VT5z��4�-AY�-�/XC�]����l�����U��B:p��V�n�\n��VB�L��&�Ƴ�Wc2�%D�*��d�nk�S�*:��E��p�q^^i��2�S2�@�ٍ�9̙Ll����$U�W4%�S�Z-��>G="QU�X\O�q^fZ��*g��Af!W�o�aU��	"�Ys���4��{ӑci|�k����o&��t�m��AS8 ���I��
gR�|a�!�?ptX>�[;��<7���I���>�Vl?��U�#DR�$����(d,�FF��y5��0�����#UV��=u�#�4vY��\^>�I20���U���'!U���4��k��5��� ±>6�E;��ex��Z��X�s���]^�Pr"���6;���FG����ߤ/�ݝ)�vh S��H�rA_�䈾�����v��U*�>��<��=ֱh�� ��{��R���@��a��>�D#7ͿPw�oǽ���9旲��1��J�X;m��z�ei���x淘�,�|�*ph��v��x��h�|e�*E*,��7g6?�������n�W��Z�0v���L���m�3.?	 D4]�*nАA�晧ڋ3�L 5�,���&ɶ�h���5�J#��^3Ұ��>�j��.��p���Y��.�_ ��x���i� X�Z�:���~x�dME4 �#�9;�O{�H �`�%��k�9���ѵ�ZK��;��������2�DY�>��M��(�y!Z�-|�?�l�G���N?ծm1������K����e8�����BFo��'�#Y!�F�[%�_7n*o�����H��յS�<ҚHE[0��\%]@-�g�� �pG?l]�h/1�	���[��=�'g�rlۖb5���v�h�:�e�r�r�Y8���~�ۣ9V5�\E�pJ����pfo�
�3<i¾9�'��;�:�{s��j�I�=+�F��M1
�a�vd�!i�pgc�p���w���a���`�5��v"ԥ�S�h��֪.���IT�:���	s�$�v���[�&B�"M�f8g�vk$q37�ú�,H��;�n���r������Y�����b����I*"
TJ�ݝ���b;]�o+Zn�_w ������*J3����<@Rۭn��jC��w%|�7�"Y0�Q�Q^�������/)Z��T������}m?TQ�N�j��#%���=+S��,�P��ۤ�X�8��,њ�8.W���B+�ʰtj}f�W<���_��F"�W8�^s]���54�)U��5�3s��2���u�R׊�s�KRg��'` _(�E�_��_O���C���Q�tВ�V��t19Pp2.͹�Iz�t��(:���w~��1]�I�FI���T��P1�\�S�X�
�>��?s��}�Fͤ~+y�KX�0�w�$��U��A�G ���TC���:@��N�mtI=������
X�2���L����ۺǧm/6�2 YK?��|>0�Gs:Ⱦ����nP_ӡV��b*�T�Bu@��Gh�Lta8�Y�
��U�!�:���T�q��R���}�0ꥮ�V9��l!�z(f�.0�-�rl���5���9���ߓ	�����T��ud�Zɩp���:ˀ��*M�N������^���-w�`��F�1x}b��C�_՜�}�:�4����^�T0��b����_jt�h|e[�B�@�|g�1�t�j�qf@#i��Ƴ�Jz����/Iaw�gN��-Jl0��wUJ��n�Α��['�a�x�c���d�%��P�	��(���G�.Zp�*ve�Cc *��/�i��Wit
=��#~���p�S
f"{�aȳ�S?��2=zƟ���quI~��m��K����p/�7�ܵX�{�C�$��E)�6k�>��
iP	*����s&ز�Q�$������T�]	M~K[�ߝ!X�ṙ6Էyö�vB�����h����k~�rcz z�"V�����k��y�Z�+6PN��tZ7�]}��TO~�˖P�a���0dj�j��Ξ32�},�9��T�j�J�w��v}��g�� :��2�ܭ���aD�qa㹃�1!��E��X���e������Y�2f��4����1}�rE�����IG���Yx3͞��k+�����j3R$�4{�����Z�	��uV�@SKh�z3s����ۅ�*D&Yz*��NN�@1�Te\
��D|m1Eْ�&(�{܉Q�<��)*n߿���!"�瘌�h�|V���Q���z��T�K���B����-����m9R�xTg��x��ؽ�"k���,*�s�5eJ&hN�C��,���C����%J>3�;�?��E@N�nt3���`m�D��ۚI���D�� �f��hG�^P�uo�ʶ@-#�pL�͈76:�NÙ+�ڎ����u��:1�G�w F6I�O:��f��Z~�g��
��%�ΉO\��}΂�O�S�T�'���B��Dh$)���ׂ\?	i)����Ç�=gV׫+)ӝ�n;�X��5z
�[�ߨ/Ͷ1���kh�:�/����rA'�����<�I�Uֳ���$��+S �5%X_�'����j�rDK�/��O�l�N���~������Kq�8��\jec'�-|+�W���_�4�:�ӷ�={��P�	~�H�t�/8R�}Fā�Ai�oV��5�@����C�(���=cXcT�*�F��k^�lh��7�\,0x~O乶x�d��k7]�'a�����|�EJ[W�u!Kx?�ڝ1,
��siH�`ҐtK��c�E]L:
	5|����a^ͽ �S� ���f7��9� �=��mr,OH�M�g	�$a��q�۹�u,k�fᦺ(k�,YG$с�����u=H�d&�׻���3>�ȡ��J�{7ӗ ��t���(k<8�%f�>�Q�Ph�Or�X�Xv�%����ߕm���N��&rʏ��~]�:�3������Or3rC��w~�釾�r�=:�u'�V�L�=���㔮?2�c����U �gqٴ�7�/�a�LB"#@����G9��7&�I�dYN���O ��a#�ʦ��3C^β�;A��<KH���Ȓ�L?� CO2	�Hh�	�S}H;ꞃ�4��(&�L��K�ٙVjs�H�W�m����C��9%��P�ޭ�����V��V�����+�p �Ƣ'���Ĵ[oS8/��}<� )��<Ŀ�ݨ�A�ꋀf�q9���c�W��Z�O�
m�4�VK������cw�9\�✩�S�Z犤�/�Vߘ!;�Mh�q��C�ٰ��Q��ݣ��(c4��#瞴��}Z����}�=xJ��ܑB-���;�}
�i�.�}%�B؂eO<�N,`�W����f�
�oW�V�*��*Ssd�޳�L8W��e\�����|膘�1��y�g �d�k	o�����ՐoC�懇��1ތ�v����`邘S����H�Q�b&���O���m����
�@���\]�'��]��t�[��?�&#���=�ת��	¢r>!ES�����Q�R�������;E�2��@m'r.�2����V?#�Ζ�l�F���'��Q��z�o�P>5�<'�Z�k �YYq��|^��=ϩ&�	��L�c����kqJ�ms�3Gtn6&V#�}8;��WI�N&C!M�s>d��I��j���)�AM�J�!N��l�����P�]q�؊���3GM0Y=1s;�;'����K[���;z?��{�_A�4��nU�aI'��,�k�yb���J�S�l�4cb��#��>�Q�}� �m����Y�RF|c��`�0R����F\[�Bώ���s�:�rR����%⽉Ń�ۏs�`�B�-��3��� �Z���0��+�f�\6z����@B5�6#�K��:�z�����Ն�����r��B�ħ�Z@T��K��q'��K3�!��ej� ��bi�"�*��֜�b�AL�.0����P�XV:WZ~�i��h��5y;�f�-��C 'D'��@�.�Hf�('�۵PmsG��=>CQt1�|[X�q�)T
����r^vj�P[0�uȘ��2�A��o��7<�Џ�� i�a}���Ow�#�����xX�Ѫ��6�<��z[T�O^%^~�;����EwI�#&�hs`ѴE�1:�}�� D�����u*�^�`C�"Էѓ�����'Z"���iш��[�^�BBC���p#\����)�$z6Y����0�3����"��]�585�ț�����ThJL���;�	��P�o�� �J�ngW�hVM�_����%i|M�wZ�$���v�l��E��i_%Zd�y����
��93�;�l��CeY��b��(1��('[EL9�g ~��惊�v#^hƃ㮫����P���ѵ4 L������$ʟ��k�e8�$��J>�.�d: 
m�EQk������J�zo��[A���q�Fg��xv����	H%��z�����R%�qԕ+	7��i>c��h��~�k�Z]�/�Xy��ߺ�b�s"ԛa�y� f�[E��&.�]яr��)��e��s~��/�{LLI|�2{.����@�+_~Y��g_)7�T{5_ ��C&w�#��U�M���d�sj��A�ϟ�yn	�bWá��U�+ a�'��&K*�/�9�34u��1GG"�%��Ѥ�ߴ<��&]�/H�4Q��������v	�"ʠ��<�vA�=�h�U�D�u�M�f����]	��HN8�W۝�Z�]���;%�Ֆ:=�{�A���1�֭����+���e%h�y�5�����O��&�_<��x?��B�8%ZᮠJ��~+r�b�З�����7���<�*�J�߯�V�\�X��}>	�x4�o ����圷���0�(Jq��A2�ʄ�z�II�-v6wı����_�}�qI�˶z/9C-E%�;�CK�̑L����=6x� [wy�(/�Xb����t�K�}Eд�흪�e\d�%+	�fr��X�pp}��v�,I��ղ��[��O�%����������C�1��c:��@���ˢ����Oc`����:-���*�J�d�Q�ΐZ���wΚ�ѥ�������R<}�g<f~�ǜ���N��-,��*(�8�h�-�a��f��RK��xf��ü�I]+adc��	G�8C��To�,�ύ ��������k���R[T��+���_��b���;BRP�_�Ċ^�/Yg/SU���L6�H�,g��˲�-tG@����gD�l�E��&���҆AuT7 @*t��K�L
�尼h�yV/�-A�N�O��41����RSWxJΔำ1P���|=���b(�D�ɨ5g�ay�A��m�h#,eW�Ej�6��(�jM�]��>�����3c�����к*�����������s�P�JL�����|e�3u��V>6�f�͟�Ԋ��!A��`ˊc�r
�j����ց/��n{��MOQ�6t����,Ω�?��ᑟ{{�W�PX̃��-����6����k$H�xg ��h�1]�m�nJ�����h���]���I�������k�">��h��X{���]���"u�d/u��.�O�7�e��.��)O(]�Rț�fHD�a+e���7Ǡ�<��4��+N8�9���'Dx�M�N��\E
�]�ȞO���%޲�:V�u�ʹ�b�ǿ�tߎ��*s�� �"s|�����
�f��3������p���=�Z��%�� q��c���x�������.e&RG1�3��ų�/�T�|0��u��c�? �RAR!���sd��J���J��] ��0�ˤGF4�5�0��_y��-:O7�O��QH��>�*ܸ����gު�y�}׾V��K�$x�9��S��T[Ja����p|�67eH�`G{�A�S����ܕG��w d�F�-�Bn^��`E9_���>����Qe�J�#���-15r�Y8���i���|�U>��e׺��]���\��k\�n%�5��
�N%Yk��<w��
�Y�I���c�|3Ӧo�����nnVk�3���
�&9�_���2V@o�Wq-�1��n���S��Y��dX�/���^x
i�a��{�@�H�_��̦�f���2=�D����ZZ�@�3�"��Qeo����Z��=g�8�f�(�o�d.�fX"^ܙ�%��42�L��jT|�췝f�oSl�t�Sl��� ��I���
�V/|N�E!!���
�(��ց��7��I�at����Yjݚ� #q��$x��֕=ԻSMT�&�j��0��*ю��#��H�ɚRuZl4:e�0��>3E?0�bSU=��C�T���v��|6���k�x?)�T@��w��FJ��'��JCa��N�
-����w�`+�+��Ο�[������ccUd�#
Rz��w�(�	G���p�!���cn��=�`�VFt��|===�~�ASp���ሽp�4a�D��y'"=ȍ�ӣ��D7ת��+!�YOʥi[/b�����{�"�$Х�E����ʈ�~�i���Qy6���۲�^]$R�4əYö.���k� ~���+A����h6��|Äu�B����&q���~U��c�l�p�Я�Wa�9{byW?��_�-P\*�B�������<���-T�/`�-éjIO���(2������mj�w�/dv�_�6 H:�2a����ID9;D��vA��uF�Ӓbd���M`��*0bW�Y�i����i��1���si�)���G$�!Y�؄��N+�G�og3��4�1������o$�]�x�� @!j��+'3��3��<��� �D���x%`N\1m@��>e�Ғ�1S[B���c{j���+N�7ߍ�Rޯv��r?h�,6��8'�"��ޱ�K�M��+�`�i�{����Km9���x� ��lC�����A�ݥ���'eX2�N�����t��;}%��͓��C̑5��񽜟�N��?39�5`�j����x�;Ip����� �Π�hҀ���u���N���>�	��?:L[�9����tu �":oG�Fı�O�|�t~(�g+�2��M�ܤu\�f }\�O<�T�t�Xv����)j��� b\���C��2�������eM)!knI,?����z�*��&}���ϛ��Ȉ���A�@�ױ$����W�SU�����5�r3���1�K�5�&?�u#��f�j�^K��ݝ���\ ȯL2��HPʷ��8��Bj3=�ϣ@�|y{����-�)��	k������V�	LX�H36��"R����O�iiK�V�:5u�;q���vB��K��c"ޓ��v�k�w
l�aÄ�*z�0��DO�rWxw�IC�k�#7�5��O>X|���E��g��cx���
��iVc�^��ݚE��!
JYT�H=��`I�a�}ҮCa7���n����b,�M��th>$o��q�7�����h�6��,'ڣ�|�e$͝���2\��e?��;��>�g��ᅵJ����5Ԃ߆�M�k�iM�s���L�O�|��\Ӧo.X���%kS�5�+�-g��ũ���Y�<�rX�ь/�:bG���,�(�rA�%�)�~�7��R��	:�ws����L�������|x&�����A��u��ق�D�ah�"1Œ�n�9D��&'\#r���qO�$�aq-;��8�3s�����;��<YҾ��ڄO �F�DH6������;8���B�ȍ�ߠL.�23?_Vx�OH�Hkm(��ڑ*93k���ÃlOK���ۓ��5��u�$�m��p ���xe�����qSF��K	����������A�n	���ɿ�&��5�%`���=�X%�mФ�Vea�&e����� W��E�*����k����V���;[k�h���Quy��E~QVZO�9f(q "��4(����}����2��AՄ�yB{��I��
���뼹Q}sh�B��9O
w:N�,�W?��� 
��]o�<��@�8��d�?��ڍwWD��\�%%�y���1���u��dM��	������՞�����/�~1,>~v�`>��Ђ&*Z2�uV�0�0o�K�J��h�����ƹ:~�����S]]��ow�卋a&-Z��2=QQm�ԡ�	аr��S}oZ�@�Ӫ`�F�э�n����M@{=r�cC׍@���xv#�a��:���v��m��(��2P�c뙊�-Z�,���;�q��^�o=�A�&��!��x^��Y���qk?w�W�s+p�t|��&$���8���W<k��!���s���=p�8>���tM�?�/�S�:6�Z1��"q�����y(��@M~�mK�	�/.'2HʨY�ڧ��?��F�ɺ��m�m4ZU�-'�,��y0N6���u�#	�z�54���utƌ)H��/Î;G���t-F�f��.^'Ro��۔,~�L���s|#V�f�࿠�m��4��S0j�ݱ�`�JJ-��Y�o)��}����[����:�z����,4B�x#N=��+^pz��t���ʆ'��S�n�xUB�0�.�(T_f�Q��H���P�ԓ�%��3>� ـi"r*����cm�A�v.~x��\�&$W�y�i.ʮ�L;�غ��NCnj�DP�Z/~ۼw<���'� :P;ZT���C�FȊwt�?��T�Kq��p^�ݕP)}uV��A�����K�^��I���o�����+@���k:xfE��Ni�'�I�dN[b\��I%�Hs�������I��?��Ԧ��W�?7SK�婮����xnu8i�^���������нJp�]�?"x������]�^���Cm�Fpq��Ӹ��
Y,�q��l�0�cA�j4�0�*��Z��"����t���J�mO�I������޸��K+J�#�WO��V�}e_�W����^J[`w�!d$�y�Ä��lX�:�HH�_sȳd�3%��֑�F|B9`+h�I�ul��_��V�����6���M'�h^9'�V~�.�Պ���q�;v���Q����؞����"� �5�@��r�r����e��$9Bo혯-.��� �i�E�}�#d� ��z=�S[�G��Ӹ��T0��Fa\��^^�WU H3]z�z��g.�!�+.8�7�[���4��h+u޾�Xon�-vbĘi�i(�y���f�>E��u.��������R��s'sL���@~{�l�|�\�.um�y�@<��_*�4��
�)Ž{��� �����S��V9US:����W[�K���y&�`�0�U�/�UA�yo�'��(&ق�/9��A���g	G��.��˓�<�S�]Q!�/���4_r����2�7M	k�ʮ�0<��t��bΣ⹭�l�4����E@	rtNF��k#ZM���3�j�Sі='{;�IŴ��B������B���h���5�����C����m�j�Fd�(J������:�J��t+ (��Ă��P��3���	����9J����hZ\��e��]��F5��:����Ũ���N(ض�q��2	��H�|I`�6���՞�O�O_2�Nq��U���C�!���5#K=`L�k����h+Ǡ^/��X0v����K�3�����x.�\��%y6�f�b(X�)`}t�]�_P�I�0��go��@��%lX�������G����K�ɀ���)`��]��cn(�v\�-H��x�6�nQxh���K��5�=��2`��d�n�V�}���f۷��**ٜ��;}���Jw*�~ֳ�{|�oOf��Ko��x��җ�����ma�-�W�8Q��i@ĺxÍN���'�u�N�0�%R���9v�c���5y�)k�R^-1_��^v�2g}ya���>�)t�,�����ti����g�t�l�cl����h�A�_���t�ͷ��X	�����F/�~�A�G�]'9j9$�;!������b������d����B(o7p�6�)@��O��m�6,�:n���6��(�d9M]X^�b�� �V�^5c>Q�Vw��8�+ǫ�iƊ6�.P�N�^���1*ƔʖQ3�D��$����@�ȃԘ(�!b``Yx���j�>�ތ؁���n�c�M]��6B�k���L5��H�{I����
΃��e��6�!<���Hߋ�g.ܼ�6�.1���j�0�JE��ȴ����]I��W�7�dV���"�i�vo�ꁄ�ˡq�]�
"�F/CO�./70�����i�O�{�O0��ըD���ed�7]<�\�fȹO�.m_��oUDF�.�g֪o6�k9z�������M��V���Tb�g��w/��&�y�+��Р�����mN��y��Lp���=�,c���>�n��*������
�%J)�<c�R�3�p��j�=�J'��ޟ��� �~�R��귒=dEA�X>���/���~Ο~�ɤU���e�V0�ҦyJW:]�H�k�Q�+�>��b�@2i�Pglniy�¾drKX���d8S�#Ti �����Pwʇq7sU`*���&S=u+��y���ݧd<f-Tnl1�`�������.�Qs&������-���g�������gaS�����T����p�̪�|kj���58��X��\��Y9%y�ʠ�X�]�WH"eʖ�
th��=��gVn$��ϔ
3�GԿ&G����)�2�.K��1��?�unP�YSaI����=�>�,��i�}R�Ω�@�@{-|��4�N�	���� �<�n��Z��}�Y�"��&�P�l�Z�g�W6f<!woo1�t�g",����T�4�H���|������o���t�ղ�|�� {Z�IС
�/�|��!��A��C�6N9�O;97-iI����D'S��p�j#�@�$����c�d�����t��x��0����5�#�O�צu(�N4����~۟>A��0�'DU�t�4�!0��o'kCr���1��a� �`΀����zcXs2ۊ��l��S���T;��i��x!đ�Z��ܸ�)0%-h��G�C�r�>Q�C����.v��U��>�:v�5�E�0�[�*�6Km!�H��<w�>���#��NPr�o"�ʘ�}�9���AvL�ݓ>�uted=˦�F;�a�Ͻ��*�Zቶ����I����e�6�*�f7�]65�6?x����A�2K�W��{��A�hL�YXm��k?��Dɬ�S�+�;\���L�(��G��ޡ�C�E��'�����p�^�ކ��(jف��A��b�Ħ�+��2#�߰I�<�� ��U.��"pwx��]Eo(��
͹���) ��%�A/������Z���;47��Ԕ��q����@��Y5h��E(�<�Z�KῬ$l��-�_��/�ɨ�9z�չ����8,L����B�R���Y<7�F#E�%��r�Bo�M��}w��0�;S�pzҵY>[���\���>���� �j�?ǖ�h��	�5[t*������Ulv(�5]�vHj�hp*���h��IY��¹�j���5��������96�Bs�Ʊ�����~'56J�5#WsV^�`O�=F�%'za��4���F�k���˗uZT��pͮ�A���v]J_���P��ǚ.C!�p6:EzÄ�����vpI[C�o�
�/��s��1�qN�p�5ֲH��v^�Ԟm��[�   �   ލp�F˸�x�rhK9�1�#l����_�)��ToڬrN�'|W�Ds��&�M3�i��P�E�d�F��FB*�@�J�O~6�I覑�	ߓc?F�KE�ַ1�v#p*�8s,Z�9lTA�'8�qEx��ϦIq4hF�w��Ձ��Ýo�,�b��<YAΓ0u��YH�T~�M�&a�l�"����|ج��)(_�f�O�jE�x�`�07M�8-��I� dh�
`�irr�����A'璩
�q��ƲLZX���h[j"�@����� f����X�'ߢ9{�h�2(k�J
>�
]�t"�*m�}j���B�I�"��+�E;�%	�B�	�LR6����4k�4T�$i��oj�C�I�n�F���F- �ѱ��:^��C�Ɉ���R��!+1Xc�6Q/�C�I�Vs��k��'M*���f��a��C䉃D~L��R�4}^�Q�D]�r��B�	��p�Q��ǘV����)zC�E�V$=y=L��dȫ^BC�	%X0�p�E�
2b����	u{�����!Ih����bEy�B���kT6pՆ]h6@��?y��&%A�X,G*�\�r�i�u�`)p!� JfJ�)Y#�M3�̘Ix(с��<!��Q�S`<4$����_�xO^3�LƷ2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  ��2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  ��i�6�|���WW&`�sK-n�h��AfىzN��Ї��j�4�rt&��,`�O��f���d-�.���Q0ϕv�Dʃ*��p���I\����҈iB�R�x�4uqNN�I�1�aD�<��2��h{�_�b�u9�1l>$F�\�L�|��� 10C`x���Ȋ�9�"�G{��	����D�ǢյO�t�t!ʌ��=	������oX!VW�=������<��)�?�M>�������`������j0����*U�<B䉵1x@YA���X#N(a��ԃ{/�C䉉"p�]6�ψ���e���0��C�I�_[.}"���̲̲�-�3t��ğ�B$�#����V��Ir��#;��N�F���^	�^T��↸6D�z�@�5���'>a~¥ܯp�xd�5k��9l	 `#3�y"����a咻   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ���q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'��   .    ލp�F˸��%�R(O5f��p"O��Q   �(bJ�q�4��y$C�c��A".
�jd�   �   ލp�F˸�x�rhK9�1�#l����_�)��ToڬrN�'|W�Ds��&�M3�i��P�E�d�F��FB*�@�J�O~6�I覑�	ߓc?F�KE�ַ1�v#p*�8s,Z�9lTA�'8�qEx��ϦIq4hF�w��Ձ��Ýo�,�b��<YAΓ0u��YH�T~�M�&a�l�"����|ج��)(_�f�O�jE�x�`�07M�8-��I� dh�
`�irr�����A'璩
�q��ƲLZX���h[j"�@����� f����X�'ߢ9{�h�2(k�J
>�
]�t"�*m�}j���B�I�"��+�E;�%	�B�	�LR6����4k�4T�$i��oj�C�I�n�F���F- �ѱ��:^��C�Ɉ���R��!+1Xc�6Q/�C�I�Vs��k��'M*���f��a��C䉃D~L��R�4}^�Q�D]�r��B�	��p�Q��ǘV����)zC�E�V$=y=L��dȫ^BC�	%X0�p�E�
2b����	u{�����!Ih����bEy�B���kT6pՆ]h6@��?y��&%A�X,G*�\�r�i�u�`)p!� JfJ�)Y#�M3�̘Ix(с��<!��Q�S`<4$����_�xO^3�LƷ2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  �xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O��   y  /  D  U  '   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=��J�E�TM�P������PŌP_`��7ju�r�d�O���<�'�?!�Ov�%ʢ���)�-#�E��-�����L9B8��	�}xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�z (PЩH��ɢ(�Zc���a&,O�$
�-ڼ1V�pU猤IV�u����B�ayR�BNj$����n ����ϻ%���OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O�����KO���O�<Fz�O�r]�pc�A�,�̨B��;W��)�1��jm4���?y���?)N>��T���GN��fg�h]$S�E�'*!���><`D��E|B|�f]�p�&��OnTh@�Ƀ ���S��;��L�Q����bi,�Oڤ��E?:���Aץ>k\�s�"O�����E�"��ƀ5h��×����'���e���M����M�@$S���ī�턙ZPyç	hBY�|�Iܟ �'����bĜ�$!DѦ@{u�@��G�Z��1DG�=�2��,�=��E|ҍ��NƤI��ןa�N��A��>(Ҹ���1(n�Q'�X� �	�i2��O�����'�@7�O�6��<��3�! �kUPub$�R�?k  ���,��䟨��\�b��&Z���T+h#�8���;n��B��@���P�h\�>ϐ	��$��>�RE�OD�G=���i'>��'Q��C�I�*�P��N�9��te�'����}����;��)��G#�e�R��-��`�)���HOJ��3g]�DF�YS��)
xѮ�3�ޏ;M�Y�'O^��'v�P����?����?ɉ��DT�p>�M��m���4	߂��'A��'�������(fZ�`�ʊ�u����ǓY\Q��rQ�:������/:j4�����	˟(�ɶW�t��ޟh��ϟ,ק� X����z5�|� , E(5۱矖n"��XSZ���d���g� ��)bH�/MªL��ЫFⴳO��2�X|R�
F�,��*##*�S�v��	$D�Bm���(w����t�@����&�'� Y[������dp�Ȕ��X�������aQ�LH<I�+�E��,����O�p����K?	�K웖fg���|��'�B�O��A�)��mIR��1�T��Ek�0�&p�ڴ�?!��?A*O�)�O��$�U\��
�F�t�q�1�W�Q\��5#װPm����'��Q�p�L�N�<M�&�J0��uv��'	��(Q׍�-~b����ҫR�4�3퉼"��h��X���Gwȕ��H�O����ɦ���xy��'�O�1`�5xq��h��Ձ����"OB��1�P�	cl����M ^V�<B+TI�	��MS����?�p������TG%R���
4.��B�$��?�M>I�S��򤙻G�4Z�'�� �ؔD�8!��ik�=�P��R�qЉ'e�!�d��U$pS'b۱'�If�w�!�X�x�-˗�V�_V$S�GE�Rѡ�D9<	ra��8=��,*�g� 5�H}`���Ȯi��>m���H� ^�4��c�0#6�d	���6�?	�°>����Z?VУ�MrcM���y"N��@5%�! �8�<��IR�yr$�@匰hGN2�~X���Q��yr� }_0:P�H�.�.0X��p<�7�	��R���q1� �F�*pd6�IK��#<ͧ�?�����kP���!�4Ӳ%s$��15!�d� ��أ9�:���`A!�D]�A��e"�-�+���C��G5d`!�	-q]��G�(�#� ��l)!��N�k�^IK#���$Y�f��(�����?U2�	�2�Н�3`e!���$}b��]�B�'Rɧ�'U�0a���@�r�I %c�Qv����d�E`Y���@��$�@L���.���H�*v�=�B�O1���M2V]�2�Uej�a�fIX��5��s���u��bt���1�]�i�=��ɽ%2���'W��eP��W�a�Z�pI�f6���IB��"|�'C�\t씙�eٖH���'�����ٚ���.�?�
�'.�TK���9���J�(L/��LY	�'p���̩A��nB�<��z�'G*�b��)��e���D�	B���q�~�'��Tc��i�#@�H��$�#��5Sd��9D�<���x��I-� s0�Ǘ(xX�2c�#�C䉗'�Nu�1��>�(����I#i�C�	���a�s@`�@�	�y�2B䉏=l��S�H,M�X5��� Q����ĐB�'J&qHt�X���b
*�ƨ��'O^9���4��d�O���h�[�D?PL$Xz2.¸2��Bڀň��K��幒�����ȓA�XSX7`d�1&�Q9p�@цȓ�8��g��*�� �Ƽ	A��ȓ,:TE�����ּ��LBR��p�OXPFz��D��$�Dq�E�A')1�@�È��	<1����ɟ�&���Z(qCD�gg͹ F0+�"Ox�[�&��Xb�uc��'5��0"O��Ѯ�4�t�hO�Np�0"O����G�N&��&*@!Y�T�"O�l!�OTe���N�i�d)w�DK�'�4���o#���v�D#)�D�86�� m��6�'�'l��Y��Ɂ�U8v� ���pf���Ш:D�p@'��(,S��s�#�z����4D�x�B�ң9M�mI'��=w_l� �1D�(xrN�T򔄁1`�*g����a1�� F�/�F�����k\r$�M4=�Q��F�;ڧ�(��"!�
m�z}������)��'r�֧� ���D�һ`JN8a'BA@"z�h0"O1
b���.3��K7@2C0|��"Ob}S���#V;�xQuOþz(�ŉ�"O84�M�!�Ti�##
V�1��'x�<�d��r\2e�1���n�Cw�O|?e�Tp���$�'�rX��:��*��˟,7��Z'�;D�di�lN�9���݉|�T!�
<D����
�Bgn.�Nb4D'D�h�ю�q9�܀0�x���g&D�,����W2�<�" Z��`"�*7}"�?�S��-$�H�Q�ݟ@��x�� �13����O*$
���OL��&�����H�F��'A�R0Y����y���1a�8���O�ay@�yReS�6��1�D.�E� �胅ܽ�y�J�%��pv��=>�R���@W:�y�^�Rĩ�b��/�r|s4�W���'�@"?"@�ß�1�)o>D�`FgK\��4�W�?qN>��S����U�3(H�ID��-p��eƚ7�!�_�yfh���6t'���d�k�!��^�2�� bSd@�x����i��	�!�ЀIЀ��!"�����$�!����h��`h�`�# $:�`TnH �d����9y��>a��㇧Y���BK#
6��u���?�����>�!��E��ى�V�2��� K�<����J�`�b�� �_�<���Ɔ!U}�X�$X&.�MG��r���YB<m��S�u:�p�㉧�(O�h�w��/�<��T�=k@-�"�O���Q�i>9�Il�'Gx���SU���#a�4R��j�'+lx��MA4.�RԐ�@H����'x.ЊvΈ��t��G�K8���'�R��I�
E�H`��Õ?C%��
�'����#�� -M8|�3�!SU�5�N�������3��� ���v�����( )���X���?aN>%?�!�C�}�� �h�3}�*��c�,D�aP��+r ���LǪh$�@�I,D��І�]�_4� B�)�v��|F�)D��0�B�z��/�aX�A�-*D�p��۴�<�Ui\�O`H���'�<��OV\6�' Ƚ��`����4#�)��a��O��O���<�`ac`Tyag��P������h�<��+�B9� �:@ht(�d�<Aң��� 〮L�v�֫D_�<1��H�t�Ќ���ސ:�<����Z(<���߂IA�|z���,u�*��K�'{��>a�X�O�I���a��a��� ~�L��@�O(��?�OH)4H�31�E
ìL�Y�m2"Or`����0^O�Q��Z�G����"O�]tcA	+ :=q�B�z4aG"O���,�h��E����.�>X�`�'�\�<��H�pO �hD�%?��Չ�A?��G�\���T�'_�X��0�׽p���j�DD9TZ92�+D�8�1�� ��A d��1�N��0G/D�@a׬A�@�eQ@|��Dg8D�lp��^_��`�u_�sT�H�k6D����٧s:(�%�O�ya���d�4}��-�S�'dX��h�^vRT" ӑD���OYS��O ��"�����1[�B����z�jL�1N��y�*PW�ƁV�"x�l��j� �y����#��q6k>:j��ֳ�y��;xI��`�#A��&�Z���'�y�+H"	�-p4�˳s�8�����'��"?���П p��^e��P��'//D)ȑ��?iM>��S���D�8�ƙ�1�!����W!�� ��)�Da㨼i�)�:���%"O�@��M&\��a�H,c�Bm;"OR�P	�<!Ш-��F�
!�p
O:�4	Q˞L��� H��mL���O�+G�Ӄ$YH��F��I���t|�=@���?��xt�	��'r <
����Q�������U9�n�qTeF�BXm�ȓ�Ρ	H�~;� ��[�PtdE�ȓu��E�F�	8 q$��s4z���	��(O��8�+�/.rP��E��y�h(�O��jt�i>��	ߟ(�'�ݰ��Z����Sc��'|\xpQ�'����׏�?.���U��3lk�i�
�'��=��O�/2&iCa�+jRT��'v�d�Iڸ
���6��f�" 	�'��а2*�T@.��L�32��PHH�����	H<��X[.ƣI* R��v��8l��K��?IK>%?��2���b�@"�Zq�����!�Q?V�*��Di5�=���5<R!���8�q���Al!�h�+�
.8!���G�@�SÐ�#X4�7�!�Dݐ9=�Yw
ܡCZl�ْZ��qO<�F~b�Y��?I��ς`�#�
��b]5�_�d��|"����	�7jެ�1*��`����m� e��C�W8��䅞3���؃+[/��C�I0����č�'`���G�;m�bC�I9���S�U"hohY�Ձ�W�B�I�5q
�����f�\R��(T6a@����a�@�}��[�c�"��D;4��B�i�~�2�'a}�AR�*_�D�R��D���B4���y�G���)�O}��w�O��yB)�97%L�2
��E�%r����yr�N�>�t�s�F7;x��Uϒ�p<)��	=܌�A��M�F�z8�s %@2��Z��#<�'�?����$^4V	�eJ��DU#�H����F�!�dȻd�TM0���8V�:�0T!�D�G2l�`#��'F��1G�iO!��.P�0(��0@����s@!�	����	Nx�Ɛ���R*�E���?���$¶"�& Xׂ��6d�`*"}BA�L'r�'$ɧ�'^-��j&*
�|�h� LWEy��ȓODP(��ݢ%���l�,���7��yIg�H�"��S ��4Wu,�ȓC���8��[�(�# .\�ȓ<*��%���;T ��r�֓.:���=A��I1W��DK$S�hq����7Fx�{��0ZӴ��	S���"|�'ɸ�`��:a4�X���C
�A��'0dl �!ZB;>���*�`y�
�'� PåG����
oE<�	�'6�5{Qo�!#T%	�L�/1�,��'d���"�`��5�Ć䳢�~�'�����i��y^$������K�P�GA[E�L�	៸��I�\�2���I�$�u�%�T�#*VC�;?*��{C�[u��cj�L�C�	�o7�=af׾c�H��b �/ �C�I"�r$d�#^� � ��ś<����$No�'t&L����O� А�`Ќ{���+�'{B�ي�4�"�d�O��#�����5!e�|$)��bЂ9��Gd�����El�� F'�)^	�@��-l�e�1�8ErL�e�-����
�� ģ͔a�(�=_��ȓe"%(À��uI���A�&Ѐ̤Ol�Dz�����9����1��~�D�v����R����şp'���
HR���l�tl����r4�tB�"O���%�V<"\Y� ��B����"O� 0��&F����a/�5|$t�"O�Uqcg	/S��qU�[�hnD��"O\0+S/�&(�q�o�M^H����PY�'��ɋ�7m.ly�l��j��]��$Qc�ds��'��'��Y�t�W���q����!�zԩWb<D�Ԙ�mB�nҔ�.�EnJ��7%:D��� 
��C&��S�U�F�R�3D����Ҿeꄡ����2�4�iS� 7����<WԨe�?X�Q����'�'G�Rٶ��3�������yub�qT�'�"�'oƔ��ط/ �0�s��*� ��'�n��pG�4�"���0u�(���'B�,ȵO�sG���$C��s�<E��'�αK"�JY�Ҩ��K)r���(ǓT�Q�,�ӬW;M\k� ӯi��f��@�'gE���d�O��2�2W�@��� LN�g h �O&W�Ȥ���OD����Z�g≥U�N�)���72z5e�N�yGF�"��P
P���	P�'4�ф�)�3��^��+E擹f�n,["5*�p��I|~�$(�?�'�HO �� ٨V.H�7DE=\�h�U"Oޱ�C�G�ZU£��f�� ���>Qs�i>U�	d}���2n��+�k���K7	^4j��ᢟ�8�	�P&��O%f�!v�6��Ҏ��l���+��V� �rk
�p���'��T{�
��?f�%R��[1A}��y�
[(c���  Y�G{f�b��'����D�l*�	Jce�#�b��aD��?Q��hO�b�x�C��Z����G�)��c�"D��Цo�$# �ɗ$B�e��!`�"�	��M+���d16�lx�O웦��h�����_
	�H�C�铧 �����<����?1�O�~��d�ϣm��US��� 4x4Q��O
v�ؤ���jW̉c�=,O�� C<�b��A� ���9���4��r&�hWo蒥a),O��� �'��\�(�e�X��Yh��H�R�%��H؞��-]���)sCG^t��� $��;���A�����������䌛nnu��Xy�T�X��i�'�?�J~b�4S��<�5͐6
��aJ�X.�0�'���+ �J���w�p���-�O��K�Te�[�Q�d�ѷX�B��U�3�ēGނ!`�Tt:X�!Dƨ�(�:�(�R!7O�8�TꐺD|l�;$�xB��!�?)���h�X6m�-G$��.�g��8���QC!�d�vNr�� �ʏF"Ĺ�7Ŗ'�xR�<ʓSi^��R��5|���QV�R.!��}���u����Ob��S���D�'�R�'��I���%Q�L�Ę������B(��&�H�!��L�g�I�O�R1ۄc�W��X�v㖲y��$��.Q }Vt�3�|i���xr��o�t��O�#.�(hEn��N�\�$/?i����SS�'y\m� `:}���dށU�ؤ��'v��R��/KP�T���;a��XQM�,R��4�L��>��%S ~��:��Պ&S���gh
'{� ��n�:���Od�ĵ<a��?��OP�x�Gl
Wv"�S�lM�!(Ta҂뛚M�
 !�w�`k��'�԰q!�
?7���5CӊoJQId��#�vp��mR�	���'�pؘ�A�f�� V��<r�2
���?����hO�c�8"L�W�đ���[�>�*�p�?D�XY`��&��X��{�V��qO
@nşL�'�l�C �~��4-Xᑀ��=�z��N�/)V@�"�'��	��(���|rq�A0)� Ib��Ú"��$��B�ʃ�T4�^�q@���way��4\[�=Ѐ�V�GE,��3c}Q����+�,���ܑ	���$]�5q��'!�	�m@�d��l�*e� ��¤Zs�t�p��I�]���#h�3V2ൂF3�HC�	��Zܺ�I<G�ԅ���3���V���ܖ'����[ir�����M��@-.�舘�D���)@G\�z�b�'���)�j�/u}*���4�r�-�@����C_�Z�$����˥O�r�!��
戟��z�k޷i��ӱ����TŞx����?9��h�x7-Qd����Ÿ]��%�1�с3G!�dC(��XC��
1�b8	Ta�+D�x��6ʓp�Nl�_*bn�C	I6:�!��?A	�&�$�  @�?�Lɰܪ���,�yRM�P��*�ꉅtİe3�b�*�yrF۲���(bJ�q�4��y$C�c��A".
�jdԂ������VG��(���:D퉲? |��ń�72f�1WV�|��֟H�I]�)�S� �Q�	Z����җグ �B�?e�P#яG�-��)�`��M�B䉬D3ĥp6��30*��9&葭��B��-P���KG��"ОѺ�+N�32�B䉆a~�AX4�T�H
s%�E���OV��>�� ^�Tl��'fR���[�~��S�C��l�8�ʹ]%[�����ͧ<C$����Ie�LK�Y���HH�[��¢;xH��I4=\X��0�	�Q���P Թt
�qq���!U����Dֆ��'���'\F��Ua��^LAPT'g:� �\���I|�S�O�p⢚�/5`�I��B��x��.�"�]�r�6�x&CK22F�q����3�?	,O.T����O�?�����˧l]
�$�d��P���lVޟ��I� =���3I+�)�'<�0�A.ǌ7|�|���Z�p����'-ܠ1��i�S�Oņ�u��
�.�q2��!.Py�OTU���'pr����� ��ݐ�%+Ntt����.[��'D"�'ݾX�AnŔe̐hq�(�m��$�F�O�8C��M��xQ,0}��Ի�{���ʌ��O���'���/
n��6��?!�>�Ӓ�ѻϸC�I�s�4�c"S-LzE�47��C�	�@�0��hS"�ᯚ�K3PB�I�7�
�� �&o�D҂ϓ�l�B�ɲ3Ӏl�P×	!Q�D���R���˓ ّ�"|�s�l�Ԅ��&T:a�#b��l���?y���?H>��Vi�����<������b��z�	�f�!�ݔ&��!���A+^���k��\�,���9�O�%��H�,N�`C�g�iK�U��mz��'l��'��)�<�,�<[,����`�"I����yb���+Q�	�a%��tV*5�6�X ����&�'m�	�1��	v���A
�Y��EL�ߎ-��$��?�L>����Ԥ���O� ~�{"Y�@o�IB��'$\)���'�4�[����O(�,8C#�<er�ѣ%F
2ax���?)��|�"��X��X����y�$�&��;�y�J�s�^���L�r���g�4��?���'����a!%0T���6��O��L>qAN���'���'<� �lQ�r9RU��K�7�xE�5�'��B_*̜a���o�8��\N	�鹢�O��S�M�䈙�	�<i��[�]�B�;n�s5H*&��pЯ���Π3���z�'�}J��Ѝbrp�(Â˧<�&�'�����~{�V�'�2��4�'�\��bH�}���Kr!�S��L��'���'��'���bF���g!�%7��Ę��d�g�O�TaBD�	A>�z�E�70w�(xf�iMP��b2!d����<�	k~�"I&H �� �ƅ+� ���XCvD�O���b��	:�1�1O���/�_�V1y�mO?=�f�z����	�J0a�)�3�e�` ��
-(�H%(�H��{,�D�O��Db�d��4�<���p��ױ����E�
?�ܐ��'#ҩ+���k�Z���a��-��`�,OP�EzR�O^�U�pI1O�/:�Ęi��`��}�t���\���4�?���?Y+O���O��Dϛz��U34 �*z+0�����38�x�	ċ@(SP˅��p>���;{�<��$��ޠ;�N�d:���Y�y�Ђ��	&g� E�&�A��uHu��EeRP���PG�)��������	��M�����O�㟜�)�e���j�^s,ѣ�Wx�<�6L�'����M �ޕ"�oJsyr�'�r6������'��)��>��D x�卢m�Ҵ[ei+� ��������Ov���O88P.շ$��勅��<PǕ�4`%h�"�N���i�z�`��mO:��{�뜼~�2y"�͖;�ԕ�k.u��HVZ}��,�e�'�&���?�Եi��i�OR�q���WT��$�7bn�	ٟ��?E�l̘<�z�H��H"9'�� ��M����?x��$���>z�Ƒ�q��N��|R�'�x����U�� M�hX�4
��lN���b�O��'�O$�p��o�0�F�L&~��Q�"O�1FA������d-;�|"O�0@��/Mx���,W�6>̼"O�љ��3p8��b��4�e*�����h�U��#1(<��ƭȺYY��'/���4�R�d�O��8�e��D�:hD�z���t@����<p�&��c��jѫ%]D���z!�a��+����}���!y$��ȓS�RI˲oD
%����C�!G��ȓ7�I��� �'�bt���U*+�≖'�`#=E��B��*^��8wF����Q3�+���g~,�D�O�Oq�<�B���.��Ze��2ffԅ@�"OH9�W�;�h�����*T�Mj"O���tnX��ҍ'=FVܻ�"O�=�wC��M�Y�D܌}&��k�"Otx ��MT��&�՟uxh� �|�K*�E�J���=��`#yZEs����0fj,��W��֟���O�����>Jh�Z$Ky�uc"O�]T�_�T�b8�Ã�{��!Zr"O�h*�e�!"F�T�Q�dw�4�u"O�LgIB�wa�Q���-][�L��'� �$��+Q�%�2(K~M@!�=Uuў(rP5�'(P�\ۧd�:[#�c��Z�S���A���?1�pj �ST�m�fp��h�!K$樄ȓ"k4ɐ���&6rx�@��H!���ȓA�vݪ��Y�4�H`�S�Vf�m�ȓ/֬�텶,�.xР(*�PD�/4�'q�J�k2�e��B��r%�O��+B�i>%�Iޟ0�'Y��{��w�B�PCh� BhD(0�'��ase�&H�>)᢯GK28S�'�~x�3�
C<d�7�T-� �p
�'����nȁ^t��F���J��	�'��s�43'
IR���iV�*O2aGz��	�{��d�ͺ|u���M
z;�I�I��Iԟ�$��>5D��S�^��D� 7�8,�T�$D�� $��l�8�0���^�ur�"Oxh �
fڅ�.O dct�i�"O$�@Ch�%\�H���MD,jP���t"O��`�/D��u8veX"/dd��|��'�h�L���g^��s'�*,HNZR��^����~�Iğ���O�PyfCKB�h@�3l�%����"O��Z���HR��,|g���"O��	w�N�I� A���įwg�0 �"Ot,�
-s����Շ�jTHH"��'���Dφt�������uTX�J��L�A�ўD)D�"�'r��RJV���ɀ̓3�@DR��?��C؂P!e�B�xl������.׈8�ȓ2"����͐"?�R�x�����ȓ�T� B� �x���e�#b|�Q�ȓ|�i0t��__�����ʥ{���ER./ڧ`/nM@ ��9�9(@
�Jo�8�	�{=�"<�'�?q���Y)i��r�V�0��2צ͏y.!�{�>��(�!�80!6&O85-!���h4����[�]�\<��.�)'!�L�C�H�B�K
,�t�b�O��n!�d�8�@y1�Z�<�6�`��Xs.�	�HOQ>�j���Q��`s�(^	Kԭ���<�t"�?Q���S�'"��Պ��H85�@����`ppC�)��	��b��>��`[�*[:��B�I�F+^Q�5b�n^��z�����
C䉒4�k����jf�,h�ņ�C� ?�5�p�4�dE���7�1O��F~"ĵ�~�D��D�(M�e�ý$�sc%�?�L>y�����IJ���B��5l1�G/K�B)�B�Ɉq��g酌U�}!��^G�B�IV�����-�����	�A�~B�	�<�Z�#��͟LF
��t��o� ����ş�Iu!ȃ#ü��D� *V�2V�1ړ9���G�$ڥ2{&)����k���b� �6k���'Na~r.ȧIc Y���A5�a��&���yr*Z�����:Ѱ�X$*�yR�S�hi#��o)`�k "e�ڼ�ȓ*��`
2���[��`��Z !OJ�Fr�7ڧw6\z�n_���0�Ȁ 5�r��	("<�'�?1�����$K�h�T�ʒ:��&iM'7!�ġq��!��?���mՌ:!�$G�p�f `� �� �+v0e�!���U�P�ր� Z��A���4nN!�Dˁo�p]�c���nt�(�W	ύP�I��HOQ>�i��<b�e+ro�k?��b�<a`B�?�����Sܧ\�e�F�J�\��E 2'�����ȓu�Z���M�Q,����!��J2V����<���B�>ĸi{� �U��m�ȓq�j�`��?)������*G�Ԇ�7/R�1���-<E�D
SzA%�����Z?VB��݋wߢ�������iu��~��|b�'���O.8 ��Ä<���+ba=zN�@�ȓ��Z%��$=���-������m>��y�"
�+�.�괢�5h/�ȓ`�j�i��� ��阮@��]��	*�?����1m�}ؗ$ ��T�0��J�'Վ[��ɘeۺl�c�̃0��(y�f\�@N$���O�����'����H7[��#�mER!�S݆x��܅Sy�m+�I�j�!�3���26OS(��H�!/�!�D��Jm�a�U�D�c+�4
�џ$Њ�I�[���iD�P,4�Z-��J�_�"�&�O��O��d7?q��Wq���&dM(O�m�F�Cl�<�.
5]^�	cѪݬq6���a�<� D�r �M �)H�i'Rv6��S"OT-I����y���ϢM[P�P�"OJ0q��	&n֥k䍁�5KH��Z�������G�$s!�Q(@k��W�K=:˓9^�P
��?iL>�}C�N9Q� �,�ڜ2CkP ~�j=���� �oª��H�F�l:�t��\Ҝm�"[�"�|�pWL=+�Y�ȓ=��XJ_�P�BE	�7bzpPQ� =D��Mc)�p� �dd��荹G��'�#?�)\?�ņ�3vuBo��B�t���x'����w�g���/���&!�ҀTb0C/�!���_�p�x5$�DD\���%3�!��=�đTg�h��D��+|�!�M�K���0U+��#�����`�8\����OZ�7C������W�M�A�8��v�	iz"~�Q��V(�4C��g�FH�+��?i��0?�e`��- �����E�L\jؑҢWc�<��B�2Uۥ��0SF X���]�<�T,ۻ~�.�R�Q1h2���\�<�`dA$g^�R���*.��("�X�'nb�}�D&^t��ץ�RZfx�Țٟ�7��|��?��O:M�����NQ����"\�4"O�0Z*�Wc�8xsK"O���#�"O��R�V-D~�tf昰p��R�"O�uJg�^�qo��٥nQ�X���"O���O?1����F��\x�R��+����/a>���c�CN�֨(5��4@�p��4Q���?�I>�}��`Vd1�@�6���'�x�<)b�
 8�x�r��v,R#LN�<��%A-.�l!�ܰo1h9	��_�<YfԢ`�lE��n�#x@�X�k�S�<�0��j]�d� G���4��1C�M�I��Oc��O��	�	�^ʈ�F$�j}�{$�'��'|"��>I�`^1<R>����P$�l�"�K�<�-<y�����BI�l���C�<yE�D��]
�E�$-e���U�<1�׮VM���h� ,�05qգM��,��<��DPdiʐc�p8��@2r@�E{b�� ƈ� ���C˼KKP�!(��W�N �r��Ot�'�OL�H7��I��	!j"��"O�m��Gt�`H��FN�k;��*�"OJ���6
U��dR�O�N�W"OD`ڢ��Ʈ�!$$S+g�[�I��h�<ԀeL�j0X���Bړ(^ْ�'�8�S��4�b�$�O��7hdAL�6A�����:�b���)6�Ke��Z�� 
�"SZ�ȓ��%��o,�V<Z�F2)�j��R��U�3�ʁg��ةL�Z�6a��Yʺ��p�Y��ԙ%ǄJ����'��#=E�D�!R�i"0�ޯ]�����T���d�@t���OƓOq�6X��"��AifHN%Ѧ!��"O��7l��p&��[`�AS�"O:�s�'�ly�@�����*C�sP"O*x3�˴'3n�R�j�w�f\ d"O�öd�xs��q$H%O(q�|��7�k��0�-�ĩC� �U�h�Y���=8�h��~������O�X�a��|>�Bf�)qX�S�"O� 0vP>Px��C��:M�$,�P"O>�##L�!�����Q�_���"O�����\�HcL|D�	1&��r��'�n�$��:h�5�7#��3d�Awo�3�ўh�TD1�4&�!�)K�9D�q�R<������?�i�&�0�@@�6z~�8E&�
���-���O~ ��@� TG�Ti��S�? "�٤,V{ �)vG$����"O~�{2i�-!�
�ħH��ta���	�h�̸
�e
R�B�1Х�0Ē���'�x\ۊ�4�����O��G���yg�L�Y��ʒ�)j7f-�ȓ_w}���'�I"�$��8�H��bO08�p�\�q_4�6+Bs�^�ȓa� �r�k�nl��I�mw~���E�y0�m�.WY�]zs��?����'D�"=E��-�':���1D�?I'���RK]�����v&�$�O�Oq�����- g�\F��t4@-�2"OLRsG��hP@Pl����q�2"O�EY���2�ƌ�MC�ei:$	3"O"�*Ղ�zLtseKN�b6�y�1"O�� ��+�l P�d�x���R�|2�2�=���:h���/\�yЪ�H�[�ԝ�	X�	ݟ��O s��|`aXCލ/5:9"Oj�y֠��%��l��"7X��I�&"O:,p�-_'=�.mxB�AH0�!�U"Ot8uj�8q�V�9��:?�]�V�'*��$K�;r!�4�֓.��1@��r�ўh1�=�'|�І�A�f&��U�lU
��?��z�>�RD�38v�x�U!�4܇�~_��e�a�Ѹ��q��هȓO����Ƈ�}S�X�(ԇE���ȓ(A|����j;ll E�ą[���G
-ڧm��u*P�U+����M?Bg����/X�"<�'�?q����� `� $M��0��,����e0!�DJ<h����cC�w��ȑLl�!�<��mJF��2G���(M�!���bni۱�A4-`�у#�@!�D�?�d�;Cf��x��� ���D��&�HO>���&��]Z�,S3�ML<�r�f�0*�%S�y�n�,R|��	
|�����'��F	�,9�bpn@ �J����;I>)���?����wG�QxD�`�\�+q�����F���`�ƋK=}�r���/E��O�`�c%�������W502˧)ZвC�g,Գ��˫x�(G|�AE�?����ODlQC$��O��!w�UiN�.O0��D_:M
\x%J�(?̕uh��t��}���<y��Z�G��B3#�1�:P����Wy�ڬ�yR�'G����OjeY���[�l�Fe���]X�-�O���&_tX��/��s���)�'Qj\Q(W�Hj5����^�mht9͓Z�f�ٵe�
yx��E`����%�\�
8˗%e��,a�gP��yNC�?���������d�4@��oe�X��M֣`tP4:C�#D��:uNϞ�f�&r,(���;ړR�?�q$
ܿ-�t�h��$
k���K��D�Iܟ�d��?�M;���?������O�����j���p���JN:�8��U�L#�q�I�P뜜��F����g�'�I�C�-CBm�"*�F���h��׮�2���.�ת���ɫRP2�Ɓ<�pس"�"$�<�>{*a�I���F{�:O�(�EGU�s?���ʅ/��i8"O��v�؟Q�j�����?��)8��'Xp"=ͧ�?y/O.�:5��'@�!������ b��rr�xn�� �	ԟ��'��'0�ɋ"⹫΍4Bi~I��)�-t!`a���;3��c����L��� 	��pb7f]>�Ak㤜:2@��D�b�š��/ ��D�b����d.ڸ#d��DI�I
������	G�'�d���D�!*D}� !^�_#����'�lb J� K`y3��R�L��,O��n����'h������~������F6#����'���71�m�vnZ���d�O����O�����&�c1�×��4�܉8���8���QƬы�r�a�&s.J �ج+�Z�sJ|
ӧ��d8 �Qȓ�,-�8Fc�s�'f�4i��?A��Dhݔa���"�^�C��%�"��(��*�O�m�c�(H��䒢 !i<H4c��'ö˓Hm����O�8ZE5	��	~��'Z���h����O蒟<�$�O��â Y*:��K6��R���	]���[���:5'�8u���6o��'��OZ��ks��"yVb���i��GH��'���۔�K�<�VYcc�V=�?�0�O[��!R%̩u�!�F�s����/�O���;?%?�秀 � ���H�c�������
�(Q"O������$e{2�B�x��08B�ɮ�ȟ�hhr�Ϥ{"�`Ɂb�c�]3� �O��$�O�aC!������ݟ���^y��'f`Őr��&#ހ�� ����u�T}i�
2L� �c�<���I�q���@�e�&��=Ӊ��>�@��O�-��^ÐtA�?#<qF��&�R�P2/�Q�^���o~�^��?I��hO��(�FU����1;"����Իb��B�I2.������u�Bt��FQb�h��Oc�����'g�I�p*�Z�
���I9ǯϔqBx則�U�M[���?9����D�O���`>�:��Ha �4��,ߵ��U�W�/�Ԃ�?�0�
ۓr��!�Խ
;ޜ(��GZ�8��%$�,��К�A��eia{����?�S�¨#�Ұ�#F�dlh�Sg�4�?����.�8��C�J�F$�*@.Z<e ,��L�1�gB�2�M�"��EQ^����iR\�@8�'}��R��"�����c~�!�d�˃�H� �Q����?���^KŪ�`�r�Z��O�C��YrQ�՜Q0�qÀ'��6��8	1G*[}$p�i�.�<P���ʉs¶��6g�?Vb�����O���O���l>��/�c���d�;n<j�S���O��$9�)� r��\�9���薁* � 
�i��	�@=����E��L�F��'��S�X��?����?iI~����D?Y��L{�υ6}\�qϖ�Tax��'|�Ov=!��Z����dL5k���P��|��O6�{��d���b�`^�0�$u���I�����\?���`�T>�I�,�E��L���ƉwZ~�IDJNK~�!}Rb���I;�ħI�.<�hT _��H���d�\=�=}�̭�G��'@�-���O�]i�u� N�>�TM���ܲ��I��	<���'���.�Ը���Z ��gU9��<��a�'=hy���M�u��e���M�M������^����_�*��FP�5�6��O�lڕV�h؄���I��<�rF]��v�o&��O��G�T�G?��l���"�A�eh�W���	���ҧ�9O~X����0���C �D�"#��}/�,��&	2X�'@콠�Ox):��Ҩ����d��n4.�
@$��^"�J?��!�@~ʟ�d�#-�����N��C#�&6�1�
�bD��Q؟��Q�W&I�$�4j�"k� ���'D�L�ED4I� MX#,V4��q���dӂ�D0��I��O��禵��m�m�5��8���*Gp���$ ��`��y��M�ë	�>@��B�˅#(Hs7c�^��W���OZN�ч%�!>">x�(Oa)�р�'�v(� ,΍=�|����N<W�,0�
�'cjU�Q{��q�K�H#�'[�eC��ţ,�<JUܡKHx 
�'���as�)l(�ZQ7R�	�'�N�8R��q�TXqI0��	�'�<��g�-��mk �͢F����'z(�����~И{RK�D���S�'�����#��&��G�;C��,��'Q�D��-_�8��3�B�5)U4�X���ON�D�O���O.́�̋C�8(�t̞-@��p�U��柜�Iɟ��	ҟ�������͟H�SB�� �(��B�O6G�<Q���M���?���?����?����?���?!@�2��+S�Q~kȨ�A
%M����'`��'D�'s��'���'�Bg0
ݎ��ʈ�s<�`1%�
6K 6��OX�d�ON��OV�d�O����Oj��Ց;�l��R�j�<BG�I3YqqlZϟ4�	؟ �I矀�������ԟ`�ɉ���MK�\�td�C��\%:���4�?���?q��?����?���?	�i�t�"�"Z�X�Bp8Äѡ���f�i�B�'`��'�"�'���'r�'�^�(�lC�Hj��#*�K&h=�W�oӂ���OJ�d�O<���Od��O��d�Ovl0P��P�d+C��`D ����玲�IП|���d��؟X����p�	ן���I�:}mp�ѳ����كa��M���?���?����?��?����?Ѧ�ζQmdM��I�	.���Z&՛��'Z��'_r�'�R�'FB�'R"��	Q�b�(�lK#|h*��2�M%Et�7��O����O����O����O$���O��^m��t� YYt�#@ $Z�=oZP~��'M�h�O�d�����r"���6A��6lcZ���'��i�Ħ9�_�fd"�$G�?��ݛDټ{�F��I�� Γ��$�)�(��7m��8��c� m�	۵0wi�t/�O���?s�1��|B�'>yR�G��IXѣQ�rZ�ā����D%�$M`�'�?a
� ,��-!8��Zq��[��p����B}��'x"6O��/5+hEb��#q|,Ԛ�G>r�T��?��(�'���������ӱ2O�j�ϭB�s�Y�"M&�H"R���'L2���I̎'��D��ԋ]xN�bK�O�,�'��	��M�"�O@`�Y��Ok3��yBM�"{Դ@d�'I2�'4r�Z�|������̧4,�Ķ�(}����r��؛�LͽC\6}���	ߟ��'�1��(KE�~��8�,0✕��U��O���?	��$�C}�Z�T_6���T/V8ꓪ?���y��i�+ٚ��i��Z͖�@���%M�&�`��'�j��Ăǔ|"Z�41�Q%:�P�FI�"l�f����R���B�O��	���`c��N�}JqPC�W,6�`�$�����?9�]�t�	��0�.X�(���E��`���#.:]9ҤAĦ���?���!N_����3�������.;R���P�G<U��
��ߞN��d�O��D�Oz���O6��,�'t~8��πT�\�����R���O�D�O�'�B�'UV7�,�ɘ_� ���W-wҒ����Dy��O����O��$αwH6M.?��h�> �e�ʠc�(��	�V�4Ic!CD �~ґ|rR�pDx¨���
P�썊��1g���'����?A��?!ϟvH�h��W�r��PD,�t� �\�ڭO��d�O�O�'V�VS�H��*�\�Q+��t-ʱbkũK��]mZ������VY��'V�'�*�B:À	KaE݉������'�J�ă49Y�<�����2��'���U���ܴ��'�2�:��-Q�t��R$d[�l��	���\;M�7������]���'��P���?��?E!��4�����w���� J�Oʓ�?)��?���?i�����PfzA�٣u,Y�E�^�^�8��?����?IO~�Q���>O����C�K VP�@���q�N|�D�'M2�|B���
��N{�v�O�	�HR�H�x�*�]c`��B�'�$=`�K?QK>�,O����O��8Q�Y$k���1����0�Hĺ���O���O��į<aZ��Iߟ��	#q��9�!��Ja&�pb�\�y�@a�?y_���ԟ�$�!���=1�f�Q��k:ڴ!�ddy�F��7��@�Q�i�0�����'���^,_��YY0�Z�N� X��'��'���S�<��ec�A�e���
����A�̟İ�OH�4��f���l J�̌���fs�B�I�����̦��۴L��H�'؛���t2W�V���ߋe_��Nݼ|�vq� �X�&�֠&�d�'���'��'|�'�D�&��{�lu��J00*� �Y�2�Oh��O��$5�i�OHM�Nu@�KT@ԥ��ʓ�OD}�'��|��4��+O,	0��8uT� P)_5A�MB��i���I�v	r(��H'���'��H��N-m�"�����2tk4�'�R�'���'U�Z��®O��d�LJ�	��kT����)�L�/�b�ভ�?q&X�H�����Γ>��<���
P�k� �$@��u��&ŦU�'� YK'�O~�O���(d��4C��X�`�0���^�x�2�'��'���'���n��Y�`L4F�4�� E�X�����Or�dWW}"^>���4ܘ')��'E��&
�L�'�.N�K>����?Q�J�05�ڴ�y2�'jR��1o߮����z��I���".Z�������4����O���Q!~��R�JU�S��<�D�t�s�'P�X�2�O����O���4Ҡ�Q�X�>q�.�Zr(}�B�ny��<����M+�|ʟ|-�E
D�Xl��iQ,��[�hT��W]D�4!�I�����Q�5���O��C��X��go�S�%�¹��'���'�B�'��O�剭�?�0�O>�xQW@P�}�S�Ժ�?����?�7�iw�OH��'�E��8�������ʚa���p�'|��C:?l�6���:��'��ɛ0[����N�T��X�vH����P���	�`��Ɵ��	��X�O�P��N���x!��M
o���Z������H�	_�s� 
�4�y+�J����Y]n`3&AX�/��i�&�O�OD�]���i��$�.��U�Ů�7j���
�.M�)"hܓ]�`�	�@��'��������4(PV\R�Y*��psf���D:�,�Iџ���󟤔'g���?y���?y"ĒȽR�K,e"<9B�����'~��
���wӐ�$�Ѐ�M-"zʬZ0eH�l��ǃ���ɻɆ(
��o||і'��tI�՟���;Oح�֋�4s�,�[�ƭLbz$��'��'q�S�<)P�I<��8��#)��9�G$I��l��O˓Y�6�����ͻ�o
:��8�����S�R�
0��O��oZ��M{�ixj�`G�i_��=�݀e�OR�e{wa�^��M�e��@����@�IKy2�'R��'�'1���f�t4cd�?w�nա��(��	)��d�O����O
����D3J�r���E�j^�19�	�|9�'o��'Lɧ��'"��$N�M��%�KT�kuFW>�:�F�i���]'�8���O��O�˓,,ɱ�E˨� �.Gd]h���?����?���?q(O��'=�� P`Y�� )�&����&�^�rD�'�:7�6�I����O���g��C׌ % d�X �<$��{��64?��Y8�֣|��w���C�qzl�&��o+�h��?����?Q��?�����.��$i�i���׎��>�f|cQ�'��'ʘ��?���Fr����x�����`�q��!�5I�	'q�'�2�'y�ℕu+�6���~�8ŉ��˄q�ɰa��2�~b�|V��Sٟ<��֟\AU�4g �����,�������ߟ��	my�L�>y/O��D=������X*Л��K�uy�>��?9I>��ܽ�@�@2JY�x���(�ؕ��]0	�px"5�iO�ʓ�ڕ��� %��
��.2x8)�t̓ r�3"�ݟ��	ܟ����8%?��'l"���;D�t�A�Y5 ��1j4RQ� ��4��' ��?�$��2�`:��Q9
` t����?���s�@ܴ����B毱?)�O%R��P�O$i
�e@#7�l����d�O��d�OP�$�O~��&� ,'A
.]b"�]=~.�l!�kC��d�O��D�Oܒ�����͓5Dѫ��)�q�F��
(+p�	ݟ�&�p%?xP�즥��b�@���$x�\����)ۜز ���&�t�'��'c
�r���,���ЖᑊO�����'4�'R�Z�X8�O����OX�DF^��uKi�P��틅�\j㟤©O,�d�O��'��k� B�w*`R�jZ�6� ���Cfy�I�i3T4#����4�L�P�2�	7_
�2L^5\Ҁa#V�u<��O����OP�D7ڧ�y2IX����@��.
ًÏ �?�0Y�x��ܟĈܴ��'g�4W]�� ���Z$)����#62�q�Z�nZ�Mې�G��MӘ'rR9gj|��Ѻ;ŋӐ/�*�X���E��r��FH��Sy�'Yb�'U��':�瘚x�H�)��Sd<1`e���)Or%�'U��'�����'��@��l�&$h$z&#�N��� �>�e�i�&6�HC�)��;�n���[�DC�q�QYC�`��c�f�O��hJ>i*O�(ۂ��(O蹚5��7.�`����O�d�O����O����<i�^�x�ɯ|��ݓ�Ri>$�q�C�GU��*�M���O�>I'�i)7����HX��.c��{�N�&,����F�7m!?1���24��9��ݼk�OO�����0閷;����5��0���P�I� �I���F��n��0�9R��F�`噗P��?9��?y�]���Iٟ���4ט'�h��ᬖd(�
�DηC�e���x�'Gr�O�xl:�i�	�l�n�xtxxj kƫ���0��J�F0��g��_y�O�B�'6R�αuQ�X�#ZS��MAP��h���'v����d�O����O\�'}\h�A'�P����'I���'0D��?��4<�ɧ��ɼ3�~�2�Cɉ$Hƫ�6��:��-����O:�����?9�$����rb\M{4$�	���'Z�Z���O���O4��,���<1b�'�v���V�4ji�6���J*B���?A�B��&�D�`}�}�*�A��j�،.��Q�GÐ5,G�nZ;�M����M��O�xr����O|������:$x���N���@`_����'���'���'r�'d�
����(*{-��2��ʹ^U�1�'x��'_���' �7�{��@  #���jJ\�@�g�O��D+�/�	CR;�6͸�\�AK�CQ�!a�͙�\Љ���O� �X�~�|R\��|ᄣʧ ��,;ա�:(68r*�ʟ(�I����	My�.�>����?1��d����ɍ�A�x�*�.[|8Mяbį>���i��7�{�	=fhF�B��������h�>T�P�'�:ܐo�I�PYp���KƟLpW9O�X�̋�<�>�{�+�:ia&Q��'��'���'f�>��taB��&�,v<d@��hm,��	%���<ѡ�i��O�����a�I�!��(\ <c�˅9"d�d�O��d�OD��S``�v���jpN�~R ���a�R�:qL+�� F��'�l�'���'���'1��'��[t�E1Q��QAqO�+10���[�x��O��O<��7�9O�i���9^�N�]/v�aEV}r�'hr�|�O���'.��S�M\ lN�+RNY���=�r/A������,;�J�4��D!���<Y�k�
��X�'UcCF��g�O��?Y��?)���?������\}�'6�)��A�q�����MI�O����u�'N6�3�	��$�O���k�@i�E�=` ��" �ٚft85o�/@60?�q ؼ:Q�|��w-ι�P�K]����=Jq���?���?A���?�����@s�;����H��(̈ڂ�'���'�T����զ��<��6l�N��#���f�:��E�Pd�ß����8s�eM����'��YÑ�M�:|v�@tʽ^f-4胰��������4���d�OX���=��-��-ڝ$s�Ƃ��TE����O��S������	��O���9�f�x��D.ɔb�p�*O4��'�2�'�ɧ��]gT��ׯ��b��DF�4)�tFOF�07�!?���;�	l�I�$q��a�ndK�)�-<����	՟��	��L��L�Sqy!�O� �-�(d)F��7���T�����'��'�N6M0�	�����O�`�D0�c�s_�p	5�O�����Bml7�??���I�c�c?���l9����N�-���B@��O8��?���?A��?����';����d�=.�\ˇ��2*o<들?����?aJ~�_Λ�4OfU3&8Z8�<����2A�N�� �'�2�|����D����O�M���J�el�I�#Α�o��X��'��[��u?	L>y*O��O�-��]�*��a�.[��j���O����O����<�Q�4��ޟ��I��ژs�HQ+�����g�?�bP��Iݟ�&��3b��f\�P�I\}�"��ǈZ]y"B�>q�<-�f�it�i>)���O��I�W�D�B+F !�.��0���J����OH��Op�$<�'�y�ڃ
�6�0DNK<~<>L���?�Q]���'�Z6�&���?݀a\7r �ڀHǧ��qchKџt�	ϟP��sɊ�m�P~r�	�����"LQm�'{�������V�n �Ɣ|�X�4�	��������	ǟx*�D=d�*,Y)��G2h��Sy�f�>����?������<5!�>2"hp�h��F�<(Q C�>!���4��C�)�S�q4��f� 
��qQ��� 4|��$ٖfv�:���`o�O��L>�(O	�j
�X*�8���	N����O����O���O���<QBQ�<���B� ]R�K't�4Ui��о3f>e�	"�Mی�M�>����?ў'��z�C�7l�X�*�+z"���<�M��O�m�G*����4���1�^�[���{g����ʂy��Ղ��'���'���'�'v>�f`�>SS���ߠ3#��/�O����O���'���Mӎy�E�T��t�.W)w�Z]�2������?���?�ĕ+�M+�O뎜�Sj��Asb�&J��{���=o����f��t&�T�'���'�B�'<iv�O� G\��/�V�\��'V"Q��O��d�O���<�Ǎ	WE��7�#O��Ӈ��cy2��>���?yI>���!Z�&�'���A��8 ��A�ǜ�e��lJb�i���?�2��OГO^aʳ��>��	�b^�xN������O^�$�O�d�O����S�rQ���l�^��0��-�?�)OƝn�Q��Z��	Ɵ\�6l�0���@%�z6�P���ݟl��e >9n~~�%L*M$H�~��D�M&�����&[��h`�a�P�'�R�'	r�'���'d��>\��s�̚H�`L0�������'fr�'����'¸6Ml�Li �B)T6�l��FI|��ҵ��Oj��(��+�� @�6m���Y0�T�]���I���&vr�-��ON�����~b�|�V��Ɵ�Zǁ��Ԉs���mq�G����T����D��eyr�>���?��)��,"��:B���jA�T�@�z�#�r�>!��iDN7��u�	�1m��!��:3E���5�C62���'��x�-+��4c�O�阞�?9��o��R���	5��!�K�S%�Z�2�'���'*"���<� �4OX h+�$�C��L���Z���s�O��D�ON�lZ|������ןm��+%g"(Qv1�Q��?����?� �i!>�ói���O�@	Dʳ��]w�@L3#�T�e�"�\�E�m�O>�*O��D�OF���O<�$�O��*�����Xy0R�ۡ&.� �<q�R��������k���l�vg�m1�� ��K�ZMX�8��dCɦ�ܴʉ��O���S���h+�݋�n�{�<���.��$��O�U��_��?1G%�d�<Y!�C�P��nH�\nv����"�?���?���?�����W}��'���e�����P� ��-�#E�?��i��O���'�2�'��dQ�z J	�#���CLA5z"��ó�i���1��J$�O�q�(��%HFT4ɜt�(�z2 ����D�O��$�O>���O8��/§>�B �ŝ!z�V�rFb�A,ty�	�4�I!����O����1�<QR�]�h��lyw�^zJ
CM�����ll�T���'E>6??y��U;=����ƃJ�Hk�!I�"��	�C�Ot<�L>,O���O��d�O�dؤ�������dA�K�2���.�O����<�X�X��ٟ��	g�ĀD>X/�L���$G;����#�
��$�T}��'<��|�Od��>&�n�jd���D�Y�Mf�Tcb-��������6T��$4�$�!)��㔎��F�_(A|���Oj�d�O���*�	�<�s�'aP��E��T\ah�W
l��ݠ���?q�hr����\}B�'?D�⠅�0U2� ݳ,0��sg�'�)�->H��?O��d
~4�L?牔�� �0KR*F#�5P�k]0@����By��'��'Q��'W2�?�Ц�J�.�̚�^x�x=Rto@E}2�'�r�''��5nZ�<��EEl� ���82PlX������	P�ڟ0�	���H��̓ J`�)�L�-�c��8(�-��A�ẟd$�������'p
=A��E�c�2h����QUJ�B@�'2�'�rP�@�O��d�O~���ip�MI2ύ�p�x�Bsj԰%�P���OFHm���M���x2��-��L��M�����K#@B��'�d�3���D���O&�iЩ�?abh�܁�C��6<��/�}���e��O���O���O6�}Ҟ�� :t��Z+U���QWNКό���'b����d�Ǧ��?���1�,�c��у#kb,�v��dU��b�?�vLmӠUoZ�3lnU~B��9֬`��$zL4��DJ/.h��ֳxU�����|"\���	ߟ��	��H�I�$� �E�-�lsB�2e�
��sy�ϯ>)OB��;��>K|�-�'TMFxc"�F:]�x᢬O�<l���M[��x������J�l�����U��	��B��@t�	�&�X �'��%��'~N�i�q��$�����b�'�"�'���'��Z�b�O���yl\}daI��!�c
9�p��^Ǧ%�?�Q��K�4囦C�Oƍ�#cÓ0L������Nz���^:y���(���Zp$��$�Q�ʼ�HX��蕥Ylڅµ�ȟP�	ޟh�I����	Ɵ�E���ΰR%�(y f��3a��$"]!�?1��?!U��	�d۴��'|����aۮGgZhA�`�&��	�O>A��?��W3v��4����x��b�Y����k_#Y��5�G�{��I\��|y�'���'�r�o3̩���s��9bG�w��'������O��$�O��)�.L��덺.�:���X��'����?����S�)F4��b ���7XҼ*1fΤ`�b�A#��ݛ��<�'O�d�IV�I����Ѣ���,��������Ο4�	�(�	\�Sxy"��Ox��wG8	���Q�~1�)��'u�I(�M��r�>�ջi5� ��!���3ͅ�1,Naؐ�j�6�oZn�Ftn�p~�a+��Ӫ1&��=�ݙE�xILmh��7H���<9��?9���?Y���?)˟ƹ�FW�G�t���G`+�m�To�>���?9�����<郾i��D�=\�!j�a�!|����5`T�p��6���a�N<��'�R��1v\}bڴ�y¥Yz�:��W-Y�X�28�e,�X�����ʔ9�i�O���?!�f��ŻP�(3�`��H�[^�x9���?���?/O��'}��y'%�C:%�m%5{,M2�<��O�)�'���is(�O�	���?���XQJ���RtJ'�'�2˘�jJ���,ť���������NI牓bK��[�:��<���������Oj���O ��-ڧ�yR�4 �c��**<�s�H
�?�AP�T�'��6�'���?��ׂΩvb-0�X�`��E柜�	�H���	�� o�<Y�� *����~�T-ذ6~p��.&X!mf�Py��'�R�'[�'�R�Ğ ��PK��9ia��+�Y6*~��:��D�<�����'�?y�dN�o������5����o-"H�	�MS�i��O1�����%aY� ҩ�<<��$K�N�(z�HP.H�	�d�I
5�'���%�L�'z��2BEr|�!JD�M �N����'��'b�'f�S���O��$� n&}`�aI�/Vz�(�fQ>j�X��YǦ	�?��Q��ٴ%��F�O�a7$W�#~B��Q����q ��[.U�v���)vTiD�4�)b��v��g2؉q��3f�ȌCP��O��d�O��d�O��d�O�#|b�l�X���r� \Kf�5%������ퟤ��O��d�OԱn�J̓EJ����@:G%�)� Y�"���IL>�ݴ8F���Ox���лiB�$�O�,��gGZ��1sӃB1	N�B��D����2=*�O��|����?��s� @[ #ԏ.Lhp�l 5�T��?)*O���'Z�����OL���H�V�DT��!_?~��-O���'��'�ɧ�ӀBB�D�UM�(��M�F��1�F�&d��x�.��R�����?��Fy�Ʌy���b��c�]	WHO-�	���'���'�"�'��O��ɷ�?9�E��4���2��@��ğ0�'�X6�"��0���Ot�v�Bc�"�ʅ�,Fv�j�B�O(��!u�7�:?�;T�<���O���5�j���Oq�T��DG�� GZ��<Y���?���?���?aɟ���@�Y�PH�gi�g�ꥒU��>����?�����<u�i���׈Xu 𚔧C;M�I
��Ӕ-�R�'z�'��Os�a���i����(U6��
�$�hNµ�be��Q����������O�d��H�pC��,A��r�U�#����Ov���O�j
�	�������A��b1T�7N�	~j���f��4�����IL�"X|�'�Er)��3Ԃ9�$)�'2�����sS�&C0����~�8O�XJSꜳ nP�rC�ܓ/?�MC�'���'���'��>E�qO\�7ƒ��T�w�Y�$��I�I	����O�������?��� �ٳ������i��kR��ޟl�Iߟt���+6Έl�v~Zw��crߟ&�����L�*e#�)�*l���8���<1���?i��?I��?9Q��iP<�J�" ��n%���'�b��?���?QN~���=I���M	�!�у�FI6=���T���	���%�b>�X��ъ�|�EĈ�,X�b�Eqndm���`�(��'��'W��7|�`Hp�ޚ����&E
Y�"h��՟��I՟��Iҟ�'w�듦?rL��=�����C�'�ze�� ��?!�i1�O���'��'.�D�mL&�)d�/T� �
���[� 8�t�i%�	
N�n9��ݟ<�����Z����l A� N)�.���O@�D�O����O��+�g�? h�%ݸzc�@��S*ʸL���'Q��'r\���ߦ��<)��Ŏ
�ڙ� �6N�@m�SM�j�ޟ8������'�ΦΓ�?U��R�[���� ���@�!���0�饟 $�������'�'_B4��k�*nYK�e�1vD�qiu�'��W��ɮO���?aʟ �&�
k�N��tK�'v���� Z��+�O���O֒O� ���E,�A�h�����Ja��/W���ne~"�O�^����N�j1z!ė�m@�X��P�$t����?���?-�M�M~b*O*-�I�(b`��E��R�|�GH�g�H�$�<	�iK�On�'��$�=P�-�4b�]S$C�,��'��X���i*�ɫGi�A�	D�r�p8����.^c�)r�aE�H��Z���	ɟ����p�Iן<�Oh��3� �~,�I0��P'��9�U���'2�	�禕ϓkD���D�_,i��<�D���86��	���&��'?A�I֦��Cl|s�Z.+�9z��2<���	0G�e���O��O4��|��C�|�	�f
�9�� �)���Hy��?���?�*O�|�']��'cbgJ
G25٤e�
_����C4`�O�t�'�07M��uYH<9RaR��Lh����vd6��������3����L Ȇ�������"Ȑ�I�y�ax�D_p5�ၣ��V���O���O��D.ڧ�y���m!�	��)�PL�yp+���?�Q���'G�6-?�I�?�w�$��K2��3lՋ�A�ԟ@�ٴPH��gc�0sGf�x�?R�Z'��DqҶ��kv�(B�G�0تl��
_������O����O��d�O.�dҕd��hh��~���CTe�I�(ʓ2N�I��\�Iߟ %?�ɉ�h���BΞj_R|a�f̬KR��[�O�Qoڷ�M�U�x�Ot���O��u�(Ӂ)U��y5��Y HƇ�2	�4R��xRnA�r J�	gy��P�\�l��ӃW@�`c+��F�r�'���'���'�������OVm��b�*#hH��8Q��L �G�OȤn�L���	���I�<-U�N(S��>Y�q@K��%k�����h�
����T�i��}y2�Ow󮞨&\ ��nC3���3R&�[Yb�'�2�'M��'.�ᓫ\��A�Pi�^��\�S'/I"���?r^������4�ٴ��'�>�� E�]6�:������M>9��?��K�,q�޴�����ؐ�9NvZ\����'&��0C��

 ��I^�IDy��'s��'.�ͻV��&j��}/@y�$Ş?]�'��	����O����O��''��$8!�C�4u֍�Ы�s�(�'����?Q���S��� IK���c�u`uأ��^����./�����<��'m�t�	E�ɷ.6��:��B�D���X �Gנ5������	ԟ���|�SFyZ���1[0�;�,cQ��K"�'��a�b�dp�O~�D
�>�����-
�*T�F"����D�O:��hn��Ӻ���K���?���ފ'��X�CE�xL�m2���O�˓�?a���?y���?!����ְ16�d��i�?�b ��X���?����?�O~���S���?O�愋�� t@rN��=� ���'��/ �d?�I�t]v7M��:��"-��򂨞*k<�tI N�O����BX��?��-���<ͧ�?Q"���8VX۶��7f�"j���?����?�����DB}2�'Vr�'�m�f��*K��M@夝�h9��YP��MW}b�'_b�=���nМ����MRg([
���wo�`& A�Xu6�����ßP(1<O�E�Ӧ¼F�h��Փ�����'xB�'���'��>�Γxg:L����'A�`�X Ě��8������O��������?����A�&#�� ���1k��&
�9���?	�����3,Y���А�GU�����D1���=sԊ�Ud�n8�D��|bT�x�I�d��ܟ���ʟP+��п(���aOE�V�|P�doWAy2��>����?������<IU�����OV��F��`��27��$�M�ihO1�8�kw��?"�aǊ1{P<x��I�_�҈��i�<�X$4M���'>A&�P�'�f�h���Q�a
�/.kd<ѐ�'��'���'EB\��k�O���x���^7@D�m�%��5�������?�bX����۟0�{�b����L�q���w�����J���'/���f�c�O�� >4ڍp$UJ�鑃S�AR�'\"�'$��'(R�F��t\�M�^�$���w/��$�O���PL}�V��ZٴƘ'Q��"��HJjQ)���6�N>i���?��?%ְ�۴�y��'ˢ�"uH*_��4[�+�iy�I�^L�8��䓤�4�*���O��dA6i��T�f���WkH�!Q�������O�ʓ.��	ܟH�I���OW�ͨEă3\X��T�/>�T��.Obx�'��'�ɧ��m�ཙ@'_�)�f�����w%�Ы�/��{:(7��Ny"�O������O���˴eD:t/:rW��)�e���?����?�������� ��,l%�͒���)�4���O`˓]����W}B�'�"#�q��`	�D�"�>0��'�-�"p/�V>OD���q��h�'��$�N�P�6e��n��'��D�P��<���?I��?���?Iȟ� FiH1�X�ck�a5�޲Dr�(�c�>y��?�����'�?q��i��%1��p�H
3Bp @##�B��'��'8r�'��a "8]�F2Ob��E9?�P�S�ġU�`E���OX��@��.�~��|rZ����͟���x3��W$� ��Kp�DƟD�	蟘�	ny2#�>!+O*�:�4Y�$���~�x�^�[�&⟘z�O�]m��M��x��B�a�@�� _)���S��I�|���r�H��C1�'?�j��'4�ϓ.p9Ҁ*�3NXtj��ݙ"��������	����m�O��@�v\x}�"�܀�\s�J�?�b��>,Ol�_����s�uL����K
kT0ȣ��;�?Q���?��aŬ�{�4��D�=�l��'�b� �.2��,���\�E���2�)�ļ<y���?����?���?�W�W�M��=�(D�@���)�"��n}��'��'��O��LB�5�N���)]�|p��I�EG6b� ��?����S�'B��}ȁ�8�&,�Pf�7��|��6�M3�O���]��~�|�^��YsO��o("a�O��ɄM{���X�	�(������	py���>��bp���kW	2h���r���j��X����D�o}�'[20ODI��MUv�e�ܯ7�X�K���Uy�����c-]RQ>��;r�����/��`$N ��(y�I��P�	۟��Iԟ���R�O����Aa�!Z=�mC|�
����p����ĭ<1�im1OzM $�ɇi�d,�@Ñ�!��|���|B�'���'e~źƸi��I�^C �֭�,6)���%A�_��P�Ͷa�2��n��wy�O��'�¯l������s�E=Ӕ�����?�)Oȑ�'�R�'�?Ys6�?T�[0@�0d*�Φ<��^�0����d$��OnH�T�����ION�:憎���&�[P~R�O3����� ��'7���&M�r6�9ʗ
M��5���'���'���'��O��	%�?)���5D�uR`�ײr�2��U�󟨕'��7�.�ɱ����O�
7��2��X�$��� A��OR��#X�7)?Y��*i ���&�� ��,9k�j�?�X$8�,֥�b_�������I�4������Ow��r��E�pH`h(����p�R�CwT���	���p�s���4�yRa�h� �a� 	m��:W��2�?������}����4�~���2KY�kY0`�zE��?9�D�~����+����4�����'n6�Iq/�O~�8jP�P�Eb�D�O��d�O:�tX�I̟|�Iϟ C�Ɨvv���&׊9�`�����a��0����M���i)�O�@��#ϻv�bV�]�2�@\���<���J���4�r->��'������y�E�s� <���;VTh3�ȃ�?���?����?	���o�pr1(�' �N���兎q�:�kGG�OB��'-�	�M�b�O#��u���
`�wO�����&�''J6-H̦���4*$�[ܴ�yR�'�A��o��?����U8��]F��G�0X��┲r�'��	�������͟��,2!��o�6J"s����R�T�'���?	��?II~�ՄQ@GJE�5��A�Kӧr1�!�w]�,��4d��vn&��IO$�&o˽{��S�Hv��ypKkR�� q�+�!�O�I�J>/O�D�գ�[��j�BC�c��S�o�O���O���O��d�<�^���I�b3	HLP�U�i���1Q��m�I��M�� �>����?��'� $W2J�
G�SU�\P	��)�MK�OR�BB�a�E��2�:�C�L�>tb�Bs��n�=#��'2�'�b�'D��'9>�)�A|3N�;Ê�D�.M2��O`�d�O^M�'�I��Ms�yB��>���s�x�f�����>v�'�7�NϦY����J l�<��tJS��4,��̓�JY0�8��k�u���ͼ�����O���O��DI�2j
�A�S�Kl�,y��="l�D�O˓Z��IΟ8��ӟt�O�l�wi]U|]��mJ-<
��P-O���'8��'�ɧ�S?=��$7H[`�B�æ��f����B�YR�N7M*?A�'aN�	h�	07�8�b���k8��Bd	 �B��	�����	n�Sby���O ua�֌B��P���#KꠌcE�'�B�'D6<�������O�Ճ�Kу]I�A�� �8Lj�Ɔ�O���%[(�6�=?��R�#B�c?q�5��{�.|T� e��� �c�O���?��?Y��?�����I� ����V�ղ<ښ��`I?����?���?�L~�,I�9O�����C�,0���_5p���S�'���|R�����nܛ6�OzD�f��&�����+ИX�
!a��'$�j�]������|�Z��SПx@[�
T"-s2�-7l��¡���@�I�����ey"��>i���?y�.�#�l��������s�]h��>!���?�O>!����\�z�QD^����u��$�O� �D�ޡ?�@1;����S9Cz�
��<!��E�(4�0Ջ�r˶��4)��\�I̟(��͟�G�d=Ot�����zL؛�ꀛm+�	v�'>������?Y���
�Òn��f  � �jѱ^_(D��?i��?���M��O��v,���z\w��M��԰R��F���R�O>�.O��d�Or���On��O
� &1���\��Up lָ����]�8�O���O��d=�9OZ@xTA2r�Y�!�.���P�D}2�'���|���;P��`wON�Frx YE��=��!�iL�ɅV�|�O�O0˓{�E�ł��>��I�FW�f�x��?����?A���?�,O�Q�'N�7{���d�(9 �t��
$WC�o�`�tҫO��d�O�扬� ��G�
���ti�d|jeq�hp���4;\�10k'�'�yW�ϊT�\eQ1l�? \��u�vc��'5�'���'���Ӏ!3 �Ss"�52��
��&SB�d�OP�N`}R�ܡ�4��'ќݰu��y|!��,w�|�bM>���?9��^j�z�4���T4T7*��	��w,$p )̞z��J��O��~2�|�W��Sן���џ�ӆEoh�A���ړϾ����ݟp�I]y�E�>���?1����3$�"�Z��X		:Ti��܆I�I����O�d?��~��1�Ԉ�c낞 q�R�(L�!.��s'�٦ݒ+O�I��~��|���uR�y*��rF�p�O����'Y��'"��P�@��rH�P �H!'^�ӒgY�!�T��IEy"k�:㟐ӪO����=h�L��E�>�t�dbQo�f���O�M±�w��+S�e��F/�S�NVH���Įs�R|�`��b
����<A���?���?i��?�Ο�����'�̉(��Ŋf��HRcJ�>���?������<)V�i���^�|Qp؉�#nVn��(¾[��'2�'q��'t��
*�v1O��H�E. ��I�@f��DȨ[A$�O�2�؄�~R�|"\����X�OJ:G��8S�J�>Bx��A'G ����I�����[yȷ>����?y��S�x���>r�4���7M̕��̣>���?�L>�7c߄B���j�*�V��q�.����Ѫ#`X���.y����|2eN���ϓ0��!č.[ꨅbUO�0C�ru�I۟d��퟈��j�O��D��^f���A�pcd���K'��>9��?i�iD�Ov���u�� ��(5�ԉ�����2�(�$�O��$�OrL��sӆ�Ӻ� Ҽ��� �-�<9��인*�B� oJ �'��I��0����x����l�	�@��Xa�E�: \�Ȣ�[9Q(�8�'�`��?a��?��`I�]X�����=m�hq���8I���?�����O:  &-�B�2�Wa�&bLt�7��^^E �O8�oĵ�?�@">��<���5WD>�A��T&$�6ݚuf���?����?���?�����$Nj}"�'��8AܤH��	���i�p����'��7�?�	>���O��dq��y��a��Y3��L9�y��C~+<7�&?	�A��>dT�)9�Sۼ�EˮX��RtfD�TSD�r ��ӟ����T�I�8�	��G�4OW8<�؄!�-l\ɚB���?����?��U���'�46-/�I�O%&|hG#�E�qwٱ �
�O���O��:7W*76?�Y�,�3����Ex`�i�،��Aa�O<�SL>-O��O.��O��5o�J<L`�!H�l�$�@N�Ov��<)�[���	ϟ(�IA�t�˿q!���a@=l�`G/ ��A} ~���nں��S�i޾�J���"ǀN@a��Lo�<�ӡ�	ktB�HГ�l�S��2�GP�	�94�T-��A����:Q��}�	˟����(�	L�S`y"a�Ov�F�!.jC� :6ǲ��''��'P78�����O���$I�z�S��U�@kӐo�a>�m`~�d�?I�|��ST��+~�j�nD9Gǘ}��%��;��d�<i��?���?)��?yȟ���NQ�Xx໶��2�F]�P��>����?����'�?q�i���
�e�8V��u'6^O�ֵi��6�z��_�Su�N�lZy?ђ�21�� 1�)ߠ>C�Y0$�4SC�B���e�IVy�O���Ҹ#k��u�ۅ^I|A���:|�'�"�'~���$�<���+�0X3dI_�B���[��e�X���)�>1s�ie7mPs�i�u9�ix��yӎL#.��Q2T��aC�|yZX��F=?�'7�����:�y"E�{-ҷ��|EY��?���?���?Y�������w�\��ʣK ����b�'����?Y��5y�V��矊�pc�
�� q�<rԝ���j�������ߴ&mL)0�4��� �Tr���'�uw�_�Uܦ�+c��sw4�JH�&������O ���O���O��D��(����f�d�ڦ��2�f�E<�	�����㟈&?����C�X��!Y�e�-����I��*�O�%oڪ�M��x��$��.F)��P�C�[�<)��
B��r+����$�	������OʓjxJ�B6gߕ_X&@J�a	]0�t@���?����?���?A,O���'��Ȑ��(�[��h�&l-��X��'�,6�/�I#��$�Ħ)����'
����$I�C*����Ʃ?�v����Y��M��O��M���47���ЀW��´i����S�B==��'r�'T��'=b��-7�zX�o��T�nٰ&7U�J�$�O��A}b�'8Rf�*c��y��<ZP�@�a�bCr4�V"�d�O��c�0�w�v�x�4��G�6��T�aF=j���i ͐�p�~��h��xy�O���'��� @�Ҷ��Ms8̂���~�Ӧ�'�"R�(z�O���?a͟�MJ�ٱz�X
���?�n��[��r�OF�$�O��O�')8�e�Ϝ�W�V�{�O�"^Qb��b�X�-n�B~��O{n����?�l�PV�Ӥ��#6'\&�l����?���?������DW��:�Չ-k]��߳6��1�F�OP���OD5o�~�z��	ğ�����Q��U��k�$=�&��Qʈݟ��	���l�l~Zw��i��۟��'`@V%�1G�*}6�-pN���젉&Wg,�2�ߧ�|�h M�rf��E� i����M��Ɯ ɧR!�ꡠD'�6������~��p��ͥbD��� 4}�ى��ȶ��X%e�t���Hvb�Q�s� �#��lR���sĉ�[[*1��)�*"���!�%�{6�)f�$��|�3K�Xn
lѦ!��hvѠb+� 6��y3�,fؓl��=ư�W�=�� �U�7��ɻ���%j�;��6�o��!��B��)�Vx	�柪 S.ꒈM-d����Ͽ:t���rd@�$��d"w�]*�K䚠4k^�*�J#x;�%A2
M;¬�Vc8؅��(�v����Z<1��׈r�`t���Y�����a�+ݲ|�G�E�$z�x��J)[�̘f�0�*c�E���Qc�?���	ŎN6\xB�&�6z`�h`��d�Q T&~}*M b��5�a��Qt(��%�*B(�b��4i��A��ڲ��ԮE2@A����o��=rBx�0���O����Ox�'3���|�<���%	�~�h�q��'s�~��?��h\��?9��?c��A~����i~������?��?��W��'���|2��ۜ�)!�Ú$f��᭐-#��	!^ބ$���	ן���w����>���Qd@��Y�2��L٭�?�Y�ؖ'�b�|��'��H������,�T���lK�C��e�!�'������I͟x'?}�'Co�J"-ʷ���3f%�e��L�	�l�Iޟ�%�h�	ޟ�����[�DA6P\�x����Dv�i��`y��'"��'��O���?��i��W�u"��I�+��Y���<q�����?y�KS�5��y�b�=(0��wNR/(�HL��GR(�?	��?�*O��d�J�T�']B�'[fds�B�U�J� "�T�Tt:آ�]���П����Z6�����{>ٰĮi��\��]����g��O(��?����?����?����򤒧f�"%�f�`�V}�Emġ	�4��O��(2�D��>yكc��^74�R�׀dC0�p%��O��D��i�	ǟ��� �O2�%�ء1X�>g���$r�Ah����Fxr���O���ڵR[d�23gZ*}�ʄ"m�����͟H�I���	�Of��?��'�"rAG	nPhP6皞�F�Q��"E���'���'���,�2���l
T��]/p�p9�'���'7����D�O(�O�q�aGC�^�̫4��1��� �<ɇ���?�+OT���O���/� ��"[^9�⠆+E>�1W��؟)�OV˓�?K>���?yg���$6�H�*<�5`2 ��f����H>���?����������Aq��Elkz��@O_��?))O���&���O���X�ʰ��#H��e�e��I���� �>�ʓ�?q��?�J~u���l:��k3��?}�\`�N�>8B�'��'9�i>��Ip�D�!W 1�u�n���hC�8�?����?�.OD�DU��۟��;����Fƞ<]�$��!|�Ν&� �'�"�'V��y���`qJ!�V����b
�C��^����%�M[/�����O�L�'a����d��A�N�% �e$,x������O��>�	4��J��ҥ�ĝ�x��G[�=�˓�?���?����?!*O�:&�}1hZ=�ܔ�!@�A�V��'
`����Ӻk�8�i�N�x͓U�.�4��՟��	����	CyʟZ�3�ȵ�j͞F��1õ�ύaPf�f#��Oy�6O����ӬF%���A�,M��Y��':b�'��	P�t��0O��q�
bAA\�\����P &���"#]1O����<��'��b�
�[}�)�����Ƶ�������O@��?�Iȟ��P�>��@W�c���SԫA�4p���q��?Q���?�L~�0�Or2t����<1��=���S(g�\1/O���O��O���|B��l8 �w�:�P
���2J�p8O>����D�</���$ޝ���YbA��O[����ѹ(K���%��񟴔'%:��K��r��'S�&�7�[ Y��a���OH�d�<	/O�˧�?����yW$Ϊ,�x��akۻ9D��M ����?�/OL���I�D^�8�mI�^A������!Q��cy��'X6��|Z���?Y�R���랸\Q��2���ۼ52&�O���?����'��{̾��!�	$�l�e�>a�D�s���?Ǽi�2�'OR�'
�O��
1�6���ɯ!��8`4KC�0��'b�'�ɧ����j�(2�& �냸C�0��Ӏ����	Ɵ�����ԗ���4?�6����Ff��oK�5�aoN1<N"<�I~����?���I�<a�F�?e�`M:�J1?�@*���?Q�������!��Q<cb$dx���1@�L�L	]SH�O��$�<���?�����W�~t�D�d�E�{Q��C)?q(�d�Ob��3�D�<�� bhw�ݝM����%��q�R\��'�]�|��ޟ��It�S*��S��*
�HRa��o��'Ly�'�R�|Y��ǟ! 	��Zؒ�k߮<�����O�Ky��'�r�'/�OS��'�?m%O�d��6�F1	���?������OV���Ovh����擿b�,�i��;D�q@)B�(^�4��ȟ��I]yB�'�\맾?���?)��Oa�P��� @2�t�
���O���O � �;O��d�<�;\&��e��-�p%�1�Ԝc�V��I\y2�'̈7��O����O&���q}g��S�ТAo^<:���Ȓ@�8M`��'����6��ģ<Q���nL�J
���%F�������D�?��WX�f�'�r�'tbe�>�/O*��p�B�2J`�1f���u!��@g)�O���45O��<����'Z����B�v�V8R`��{�d�Hׇ~�����O��O
��'��I�X�Ft:���� [r���*�6)���	ɟ�'���Ce��$�'�B�'#t3ǣV�r!W��`�]��'=��'�>ꓻ�$�O���y��B��V�ʥX�`K�e� ���'k�I�'����Ib�'g���Ŋ�$]*(kf��C�L������D�<Q����d�O��d�O@��P��-�VM�f����>����� ��$�<)���?y��� �db\��Z�6IR�DS�Y����?(O���<	��?I��tU� E�ŉq�]������,��!�	ܟ���IBy�OA��g���%D��`2�U)Y��L�k@�����Oy"�'�b�'J�9�Ο�牰4��
�HQ�g)fT;1�mD���Or�D�<��7���ΟD����X*"�W�@���P2ɇg����#Cy�'#r�'���'#�'�C36�3V�T�Ya'�Y�B�rS������M����?���?1�\����@��h0haAj_�G:�d�������֟d�b���IQy��	LS�aR$CE�h��M*.�+�R�'�R6m�O����O��ĆJ}^��h�ΜBv��� ��NI��l���q�.���O�RF�_o�j�E�&l�$MKC_�7m�O��$�O���x}�U���	�<9��x�$�bg.Q4��'G$�'�bˁ
	�O��'0 δJ/x��C���Pi� �8���'d�,���O
�0���vR\V!x ��mU�#˓a���<a���?y���ɔ$Ir�<3�`��!�ԯN����E�'���'��'���'h�"U�)v(�!�x86��w"ɂW$�R���	ğP��J��3���DA���XqQ�G��x�	XFyB�'R�|R�'Lր�~҉K'%�f`���1-(�ʐ逫����O�d�OX��d�$>-�bO��snQ���zV�P����,��U���(�	�-n�e�IL~�+��=��HɣC�#(�
�������?9���?�*O��dRa����H��d���&�р6^�5IB���L$�0�I�� ��E�$�H���̈ .U��BO�<�2aP���O�ʓ�?���i�����\��1��d��O�Te�����M.r4b��ʀo��'�rc��y2�|��ɓzviq7�M7BOI�%3N���'��6-�O����O>���[�I���	1��Ek\��Hʫh�,�$���`��ܟ�&������T��S`�"�p����.#b�LJ��iK��'9b�'�2Ox���O��H�Ra�@B�w^~ƤL���5�ą�S��<���?i�w_�F@+&���8O@�H! ���?a��O�'���'��'��3�	�O���p���,TH$�_���HI�X�'U�'�r�?ہ��?kZ�hr��9Za�4��OH��>������?���1S6R�BD�.Ԕ���L]:�����<�*O>�$�OH��+��B�?ə BR�.<`���ƚ� �<����?�H>���?��,��<�����3��y�3J��N2>�+��;����ON���O���$>�����C@֤*��ޤ�����d���	n����		���{~R#ڽ9��
M�Ggf��&�ո�?��?q,O��d�v�����ɘ �Bd�2�hH�E�Z9OW�e'�L�	������<'�`�'$��PBPCó]"B5�b�Z2
q�Iey��'1.6��|r��?�FQ��6C3��@k�'��=��"�<�+O��<�)��@""�T
��"�V\Y�V�?������'
��'1/1�4����A��O�6����\�q�6��<�������O��M�,�J�����pp���P�^���'��	�`�	���'��8O4�l[.1�<�z�%I��<�b���O�������O4�$�%�f,�VA��pG� +n���O��D�A}����'�I�
�nm1½�EN�$p��@#�<9�ʦ���?���?����D[c��"�a,*�6,�XN��	uy�'B�'��'R6O���QhH/�N�C�	n"��'zx	��O ���OF���Ob�'��ĭs*�{a�Չ%���-��?A��?Q��䓖?Y)O��4�R�2UyѦU�#1��b���ʓ�?���?�K~r'Z?��I%Q�5��În�6�K'$[.��H�Iӟ`�I��6��y
� ԙa���hBAN�8${�l�5�'���'���'�B�'��'y��'���E�9vK�MA�B�\m(MK��|��'l�ɺ_&"<��GV1��Sr �4�x�ɷ� (|hٰ���=#
�t����vbP`�
,��C�'�u�g�����(.�8�/k�a@�j�-�ēOV�d~�|�oڋ�?����?�����
T%�%�]�\�R�F;`��?��K�lM��!BT�CDfu�iE���!�6l5X%ۯ*����%�'K*Y;7������JBR��(q"��I��\8�ֵ�8a@��	3ڹz��͂9�H��AD�Da>Hp֡ %eZ!����6	l���g�m	"h�`��2�0ʳڀ�5���S�
_��[fI�	NΕ�f	#9�{*'	�̡;�eQ�]�����	���3�O�56>u{�Q8:�,1%�|���Ȍr:X�VH��yg����BϞ0���X�N�\�n�x��4s]ؐ���:@�ӥN@z@m�ğ�lZ+x��`�VP�1c�HBJn������H��;a��	�b1w*�Z��$�`G�,+����0��hA�!�Y�P�k��]�
SLC�{��E��EK
\�1�TF�=/k����P��dQ�22�'��)���>���>�8�)SČ�!��y�ъY�<Io�>˺0r��JFrp���
W�'��~J1I�5��8"Gΐ�q�<�h��S?���?A�F��$?�6�'�B�'X��	�h�Ia�
�$E���`�&ѳN�r�}o΍��a�����'��) �Eͷ#h|8�����`	������	W��i�Gh�3�I��sdn�\�(G�ˊ"%��Oڵ�!�'-����	��"F}��'@H�n)���$"Od�{G�R9[��]�!�0,�~8z��O4$Ezʟ�˓l���w�� � ��N�S�ҁ�e�I8y���'Wr�'��I�����|���&l��G2u��l�A����hq$cʡbQ��Z��B=��<���;U?���	1cn�A�/�r����Sa+,I�:%  ���<�ca�)���ʂF���Ф��'W2#e/�2�?���7ғ8P�
U��!䒨�&�#a0���aւ�;"�νe����Q,G�̚,�O��'��I*A�Z�ٴ�?����M��!C< iH�ؑ�7H����t��O�I����hX�Iß'��n]91��1�)D�z��ȫe呟�dN��Y��sŭ���鉝mQ�4KQ�� )Ð�b��߯gǑ�`�r��O��$^K���\;��z�(���RשJȾ��I�?E���@5rD�A��$[���8I�V6���ذ�)§'Ǜּi������E0����ᑡA�&�p���<�㡓�e���'�ҟ���'ћ�&UZ��C��]Qv03SB�)Th��
�C���HWb�* 
C�ԗ68|p��O:�O������9Ct�%�K�o�A��Od}0A�I7:+�4�)V&t��I��aQ ت`3�e�����)��d�䝅Y�6y ��F��$�, �	#�M+�i������O����	�t��=�1m3�xu�W�i�N���O���)lO��֭ضw��Q#��������ɒ�M[��ir1��u��dE�u�LU�F@��iq?	���t;�+�7�r�"&�G�}�%�ȓ!��P�����K�.��ҫ]#PZ��a�lΖk���tS<��=!�eZ���ŮH`YP1�'�Gi�<	�홚K%��c�+�;	�h�[�EOa�<Q�ԭL���Iޮt)\�v�GK�<Y�.��Y�T�a�i(D��̸�&�F�<q��F�0D�t��e�*&?�HX2"|�<�����{��,9w� ?=ܑ�f�t�<1e���!���2��5V��x*��j�<�AH������9���\�<9rI��M��Y�n�5��Q� CX�<�$*�+1�x�ʓ�Xk�B���a@W�<GdX�<���c% ;1��I��O�<d���bļQPIY7���I�N�<�J��f�X���1Di�%�Sj�Q�<�"��b�Εa�Ŕ3�6H�̚S�<��]"���C��e�N�+��U�<�S��yRy��@W��qB!
[�<���ҳcm�` 7�
�4T����Iz�<��ꕚ/�|�!�8in2���R�<�æ�=~��j���\
���A+�q�<�S���LY�ћ�hZ75w\�B�#�@�<	tN!P�, (�'	�����H�x�<9D���"�@ 
e�i(�倳	�y�<yr]�co�E+У�.�qp`��q�<���-2H��`�;E�X��5St�<� �I�����rNf�]�P���QB"O�M���4P�>�@W�L���s"O��rB	�(8v���n^y�����"O�壠�}�ZP�Q�H-�B"O�E�`�D5�h�K�d%��"O���dHޞP|l��l��ZG�eJ6"O�6i�
a�@�1�$�E).D�� ㌊]7!���O8f<�%a D�hȧ�A9/��ʳ�=4���!D�XUϖ����а��:w$����(2D�p�"3Cf|�gO29��� ��,D���pd�f2�9��Ɍ2.��h+D�|��+ܠ^ܝ��HF�k��];�m)D�,��f� Ȍ9A&C[�d�ʅ�ǩ-D��(�F�~Gd�q�oL!22(8�	+D�Ĩ#O-os��iK��923�"D�\���Ͷk9Z�	 ��M��j2D�� 4��T(�c���$0}*İ�
3D�83�&@7
�TA��.��`S�գ��2D�@�+�[��(k�)l�h�3D��0��E�S�fp�	}Shp��);D��x�NWxW��b���*�J��l'D��@RAV�t���І��CIV 0�O8D��(S�@6x4����(ѥO]D<�W&4D��bO��]��P�/�N^����2D�,�L'T����)�%�\LH�%?D��L�7
P�K"�ěn#�Q�,/D��S4��#B���s̅��۶1D� ���-<�IQ!@3G頔�
.D��Ib��.�d\��^�w�@5 ��.D���B��KQ�=��G�A8�R�!D�����]�t�5&ɛ�D����%D�����׮�1V��N|NA#v�#D��bÇ,�:�ٖ/����=*� ?D�\��L�;q{��t�AF�M���=D��R�d$F�}##.Y���Y�@ :D�p��A� Aƴq�Ԯ'��hpL<$�h��	�'b&�QC��y)�h�I��y�Gͼ-�<rU/�O�������y�%�63��f��m6d�s����y�$��t�
�� #J�� ����yR�VN�481u�р{�����4�y��$f�RQ���s������ŉ��'������I8���f�#K�b�8����1���x3�*�OXyg�P7*I����'�ȱQ��94�`�E���?�v��YXftZ3c�39��� �`�'��8��ˍLon�j��|�)�Q��5��o�dsA��(�!���2dN�"�n^��`�!�<�R����<U�u�ʀd�T����wlRA
Bg� ܂��f̾b�=�<��&L�`���d�*>�A�$�ٌ;�V}�`�U�h|����'�ݘӬU�TM��W>c��	��dklqA�`ˡ��*A�Ivu�h��VW؞4��.N�����FU�Jd ����L$�����n�~Xa�/�S��$H==�xK׃�+~':�z7`����)�7�r� �T0#G#��g^���M{�'m�)A�$
�F ���%E�-��'L��q�B�r������>X̙Fl[�%�*d�pμQ���E�c���y���6�(�(�ѣ
�	u��XP��'{�tm��dx�������;$8�W�_)Y\F�Q�go�5� '�
B�m��Z?�N�pQ
#�4��A��	�?T^hh�闤2��1x�/�z�X��U?�%��_4W��8˰bÛ_H��85�F�][5�3/8����I�P��=��ԟ�7�C�[A��H���E�m�I&�n̓�'7^訫矇O�LZQ*�>}DPB��.�uv��/[E�|2�*��H_�l�1�I��f�����3S�*\|pºib֐34�U�{8XʒŊ�BL��W&:E�H!�ǂ�*��EI�J�9����v��(=jPH����Ũe2ʅ2>������)?i֝0kV���!�V�V��bمZ�ܜ�&�\�U���[ �u��i�iN�������T��:,8��3�h�!� 6	���C$����v(�W�WHY��J�>@E`x# +�2�f�A%���
�����9;@X9
$س���3:U�J3V�V����@�<N�r�#�ʠ7vj���">�I �$�U'A/\ݚW'�9+��12͒(Qt��E��[��Ti��APe�,N�·'K�*��A�2� ��6��f�jJ�d]�<3t��q��0hצm��Eϖ�G|Bd��d�h�l�@<ᳰ'©9�� 6�I#oo@�xT��}(����K�`֒,ʆ�ċG ������j�0��FċE.��a���q�t���dH$f�q0I\�'�蘥/�:j0B�9�Ă7�0�D^������VX�K���f ���l��$!E>oX	) �P} a0KF/KZ�����C H�?]ʂ�W,3����&��+��[����U؁`l"P$�#y�}[��K�]j�9h�a�#L���:.^r���L�P�Zq�+A�-�|��#�T4�j���7K��˲跟�Pv��?#<��䜔,9X�`���4T�=��G�I�M��c��q�tHs��,�r���rV��0!��+�Hi.OkL@*o� a��x<*���o�}���	n�ڶ>c�Z	&	�0/����@�5��F�U `��4��"�o3�K+O�M�rlG�B���(OP��$@�5_J��f��#6��hZ�I��D��ˉ�Y�j�q�F�O��!I�t#�\����hi2�Y���8���iR����&'I2��r"�	�[�fi�e�I�|u~�2!�%[��[N���U	�B�$L-X������>��)K�3�r�
Gm�;�����Q�N-sWcX�v�x=���	t|}��ȋoL8��P�7e�a�7GVhK�!��B}�-sp�'���8�D5"�F���]
<�A�%�?CVL���u��C�4:���"���*0�ԥ�5_��	�j̨!�%���|�w��/?�˓{��2��KA4�:jP�B�|��א���)=��S�)X��%��CRJ_�Z�����)uӶMbB�3{.v��P�kk�C��)tѲy1�+D�Z���`�j�c�`�)qR����b�$�3膆
�$2�Ѿ*V!�ĝ�#9n䀥�Ȥ+j��Ł=U{!��ˠA�&l�1d`�AB�	!�'괜{w;dfn�c�G�8R!�d��p���X�X��ꊛF��	>�<��b�}��ԫ�� 4`L���բ|�d��o:�Ox��m�>k���c[�?x&��Qe�s M���X��y�#�3@��P{�|��Y���'�O����	d���&(�S�o�����"_,|�!��	^�Su�B�	Y(� @�h^�G�b�r��ݢH�jر���m9T��ny��9O|��+4d��M3bܮߪH�"O� �ԍQ�>�e��	��|S�;ON� �m��W:���))<O~q����cF�5x�Ȑ'�^=q��'D� �7
�a���Z��	���pp�&y�Qx����#���Βw=(�㦃�W�^�ၮX(J?�#5��#�b  g�G��x7P��$g�6`��@2��sV|x��w�:M���&R�1Õ/P�/��`hӦ.%8Ir%�2���s�d!��˿xB�=��� t�ՙ�m!D�42�C0t0H��M�>���q��~�㇀�'I��ڳI	\x�����=�1��3x��s"�<�O��!&o�=q�����A8�����.Rn�:����w=��h�S��yRe�k��e�q+��/$�u��aQ��HO`ͺ�CL5s�0�|J�"��y�NM���ʦ�h|xҎ��<��O�%z^�h���1j��Y�G	�	�I����e���\�k�p�A�,�!�?i�Eѷ/m�p)(��D����X�<��	:$4uj��2����*c�?of��c�%3씢}dg�m�Uf��;�d���{�<QĂ�(?�� �O��HΦ��I�F&P��Ӂ���	��H���	3l���`�G{�q���'j_xC䉖m��x0' D�=��m��a�7����h'���=��jJ�w�LL���D�&�Lx�J\؞������D����'�-)Y�!�z���g��xh����'��x��ʮrB���D�I�I[h0:�}��R�\ Wc�R�O'�T�2�V)
grDx�E�qF�,��'�epR(ܠ.��c��K�Za�,�&@��$����>Q2�>!��.
\��$�*d�X���_�<1ƀG�f�����ϥeRB�zCo�� y��h�X��Ɉq�E�2bF�z]HQc%m�##j����+h�Y�';�H���Զy�Lx
a�@U��i+�'��(����H:A�AR��ၪOLR�I������ܽkrPTi�N��(�phH��0E�|�a�	�� 	7��#G. ��ꂙ%��uy4
	�u�<̈́�8��R�4.�$A��-�$'|EDx��Įw&|�ge"i]�<��w�E,6z�E+t�O�5��}��"O� a�`R"0����;�<��V��o	2�q2A���S��y��?H�0���E��Y}�AHw��y�!��1�Ys�*!X�r9��y2�Q4�� �EkFaC�y�	��E�����ɟ_�ȹ`q��0>�.��5�(̲$��#z��DH�GۋS�
�j!턪G~�Ѱ�'�
���I�7�S�O0ZM���D*
? %Xfi��� �?}�%�R �z=SХ��
��!��$D� $IΘQ�Aڰ�W�tm�g �"C���I����	�p핧�����2vxH�G.����0�ҹ*&!�䛎{�%��NG�)��۰.�/~,�ڢ[�z��2��;����D�?R"6Ih�&̀/�4��(��| ":~�:��Ԉs�Ւe��2<�d8���iɰ��ȓR�`t�G���Z�3�&�����鉲4������BY�O`�0˰$Z; �.��D��*?�0�
�'���C2�M�|66l�ӫ��?���
�'?�� ���Y��)��U���R��yB@�(_�I�F,�?������>�y2B>�2�E�R� �Z1�^��y�c@�2yJc�k��J��PC��y��̱O"��3���sۨ�� ����y�n�[���!`��0c$\�`���y�̌ޞ�;�n��`-p���'�y�.}�*I�p�*��@]�y¡��TH���ܩ�
�9�ʏ�y�Ģ`��u%!�l�~Ib����y���i�l��8~.a�q�͊�y2h��2 �Q���6m�� �q�ۧ�yb�TnX����ԚcJR��Ce\��y2c��*�$j7��!K�h
s����y2�L�d�P����Sl��r��
�yrʒ�^r�ai�"_4��I��yr��2`,0�*���W-n�!�W��y�M�=D`�ժƅ@>I�*Ԣ��ybϻcʦ�sr�_�F-�����#�y�Q8x\b@�6��c���4�y"�=^�eavb��S���s���yr�M�X%�P,�N� ��A���y��W<tO�u�7���2F	:�y��/qM��MQ:��&� �y�Z�L�T�R�O�VР�!ϕ�y"`A�W4l���'�ډP!`J�y�
�L�Ā�Q�cX�p^��ybGV��Y!���=B0��y�dI�0�x����߂�F÷
�""F��p�l�:���P�'[�;T��z��J�J\tR	�'����mW�T8�W�ɼ'�<��'�H�2[�4	ׁ�3 2<x	�'��1)%.Z	?�,���`\��y�'�\=�t�M�5����%JӿF���'Q�|��� 74d���9k��	�'c���ċA�%��s�N�4l �	�'y�P`0�P��	5�ݦ,�Bݣ�''p����7>��XRCcR�x"ld��'�z-b��TA���1%��'�b1p��F9�Q�flϬ)t����'6�L*��7,@�Rfa#Jz±��'"&��A�֙29������Y��'6tq��P�B�!s��Ї6h�		�'��0����d�G�
5��Љ�''<�@` �p�`��f�H�>_"-�
�'厤;s�����VnX�80d�P�'�h�����S�h�k6|S^4#�'�@�Ƥ��;½��/�&T>��'x`@c���5,(��[�1��@q��� ��yg�,$�@z���R�L �"O�-���<U�����MśPO�{�"O>T�Q.��v�|�(���8�1�"O��遬ن\���#�kP��`��"Ox4b7J�Y�4P3�k&�2�[�"OTA�1�<'�|��H�x��	�g"O��R#.[��y�ef%� (	�"O��"~v�y0�F~MF�"O�xGoۡA9��D�]?'����P"O��x�"��1��)0V�ǥ92�B�"O�,�1a$ c�I+�x��"O���e��<nϔ���"�
e���;�"O|ѐ2a]UU�,�9��t�"O>�фA��ꡢP���^�*p("O���g�(>y�g�0�j�:'"O��a�U�e8�$�ʬ{���b"OP=�-�

v]�ы��K[�	ca"Op�I���S��r!V�nA����"OfT��1f۔5Å`\�[5�5�U"O����-ͣY�� Bb��"#�l!�"O``Y����w_�, ē�`p$g"O����SET��:��T#�m��"O�d(���1#}�$��̸r�"Q��"O.]@�`�	e�����2r�@�=D�(����4�.�XФ�tҔ!�*'D��ۀ��"�xr�k@J�X�)&D��S����4�rH�� �*h����M$D�|�J�\�&x�nۯa�V=Pv�"D��B�6P*� `#���P�&F?D�4�aD�j�0�1rK�7K:�ɰ�8D��p��uA�I����32�Q +D�Xz��>"/N���NF4w�.Kd�.D�����"����+Z�.�ܥ��,D����4(����f���M��G,D�0K�fEb2ֵK�B�(ش����4�I�,Ф��˓VXt�b��q��X6��6db&̈́��RPd%�1+\�b�@"��ބ/ĨMq�ۑ��C�	#G$e�E�D,�TMz�DF0�z��$.~.r)P�{B�I�g����K9OTf�8��y��U�p�$aīJ:,!��� ��DÊS�dx�{��	6|����$�D�h� hU!�Dֿ`���`g"߀;خ��T   >TqO�Lj� ]8���P�q?�	�ӎ��rRPԨ��5D��Sb�
-8l}��G�69!�(p��%D����
$�"�"�w����n9D�D*%�32�B��"m�
�6��.9D�{���xSn	�v�[.Z���)�l,D��J��Ɨbt�ga�K��1�W�*D�xbe��w��D�u�;���S׋*D����*A/��A�B ��F]�@�#D����	�V���a��^p$K'D�j�/1�lx8Ĥ[:�1��#D����$�~�ђCؠ5� h�,D�|P��.�9#w�ֿ�C��<!J� ���H�S�$#�^��R�R�=+ZP�W�
��>�Q��>)rh�$VS���e�8*���Gˏ�"�6i ����O�9@���&5�B�c�ؼa�ؓ�鉌O:��Pvn�*?a`����8B�(��xeX+��V|�e�BݕEH�X�S���&Ӡ)c�oO�p=��Y7R��*�mˁg4BQ�mզ5�@��33�4l:��^����IO�(�eۡ'�R4De5H>���.lTI� �$�c�j��y�NL�Gh�3KZ"��|Ű�~����y���9T�(`��.�t��6GBrJ}	݀��T��.)�zt�2Mi� ؑ��D'�p>fKZ�s]�T:�G��]V�+�+�C���IϻS���y�aݜB<�	9��9�g��w����]1O��;wm���R��&��2�%i3�I�V.�8qa��c9��� ��<rj�$k7��3W� �У�a_�CŪ�0r�$W?r��2lZ��$9P��.c��Ap��'���d���j�^-A��
J�<@Ehƛ.v�8����"4 �͢���34Df��`���*^^,C��<J��=BA`n�>|H��֬m��Jc��x�[!"O LZR�P�5Ѡ�,�- ڔE���WnX-����FԒ1@ MXV�ʦi�M�[�؉X6x�a��$��U&e�!�qW��ˤg6�O.2�E�lE�2M��3�
ы���_~�ڗdO���|9Ѯ��?���Ǐ=��e�4AٷSm�Ј���{̓o�jܲ��G�	� ɶ�O�4�-Fz�`�1�����D�d�eX�]3ZK|Q�ƿ-���q�]0|�Â�ի0 �ن� Y���"�Gl�X���I;��"O2]�h���!�'���	�r%�ゞ9)ڒ�st ��z�vWW���pC˔M	l9;��~��Z�G n�fdh�́�+ P�q�
?D�`(�� pmΕQ�Z�x�a��K�j  ��T�1�,�J��(��`*���ON�W�B�d�(`��Gz�E�厏� ��5��ߠ@>��G�9�O>��A�A$9.x��V7]�f4:&�I�2�*|	�� ]>�uҟ'2�E)ǦҷP[� ��N=,f58�}2�;pA�)��ɟ�pK"[?��D|2��(��Ň��ΕA`��]#l�S%P
Zp��!`��?4���J	����9P���G�'p>=���P�2�$ �2��x�'l��֢�C���)�I�'�><��Lm�0�,��y�O,�m��d�-5\�؈�h�&[����'��yY�� i�����8~<;����� ��8O�s察�o2~��'BܵO���{썒EK^-j��f���2���&|�|�#�M�O� mۢ���.V�����d�f.v�ZQb���Hh� [Q��bq8o$�I"kG�>���zr,�(`�d��/��]1���B��p8�e� 9�
�%�>�|�����i�v��+߉0�R!���*%e�P;m�/@p|9�Y'[��˓A? ���L�$lp!�BY�c\�dYt��ʧf���H�?]�4��MW�o�޽�ȓF�5�$��oRQ&��$I$"�i��I3°�t.�3���I֡	HEȟ'�D��W�H�W������

���'uD��I� U��	Y��ۍ�(�8��>�D[�_��ppu�٠H�Q���⌇��q�@D!^�hr
7\O<�'�N���ԻA���"C�H�;/�`���=G�R Y@�rTa2�<� c(J=|�슔���O`l��+ q�����TN�-��	s)�{�Di�0��y$ބr�ҙ��B�P%!�B
��Č ?������+����*�"'��T�v�C;�B�	�iX,��^�(�xBs�L�k�B�I	]72aY�'�d�v@��._�ZC䉚����@�>�Z,�%eڍj�C�I#Ir�d��H �FH&�y֯�t{>����9
i���!Y�����%6_�i��Ꜣ">!�$ݖNMȴ���ӊ"���C��F�"2���R��yj#|֍�#Q
@@��i��/���x��J�<1PhZ�FY���g��-u�0a�����<)%ێy~���<E�$#VE�F 
�d��Me,]!�#к�y�h�"_���`\�@���&G�������H)�w�'z�HZ�i�"3Nd��ۯc%n���b���G�>�X@9r#��AΈ�YrBۖ%c�L�ȓC��8v�ՌH;ry� 
�S�2MD|��C���ډ��	g� K���?5v�U��!�@ Pԛg�[�|W�DsBÇ?�!�dE:0	�Y�R`N�%��,J��gN!�$�+"�UY�"�$5�^A���),>!��O�'$*���l��5�
�tH�%)-!�$Ѻt?Ji��C�9��D�&�P�0�!��<T��#���D"�q��hޯV!�d! �Jt!��#��'H�PQ!��P1f��������̔=����&D��j�ř2޴Y��D�W���"!�%D�T@�,	�)q-�z֐�X� 6D��bEǙn�xi '�L_�$���
3,O�ђ�N[̓a�&ɠ�hPp�6�O�f6�i�ȓ#a�lr�%�,U0���H[@ԕ'�@��)��ا�ONBe�"N��.-B`�?0���x�'����]�p��x�$�A�x��}�CF7���]���%��b�#`�t�2�Q]�!�Ģ;��Y&
^jܻ�fY��CK�\<� |Pq�[�:�F�����*p��%1!�'�V�ˎ{"�+<�(�&�B�iD�qPđ��y�HZ>?�Ё��&x2(��C�yR�FuHI��$ t�Hh����y�eɒJ��Ⱡ�#o��i#�R#�y���
X�ZesfKZ e��Ms���y"�B�n�2!�A�ψ�bՁ�+�y"M	w�P]����5	�Y�����>�G>>'�Iba�_�E�@�r�	6@��Ȇ+Y4!�6�t�T(�p.�ݱ���&(���`�G_2Xj����|��2E��{I�K�戃y�!�PSR�8a �P�H����Boy��JK#+���K��s� 0��&W�C\!�q��+E��'�B��"`��q���-؃i�T���O$���F�l�lSϓ<��]ȃ玫sDL�{eJX�~݇�I�n��C��G����M:k��(;�A"�@0�'�z��U�!��T &�Q��|�Y�'�$���˸g�����3�`b�'�.�k��G�T%�Y Iͮ%h��
�'�	��	^x�,ȓa��#/rY*
�'p���l��c ��L	�&� �'��u
C���hwL����=�@��	�'Z�t�v���~�%�/j@�};	�'(x�j��F��:i�bO�J��j�'�.lbu���;c�}j�Ë�r��
�'��EÇ �,gh����� �	�'%~��-�G�^\���3��H	�'������7H1��GMq,�{�'��lB�$Q�'��i"'���'���8�G>UvHyDO��
8vyQ�'��d$WaD�8��ً�����'��}j7��#x�>��*��tr�0��'֝�5�۪I�M�aꙚo�j�{�'�Y`A��� ����n�@ɇ�z���B�Q>k��p�+�1\��T��#J�U�1�A�;�FY�ǭJd����u\3[P2���0� 
��Єȓ\��ɓ="@08q�>w�F���h�l!�7adM�X钾r0���ȓH��`x��D�����jN91�f���H���Y C���!��;']��ȓ?�=��lɣ\��!) �9H!�x��6z[�Z�hN��F�ڼK1:4��p���T�P&i��!�Sj��M����ȓ.fŻ
5gٴq�t��p�P�ȓeY�!�T'|e�YUDě;>nX�ȓl������S ��d3"E1PE���[+�`��㌬0�H�`�M��1�1�ȓ[���Yӣ[�{Z6��0�;?���ȓ:b|��䈑&d܀aDŜ,�*U�ȓyؔ�����'>�"�;$�]1����ȓi26�A���> ��K�!M�{��ԇȓz�����\�g2�	cc��E���H�VЩ�̨�,0b�j���ȓn�#Ɣ�`��=���E�����t}k"A/�� �ˈ�-{����j,�Yw	 4�u��!D�GL�`��Ӿd���h��$���REB�m�!��?qw j�B��,~Dd�7k�B�!�Ǐ\��}A%�@�Z �)�ȅfj!�$H)yp4�q,� P�:�BGJ:�!�$"w	t��爒�b��m1e�X�!�P�,�FUXsn��h[aKG[�,I!��9q�l�b�3Fp�[�e�4�!�� Hl*�=R1b�т�f�<�C�"O�;E/Oo |��C,	z�,��"O6Xs�j�jc��Bf�Ši���"O���jTq�"x#���/t9�|0�"O�tӖ�|�����;��
�"O��Q�@�$v����f�v�c6"O�Á�Ө<�i�¤�!N,��"O��B�F-	)�=;%��EG6A¦"O��5+�A0Р��э,;��*�"Ot�VZ�6�C��.u[S"O$u�@�������Dn���F"O��j#e�+&L�6�O"T�踪"O�Qf���Cm�=�!۷_�ѹ"OpU�D*^s�� �T��-Ht�R�"O	�g]�T�bH��ơ77�[�"OX��G����s��`) �²"OpY�dES�l(�b�?."�0U"O�h�wd��N��7�*u`:�"O�1[��('J5s��Bpn���"O:s%h�c�D$�d��{P���r"O,<{�EO$@ Mz����=��b "O�Q���Y�u�\C�2x:nx��"O89�Rʜ3&�5Ue��.M�"O4�[��6pr*�T�	�(t!�"O@@"gN8��y�5�T�HB"O�]0 �H�W�С:����a�����"O�X�%`f���=\�(���"O�X0�$څ[�R�:�G\>H�vLq�"O栣�G�41�2�&�4:�\�"O�����څ
9DT�0����!�Ě�X��T[�0aWvU�f�
�!��7~LZ	��+�,W%��J8<[!�SL��AN�VU@�K</P!�?J��h��MލKĤ��rJ��!�B$m�  ,�L��@�`照q�!�P0#�:a�-�>~��r�E0 !��
h�ʈ�T�~����G�l!�S	�4REZ�Y!��Mg!�DI�@̼䡶舤|�^��E%�$Ik!��~��Q� AC&	Ӥ�]!�#��\���M1
 �fC�	L!�D��$�j��]XĲ��%�\�6-!�$�B�\5)AB9�~�"��ʇH!�Ӎm�n��͜JH�q҄ޟ@+!�G�+����)Ý3`�d�,!�dݠbށ�(�E8�CBCE�#Z!��زIT�AegS�J�&I���0P��NU(�%�oD6�Kb�G.ij0����� �s��$SG���$�E�ȓ�r� a (p	�5���NY�ȓ�J��	Q�m}���M�7�4U�ȓuuF �FIO�\G\)
�o\�'��a��n_���	b�L�MY�i��܅�'n<S�υ*��k��S�u$����l�Z����K% #�1�� �;% HІȓmV�Pt�P�@a����I�ȓK�	J��_+E���aKЖg'�0��Vb��G!>1T���>0Nh �ȓ~��9�ҋ�,@��!I��E�ȓ" R!J�ʌ%L��"��� ɇ�m2�( A,<4��\,��T^���FN�f̂`"�e�E��ȓ��5R6���ы�E�z �ń�����y��&�P|6%��S�? $4������)v���];��bG"Oz8@F�)J�h�Dͨ:}�!��"O�sĊ�mҰd2�2v`1�"O�S�j�Y���h����Ҏ���'���3R'Ӿ�uS��/̨ɪ0M9D��jA-R���Q�Q���P���!�b3D��xtAј1��{@+ƼR����A�2D��d��5�=��"Ȱx�^5Jgn-D��0�"ݙ'���ʷƨI�Hi*�*D�@����p���qe�"\�.�)D�lS��%䤙ʁ�b�ʷJ%D�dۂf�(�
�@�OZ*'rؚc�&D��+�B�9��K��9XW�P s�.D�,s��=8ݲA��R�z���j%B7D���M_1k��B3bV&^tb�4D���w�б)I>��qc2(o1D��lD'�J`��? I�%��_�<Ys�'0
f�J􀅾&) $�b��ȓyD�d��?�T�1�	�D�ҕ�ȓ<T�3�֋UZPYb�!R<�
}�ȓu�L����Z`��"Ԅ��$\��ȓV���Hp(B/�q�3��=\4v���24I�q�IlM��/�X�ȓA��b!�
'U4�1�AET=��Cbe	'a�L�� -nV]�ȓ�za�%f�� ڵK�)��|��8��e�\d��On�:D���T�ލ�ȓC�����������S�Q>|�X��+p*\BկB���X"��>}�R\��c�,Hw�L�t"Y`ň�`�@�ʓ}evm�f@^D�@��#���:C�I  ����S&Jv>��%$I�C�	�p�lT����@��-�WA�,��C�	`�q�-��E���vf�>x&B�ɖm)nMp5HΜP~��ұ*ӿt�C��3��)�*t�NIS/���B䉭8�0\i��]�(�
U���-� B�	!>����.�z� ��ID�>�
B䉪'���#�ԡm�����ˁ� %�B�I-/z����	�:6�I���8e��B䉱"��ͩ1�X��m��&ǔ��B�I����:��U+e�M�#�� Q��B�ɽ�R�o�V��t2��N�~K�C�����▫�	R�ܴ��/��*�C�.� ��%,	�^�t!%B�RC�	%Z�: S�3�n(���"4UxC�I�w�K�/�5H�8��-�� ��B�	�i��p���\;8L���6	Y+\�C�	G�(KP甑4.�Aa≃+��C䉺C/�y��ŏ�Da|C�f��}<vB�ɐj��)�1K�5k<1@�/��-B�B�"n�	�f��/����	�0|B�;-�(�%��32�C�ņ�0��B�	�;>�"��ŉW��Y��$��B��, �)�홛E����V�)Y�B䉭?Y��	P瑜-��hQ�ݙw��C�ɔ/��I"c���#��f`݌L��B�I7�2�`��] �9ae,)G�*C�I8<��v� 
!�m;'Z�:B����}����N���`Ù��C�I#qyS`�j�Ы�bZ�ZU�C�ɯXT�Wm�~��Ybv�� C�ɘ;]�r�G�6Nֈ1s!H�3��B䉥ZM@A��+���c"��0�B�)� �vQ0>�3��^�G�>��f"Oԋ���"�9���șK�6�Z�"O����mԖw�D���
o~�U@�"O�аq��!"1sv�<f^�5��"OL�+GËA��Ke,�O�W"O:Pzu����p3,�-���"OҘ��퓾|1@Aa�
ӹm��ś�"OL3�'�Y~�`��_�yz��{Q"O��H�`�1z歑$�g��!"O쵢�@+du��*M�U�q��"O�%�#�Ֆ`dF%�O����"O쐁���I���q� �4o���p�"O~l��Ŕ�8�p��nO�>L�x"O,���K̻e4��rnD*V��Q"Ol,�a&ʗeP�L)�l^��>�!"O���5��lj|,S�K�q���"O��Q�!I��е��"�"ORUÖ��(n�2Ɂa�C
*�:�C"O�=�T�H�x�F��Dd=�$t��"O:�� �R�o�����	B�Ne�t"O~�S��
,/�&	�3ⅵ����w"O���V�A�4|EA޻d����f"O&%A&lA~w^,��O]��t ��"O֠�� W�`L�M ���*J<*��2"O����&� .�q �%#&�]�"O�!��M�#T8~)aD���,��Ա""OP���uv źF��&,Jr"O�%[�y��&V�b�"O�iAk?J̜��^q5��aƞQ�<�6�۠S����aMF��ye�B��/gˆm��*�i�d�"��*K�DB�I�rrDܳP�X�'6Y�G��!F��C�I/�|�`��O�pN*!)&�B C0�C�	�dt|��!$�H#e�ц��"{�C��,EQ|RRLʦa-Jh��"R;{sTB�ɮ`*<Qy���/�HP h�!"��B�I�@�
̻�/8=�T	�b͜~�BB�I�m�Q�T!^+D�IPi
P :B�E��9��j%v���_�\7hB�I�=4�C''��j4��9���0:B�I�C89఍�Li���5LZ�vjjC�I�vT^�Т�W��ܥb��V�� B�	C��e�aR3��љ�MV���C䉶>�|�y�o$j��@�O$C�I�i��e5K�(Eh�O�;��B�	y��싷"Β)p���M��7��B��1b2t�2��*lL�����M|B��< �r�;�m��vp9d.�bVB�I�I�A@c�f��;�̒-ĔC�	8y=0� Bb�&������
}&B䉚k��$HZ�y$��
���?�`B��I�>���J	?����'�@�%��C�I=!�,�
�!P����#��`��C�ɦ+�#ҥ	G8�ȴ-�ʹC�	�>%����N�H�X%���N���C�	�m�� ��2��&PCI�C䉳s����!i-,��`X��+�(C�ɷ;���3h�Z����ڰvN`C�I,�61ԏ��4���X��p;>C�ɖxt��J�)J�k'���X �>B�	�R0�,`�O�F
�$�N՝e�C䉢Bt�Sq��(�p[��GG��C�I1C6���i�_�\ k�>dvC� ¬EXu�8T�`�u脰�C�)� l]�T�� HjU��ᓋK��9�"O
M83f�5D`� S��٥(���T"O�%A��W�`=�X`�݁v�Z�"O
�K�E�k�,@�
L��BY "O�LC�Cӝg��!�L°τ���"O�$��똏pjae�],���R"Ox8�I��2�V��tע}J+�@r�<+�+LvTIrP$�>���7��r�<9⃔�c���ؔ �zl����B�<!�o
��|	ئ��_�`��X�<��B���e#�$��t�D��x�<�c�Hp�|劶[�4�y�Q�Cr�<��fY��&8z�h�Z�f Ѳ��m�<At�8JP� �W����&?T��b��B+v��Be���h�T�3D������S�91�J5[�ʼ�!�1D�0C�M�����Ɲ$L�T`�*.D�� ���;� ���*V>WєpE�+D���MߣRk ���G�.�|���O4D�� 1�7
�P�J��޸d�
y�=D� �b̂)l|%:�꘿Dh�� �I<D�D����	f8!�� 4�V�9D� �f�#N�l��1A�
n� 4�@e%D�1��ުg�2={vHT�m� \�C D��!�P1V�zia��7��平�?D� ���W�/Q�$���6Q��Ѓ��=D���ů�*���3@��W|���n:D��+t���U�B��/D!�֌9D�xH�*ڕPH1u�[�����-D�ZwD2=,��f�ʯ/R��'& D����m%W�:�c�I ,,���4L0D�(*�텥?�򽠲��U����0D�!F�-��J��EKt�z1�+D��s��B�C2��Sk���`�k��*D��6
C�ri�}6�S>T)r�`�%D���DΛQ��E#��о  ��g�'D�p����\g�y	�.�l�W�#D� f]
�j�m}Єٶ'!D�D��#�M���s�'	�,�Ve�%�$D�x3��ȰH�H�1@I ��! �"D��JgB�Q0�0'��p
(��a,?D�\#@H _�"��E�̭	��Rb D�[��/��- �]8��u�7J"��<�w!�x;r��փ_�=�b��c+�B�<���<^�(+LT�o�4�)�j�s�<نmU	H"i����#x��91��o�<)T,��p,�i6,�*4�l����g�<id_#`�)��� @���HHD{�<�,O�s\$��1��I���� ��P�<iD�D�>v�0��狛A�V@#�n�N�<����0���I�O����9s	H�<	�AǫL��X�2f�)2nM
t`�G�<��AA�3�q��E�L�lhc�\�<�!V2P�d�F���)�L��a��V�<��H�K�P󵩛f�z�"�W�<�#G�6AiX9	С��de�"eTV�<)����j�Vn�G}�X�S��N�<��gN�	�4 E�s؎���eI�<qTGd�V��c�XݐQ�ƌ}�<�4�uj����b߆� A�Cw�<�#^�Sޥ�q�ЦaJ��ԤOX�<A�b��f�"�VND7_~]R*M[�<��JN�2���r��!O�1xT-�P�<�0�]B��Q��)9�ڬ"�'P�<� ̱���
�+S ���,]#y��,�3"O>0�dLсG;@3�O�^� �A"O`�d��,���D��ܸy "O-�6)�F�(؁���$���U"O=��.{W2� Vʆ���,�w"O�$�pl�&ϔ�TdP�r��,�v"OHar򌒢����F6�<�"Ot�k�H����y�+D5��l�g"O,�(�HЮ�F(S�M�a�Ѕ��"O.�x����"��<m
&D��"O¤څ�ѽ��AH�L	�S����"O"���P�C� d`#I�D�ȥ�0"Ov�C؂!}B� D�Ѭ@u�$"OhhY&��?�(x�`��3�<z�"Oj  S&��6��a�׋2���
1"O�h(Cʺ*��Ő���,at�Y�"O���RL�"EO�L���50T����"O(M���:����P�ͪgO0�@�"Obb��C�qw��� M�Wk�$y�"O��Xg!Gp�|�9#��>K,�1A"O*�����C�:���J�1m;��"O���4��I������#���W"OF0�g/΀�$�dO:+�x�q�"O���b���3bh�I�+o�|0%"O����?���a�`�!��)�V"Oly懽x�`P9��Z9��ҵ"O��saG���.�+l��`"O��`��ϲ4�l,9����[��	H�"O��p� �jB@����BK�"m�!�Dگ||d�����Т L�!���n�Ǣ�T�����kM)a�!�
7�Q�rCF�jg��0�A�a!�ļf`:�;Q!�YZb��C̝B5!�T )⍣w�R7^���(X'!��@8ֲ<�d�U�$?��a�N۽!��V!�8��Ņ�4>9�9)0+	�"!��U�4��P��#����#Z��!��!#������<ePv��P�$j}!�d�q�¹�)rN�\V��"@y!��,d����%SM��a�螴 y!�$��t���0q�NL����fV�o\!�$M9FbI�F��]�Y���S�<AfRE��5��"��6�ԥ���LJ�<1Ҡ��5�vm�	%Hh|�� E�<�0 �/\����Q�ًl�r8�d�A�<IäHǶ�[�Fؾx�䛦+W�<�$OD�'E�]*7��5�h�ӲF�l�<i�(��>ܒ ��� �9'
��w#e�<Qn^�*� �X�څ ���:T���g�M��b!��߁Q���%l)D�D���2H̘D\%/Q��(D���[���͓O�>E��B3D�x�G��⠬��I<��B�+6D�0r�F�8n�>(��Ŧm����D�3D���&�U�bG 5�v�G���p��1D��1ͳf�&(�u���,��|�H0D�t�!��(A꒤�9"F���$.D�营!?{\�Á@F26�l��*D�����^��	��b�P�����X�<��̩flXcpZ��l*r
�X�<�BO�M|4x���3�1"��GW�<��e�!�ޤˁ���,,DT��FQ�<	�"�&��dP�@�:lb�x��,�L�<�g�=O�Isg��;B�<��C��m�<� �Xb��G�8� ���.\�r(��xr�'���U3[B`4�#�g��x�'&,x�S�V.Ԩ���9	��8ڮO����`\� �AlH�~Kj��2�H>��6�>�M�"~n?N��邬�.0n<�{'�+�.C�Ɍ1/
�uL�-&�r�@���C��=0#6�Išò6���@��@"O�����-*������'�H�R"O��hTb�p~蘂%щN�ܸ�"O����L��fF���ĕ8 ۴���"Oek�.<`Gt����~�:Xq%"O^�ˇ�לT�x5�۠YXp� 7"O�ɓ�덝R��L���\�1OP��"O��FX/+&L"�X0ZX��"O�3�e7����� ��D�(��6"O��Qt%\�zO�š��B�Pй�"O�8c�a*&:��R��HH����0"O>��s�M3
@)�e�f4d!��"OZ �`kA<nT���,|��"O�R�l�aNy��!ӂ0x��ڳ"Oj%�Zh�r�V82e��F�Qb!�ۢi����# Q:��@��f�k�!�$�(k�6��稛9i�<��tO"C!��#;�v4�Sb�/e����O~I��'n�"� � ��x &@�$l2��'�X�`��(	���%L
3- i�	�'z$@�$.|�`� �� �(���	�'W.H����,0疥h�k�&r0$)�'@f���X :0�P� ?L��a	�'˜q�#�3
�
��2��u�|R�'ުI��AтFʦ��b��>pTΉ�
�'�\�P��%dUb+Q!���I	�'	��y�C]�Z�LX�Q��X�X���'�ٚ�Q�H:�1�K5L~R�B�'��,����:4���DMD��X��'�V�zgg��"����r��&0\L5�
�'
�%��ㄲ]�Ps�!�$^{N-�
�'�9I�8�R�x!RWQ��1
�'|~��<u<��9�hXO�
�)
�'�8��7H�-#����oǾM���2	�'�:e,`|$�Z!.ԭG��z�'��Y��\�m8t�×���:U*�0�'Ƽ!�3%��)sPݩ�Mט{���R�'A�w R�EqP�	�Ʈr�n
�'�P��G�.:^({ӊ��n�Z� �'�Șs$�.l�0�2�ȸR��u��'霨0�7��0.�;� ��'���s�Ͷ�t��J���9A�';:x�5���
$�ŬҩD8V]�'2�Ч�]�|,�/��B�~0��'~`E˴f $�������'���kԍ���LB�ƕr�6E��'��SF��o�L��U͐^N��[�'��D�Ш�-�I�a��VFޝ��'tvX�W'W:G*]P!�{�Xp�'�5.U'BA�УX�>��=��.�c�<���1ly��r2�O�u�P�15_�<!��B"��S�܋��\1I�o�<a�"x*u݆!.�s�/R�<Q&`�-�0������h�*}k��c�<��$�	C.�A����4(�\ġ�ND�<9���'L9� Y Ƴ=(�	RC�u�<Y��V/#� �Bɑ-"�ʙ��}�<�7�n������e����a�<� ���ɵRh^t8È	�>n��w"OB�8������	�<���c"O�5�c�;C��H�CЀ�C6"O
ݒ�Ոx�r��g&8���v"O�`邃~X�Ks�Kg��a:�"O*��֠"j���:$(�"O�!ᑋϤn}
�fLZ�G
ʘh�"O:�1�A@�N)��j�	F�M��: "O*y@�X�԰略�l��@"O؈��R�����_���e"O
h1�
�<U�F�s!��;Q"y��"O���ǒ_��kť܊SJ����*O����h�*eDD����<��
�'}6��𧟼�~9��. t��	�'^����43�t���^��bղ�'�a �c�zW8��C�̦��'�
�;ì�	��$	t�M6���R�'R�� ��A�5��!�NL?Pb*�'�J	�GJsv�0� ��KZ�a*
�'��Z�M'o��Q ��4=�^��	�'K<�J�m�� �8X��!�:8*f�C�'~ݐL����9��م7�؁��'�Y�C�ɏW�`��F
*&4A�'�B��e��%�rm��h�(����'�x��>_��A�ٽj6��'���
PM�0d`�e�x��x�'|���0g�>h�5k���$U��'>ą�7d4�ԭ�ħ9/����'�Xi�CB�I7�k!��&���*�'�J�;�ƍ:^�TU�q �� ����g�~(�r��"J��9�aɗ
fH�ȓh�f��whХ1��@�&d�rA���ȓ��!&���v/��l�+F��̅�V��H����� ^*'@��7`�Z����� �*�-�7��M�ȓ�ֹ��/Y�r��P�3�ɞ?^�E��i�6|H���q]�hY�*@�Tݞ��aM4�rr��L�T!鄨�!y�نȓ�2LpW�H+*�z���B��
��ȓE�H����!!�ҁ��C8N��ȓ�<IR� 2H0�,h�h���"O(�b�F�3P����ʅ���"A"O�Er"�Y!D}�)P�K$|����`"O�x���_��J� 
#w�`4�b"O�A�&�8y�̙�W�M:)��u�"O�`)��/R�0��ꎔn�Ґ�1"O�����$�J��zѰ�J�"O�"�f���q(ȾZ���"O����e�� �%Ɏ�v���"O$Mۃ���R�N;��C���"OD��N]	]@�гh�.	��9x�"Odع��5^�p#IȻK~z�+E"O�Ւgꋙ"�UcG	�CM�p��"OFH�ъ�V� I�/�EQ�<H�"O`�H��\�:v}�.�]bD�Ѕ"O�xC* �5AV��ä ��s7"O:I���:N�t��4�2<GЄ�g"O���1Oߓs���veؿs(�! "O�a�eE!\yH�#'(ޡA�"O褒�ʂF�
9@� �N�<�q"O~���,O��D�ҏ�d�Y6"O��&"�!*x �e��W���"O�\b��З$4��.H�P1!"O�����Ș{�Tm���M�V�x�"O� L�0��;S��ݑ��֍-�z��E"O2Ԫ��� �t��sO�*Ǹ��"O�,�c�wD�ha3��I�"Of���B��p�`��#���x%""ON�x��+h ,��W�N9n�0�R"O^t"�� �S�.����'0��a�7"O^Ԃ�l��ZD��f&ϱ^�0 #"O��HL]+t��`2Dԧf���J�"Oؙu�Y�b�VE�T��""O  �	sޚ�ۑo�9�Q�5"O���/��CB~��G�X��x�"O��`u)�*x�|p�,�Zǂ1�"OZ��*z�*()`K�(#��(Y�"O�)�K�W� pDQ+C��j�"O� Y�o��]\��
��,A�`���"OJ�	�����`b܉#��р�"O��ӱ�[����oK&>��y�4"O������Q�4��{���"Od���͒=XHɢ"$AFt��"O�����,R��q��"�a)�"O�b�I�X��t���Ќ���"O��B �>(>�#-��8�z�"O�А�ƥK*�Q��� �2�B"O|����+P����,��'���ʢ"O¸�e�S��{B�2N�v�I�"OTAPr�L�truH ��AY�"O&$�s��00�!�e5}�m`C"O�p����>c%��AjжoA���"O��+���2\�u�5J�"�m��"O�=�f���JXp
�>jْ�)"O�=� $p�T��B�J�M�"O*���ԲU�X���a�H�ٓ"O���p��gjl��f�P%l֤�`"OJ�y��	3�A�v�.P�D�9#"O^5P��U�%Bq�waƠ@�\�H2"O�`S��J�-�.L�C��P�X���"O��0d�7���*�/�35Z��g"O���ׅa@�KN.H�xw"O��0���a� yd�A�"O$0����&�UFݾW�&��"O�Tc�lE t���e�P�65c�"Ob�2�C/�a�NǚC��Q�"Ol1з��$���$K�-e�t�8 "On4)TW�9�����.4�,�"OZ�����d�N(�Pd**6���"O. ����=e���C@�L�x'�H�R"O�ҥ�"`�RQ���4C^�@"O�dh�IľU
Y2%��'�x "O̩�wa�Q?�y�n�#G\�ڰ"O���N,T?a���.QZ)t����	@��<[�%T�9��ʟ��P-���:D�p�S+�`X�#�@[�LAKW�:D���R�C7n�1(�Q=92�"D��ʶោ}��mB����V��2է%D��A0$��f}p�x�GK!���TO>D��h4�T�Z�,�Rb�Rkr%j��:D�Ġ�M�)n��kӎ�vmX��=D���# �/Nl�7��=�0e��&�Iz���x���9���E�&����G�?D����d�� Qd�@��vT��Ao3D�������6��2�(�<,�;`4D� q@J<Q���iF���>G�)9�'���D�|c�-r��KB����
�'s`���Ȅ,AB\ё��!9Gδ���� ı���Z�¢�+v4U���<a��4�p��2�Շx�v�Q�`��Smf#ǘ�8���JN�b���?J�*�cD�� '�B�S��]Y���KB`�P�)2pC�	�d���9$����|�b�i�sOhC�	.?��q��-a��@���;@BC�ɀ@=�a��|5H�iRjX�fY�C�	{��]"D �
s�����?�,O:�=�L�pxe�X:4�b��e�rR�͓��?�%���[�Ni����;7�2Y�6"�T�<Qa!��\G��B�K�5#���-LS�<��!�������= }#YI�<�2͜)u���bG��fB�qC|�<a�%�L�<�C$�1l�^�B�p�<�ǥ_Q�ə���.��=�`�';�yd�oX�	1
֮j�Y�dKgt��Slt A�pe�-.!�aZ3�!�$�����c S�^�ʍs�R2�Py�Ȏv�>t3rAI�M��4��:�0?�)O~���A��Vp^T��6=L.���(�S��y�%6aY�����5,
Ή-W�֍�ȓy��E�8~����P`K n�ȓ��lI�I!Z�� ����\pD��ȓ �Z����K�y5Z�o2
�� �ȓ"��d:�j���U"B�\.Du�ȓl��ȗ��*{��p�`ʕ���}��D�t`���,"��S�/�&&$B��cH��g�[�.��"�;(�C�Ɂ5d���-�>��!��B�-�B�I���5�� �	 NC��hO>�*�%�"�4�`b�N�\�i�N'D��&�ײo��y�- �D��#e$D��C�O�d.X8V���C�\��� (D��@���5�z�Z�Λ�c�Py5�>��T�j��A.ç(��� �aI4,G$M��S4̼XۂQ2p�pR)�.>f���hO?�a�Q���1[���if�6?9��������EL	(5�9Җ�^��@!�"O6�k �\'bfD�X5O��4��"O��@�a�3T�91�͉#{��#"OZ�AEB0�*�#�A0 ���1"O�01�	�Pn�P���wLy04"O"X�3$	�ZXv�9 c·T<-�eN/�S��y����/@��e9�p�V����'�ўb>ѫ��/]T��R&-tI" M;D�8���,f��7'�>���DLx�<��� 2��7�:(���g�I�<�fZ[	>�b�,��� I�J�C�<	(ۚdv���vlX�9�G�A�<�уY�p�=h��;ԁSQ����'F�𙟌�r+�>zO�yI�#T�ՓA�1D�Pq��t�ق'���tҜ�j��2D��{��Wj!�1�PEb=FK1/D�0�$H
o����+���0��,D� ���s0�8�R�fE$�<D�8��!;�$đ��[$D!���:D�\�⦆�k�BS��.{/���`�:D� ��oK�P6@m��2@��1�7LOl�H�E�+� �P����^�yB�s�Dx��mL�'�� ���y�V
T!��c ,H�P�U��y�L@2Kд$���8�d�y��)�'x ���TTH�c�"w��A�����m��QP���8��Ї<tܕ�P"O� ��;V�ɢS�l0�Ԁ�r����"O�`��!�>O���-˖$?2��1"O��V/��f.0�g�M���u"O~��(i�N���k�n�P�Cs"Or���VuD$�!Lڏ^��yI��<�I>E��'Ī�q����r�"��e1X��O���;�)§#���Ȥk< �&m����Td�}��Zz욤I�/J��
���n�J�ȓ<� �cK\��Ij���/V���Q��H��*TD��!���"2=��/,@�sRaQS�e�1�XNK ��ȓ3,><3�O�D�iY����jH��z�^8
7h��+(��1�߄<ܪ܄ȓ9&���%E�!�F�G� ������?ɡE�{�����J[<{Ƶ����L�<!sbߔw6Y���ґ}D��Yfg^�<i3�֊mx@���(R���'n�X�<!���JhI0ύ'�hݩAfZY�<ɐ�G?Qvn���#��:O���wc�Q�<)UA�l#�̣�bƙL�\���K�<�q�Ñ�#�mH�#�h�:A��A<�#TPR�@�N�pȐ��P"T���a��E;֧C�*��İt���^��Q�ȓ\5(�3oҼX[�@(j_�+k���ȓ�
\����.��ˀ���-�~��ȓ.�Zc!�]-�j�%���jU��-.�)�$"�:TvjQ�q�>
��Dx��'��p�e�̘�af��l��	9�Or1QA�ֿs��!tiϥj) ��"O���'P D�vp�`(r�9A"OU��[�R0��N�bE��n��yr�H���<�H�'4Vl��!Y��y�B܄w�ܔ3���1��]� ,��y�gZ�j�Jy���-rs1钧�'��{��_�����H;��@�֩�ykJ�Qٶ���J(2�H���ψ�y�"�b�d��"��,'�B-���ד�yb ̳z|�S�"0!J�*U���yb���$�q[pFX^Sb�
D�"�y�*�:"b�23�)P*�T�����yR���
��ȫ�k؂�F�@S�+�ybh�n��Ʉ�Z�8 
\��yrH�R̐D���|DK����x��'�Z�&̞� 3X؛�Bܳ/���k�'�t�[�o�W�
yx�@Ι,3LtC�'q���o�a��fhL;6��|��'6�LP ��G=Ȱ�7�Q�_�����'��Z�_�+^��N@�l��,��'��cDG�)~0X��̫x�*�B�'��x��) Ii:����o3�5�㓙�D�OdM��L,h����o�#I� �(�"O6��B?玘KWnS%H��Y&"O��f'A w�U��=J	$1��"O��ddH�#��M f���P��Q�D:�S�'qۂ��g�Yj"��Z�ߣvv��(����ێ@鴄�צ�!�4��(>8�ᖩ^�/=4b����
XD��d����օ�W.��y�l� ��%�ȓM�qz�+C&s(&�1C
��Ț��hZ�8'	7ib����4���Y�I5���X��V�&kf�pmi��B�5���Eb�qVfX{�@��..B�I%�X������U�4䂤�S�T�B�ɀU�%��&�4_E<M���
B�)� �lb6����&=��)��|�VU`�"O�UI�O�3�1S�g��X�j�q"Oj@+5��n�f(#A,;W���'e�'�h��fաUU��ۆÅ �ȅ��y��'��y!T?U}����a�v��-3�yR%�`U�#�I�jR���yb�Ɛ:F�墴��
3<`T$F�.��'U�{2�ea��CFB%c^�(BL��y2�ثN�@*w-�.N.E�&A	�yb)@�wՒ���DoG�2�d�7�0<���$ڼ3P��t`X�Fh|��ef�
��X��	#:���a��I��P�	��C�	n�r��̉�-�h����T48ϸC��/����`O+6 ���$_���t��`Tˏ�5!�	�kN�p���c�6D�l�AΟ���=C���ht+ֆ4D��[�'��9���1�L�a���#4D��RǬþ_�ȡ�RN�sS��邤>D�TxB�S���Q,UeX���6�!D���b-ϭ{�r��-
o�ԅ���,D��gd�9Q��`��(�1ҙ�G+?�	�c}��QFG[�U��)fڵx���ȓ.[�xR��Z�#��I;0��2\�ل�$�~�Ȏ�j���o�kM� �ȓ��e�#�D;bS����`=��@�}0c��*!v��*� J�h��ȓt��p	��̑I��l�F*S�%�x�ȓDF"��E�ŚV$b�����1o�����V�9��ū	����f�-f��e�ȓfL!��*�*lb�C�'�&x�(H��PE�� �X%iFY�7J�()���ȓ]�ء�q��>)^��n۫t�1�ȓ#�@]BWc�S��|p�X$J+�Y��P!��c�B�4�� h�B�����g��ܐF/�S38@cb�U<���.��)�?�=�!G�(g�]�ȓK� QD�"J��)���$B:���ȓR�±S��(w�Q�w��"�����z���`��/0uQ���ܗN����ȓ/w� 	@�ɮ_�x�hu r���ȓ\\) rkN�7�@�yЭ� D��a��+�4�,JV�ɰ�N1xP]���!u�߿n`�\�2��de$p�ȓ�n�# �����,��ȓ?�l�BmD�G:N��4���N��ȓH�J�sPM
>TEBSE�'�L�ȓ8�6d{�jS�B���&���-0���E����%�2WVDaG�C32̆ȓM��Q�q�Ӆ:�0Q��2K;�\��m�(�	��\*y�l;$@-s(����[
�4j�*f��c���c/���{FŚ�'`��g'ی/�̈́���P;�F�#�Y���_1��1��_�����	�kBj�z��Ϊ`Յ�j�����5)X���n�k[��ȓ?�:h
�mR�&�:�J��W)u޾$Γ�hO?5�N�D��xh��ъs
�W�<D�h����$ȵ΃� ۶�"P�-D�8 g'L=<���9��#��Q1�,D����Z�m+�)��˫� �1
*D� ˓g��~"����*J���ɥL$D���T�[VPs��05�|��S�.D��`s�N�l�����͐I�E���^�����D�5���b�Wk�( vl�S�!�� �\�d��#(.T�f;�n1Z�"O:��A$�z���#�����1�����i��+��ȁ�+r
 Y��:,!�d���${e� rD��)��Í
!�Ă;2��ӵΗ&_b~apN�!�Ç�<a�0��Mi�|�4��6v���:�S�O&�+��Pdt��tIH<0OFLi�'�TsՋY�b�*��S�C�zt�0[�'��M�#�3&N ��u[ab�y�)�S2:��jP�@(|=���"iqnB䉶PgEX���B/@�s �V8u4B�	0�2U�2�4�lř�(��M��C������S��aȎQ��A�-nx�B!D�pG✃�0u��K���0` ��?D�dIC��,aJ��5Ɩ�H�:�x�+ D��R�ϑl+V�;em�{D�@2�=�hO�� ������-R��ԦͿw��C�ɑI����E+(ČM	�Ÿ�nC�I0BĒ� � l9�U��"f� C��d�,a�Q��B�!P	ґp��C�I~��0YS�Z�
�p:���*+&�B��^-���㝉e�r�h��[YnC�	�y����5�"��e��c[�C�	?H~8�p�O��V-�I�B�WE�C��.n� %�ׇ 9�6$�$³PЬC��)QF,H����3������x�RC䉀�Х�&�� �5yӰ�hC�	�f8lD���C�v��4���Pj�6C�	�`�|� �(�6$Dp2M�,xyC�	'�.��܂E��y㵏L�XS�B�Ʌv}�Ȋ�G1�9J�h޼E6�B�	[���@��6rua2�	
DJ�B�ɲ=N�A@)P��TM�p�/}xTC�ɧ���X"/�m+\���h�C�	�F�l(�ʔW���N T��C�	�N������"iL}�'���"O��@��[��ؗ�E�e�V82B"O�A�2H�Д�2hQ�kz���"O�y���σN��]{�'��X�ۂ"Op�Tb�/M�(��Egޖ��0"OL����ШY���x3�0���4"O䬉b�'6�b��Y \X�i�"O��� �G�%��!��c�.S�D"O4�q��A�z�mA�a�S�<�y��	K�O�����&�hh�7�O!?���x�<��o�&"�Ȩ�ӆ����d�"
l�<������2�-P:��3�L�<I&�ҫ��0ذ�n��1��KN�<�2�ގ	5�<�Q�Չ\A%ӷ�M�<���	�%��hH�&�Sx��b)�t�<�qJ�9Zθ`�2���J��@��Rv�<s�H<���K�O+���lh�<A��K?�y���>xu��3���`�<qp&�}� p��'�(��-D��pr	��^XXb�B�z ��ǧ �hO���Y1�W2a�ҼW@��C�I,;�n�����(�){�$R�C�3`���`�9�x3AŶJ̐C�Q_
9��/�"l�d`�J�G8~C�	����$��{z%�Zhq�a4D��p��9܍!d@�2�����@$D����+�ISR���#S�}i�Up��"D�4;0����qvmO�U�Q�G�3D���C[�?���aSd�9?V:��2D�� ���P4A�hԒ@R�>��y��"O��S�Q��`�ϗ�r4i1"O�i� �˿b v��1��R�t1@�"O��%IH(pR�@�)�<j~�P"O�kc�E�J��@��CI\̰!"O�h���yEr8�Vg؏ g!!�"OzͰ���)��|S�/_�}e@�@�"O� !&�A ̒��F�0�'�'x�Br��*l N�j�+��"�J	�'�䢵��fp+5���^�c�'q�l�� ��k��z�n���(;�'����&�ɿ)i8p��-� �n�I�'g�d��5&R�J$�@�@�$a	�'[,e	� G-\Δ�bS��3�xIX	�'&���J�6�B�[�)�%x/�-:	��?�*OƵ��f�>4?t ƃ�ێ�p�"O�ӵۜn�0�#š��V,�f"O h��JI�N$݋¡�!M�8���"O��x󤆥�z��b	4M�A	"O���*A�X(:��� 1
��g"O��C@^e��8�"��*(B5�`"OLH���'p��d� �2�*=�S�'!�O4H�t�m
`�8Яx��M� �!�Ą�G#F� ���	B�ءRub;|�!�$A0����L91��H��j '�!�I��I��dʼg��(
�jV�Uc!��3�^9���@�0�gQ[O!�DBG�V��s'�a9��P���pK!���]Z�d��� @3Z���Mx!�dG4�l��&��a0А!�l��&�!�$Vv�:��@�
��x��#{�!��ɾ=P�pr��U%��1��+t{!��
p���S0%�-v�VU�(�wd!�D�9*2�� #�4����^51u!��0`�����3�2�z�%�:i�!��ٓ+�pU��E-��#2E�/a|B�|2A��q��Y�.\���(R��T �y�̓0>Fb���Y�MUP-�T��yRo�+n!r�%ƽt�l�b��-�y��T*.�a�Z�:�(�CU,�y���:�f�y���3J��zR ו�y2���rv�"2N�����L��yB��TAܼJS� �}��-��� ��0?�.O"�a &��^R�AP��C�1��Y1"OR��ꙣ_-���"���ꩰU"OĐ��MC�1�d�Shښt�za��"O�Ȓ�� -��*�F��u��Dє"O8������\������1��H��"O,E١n���$@�I�1��q0�"O�@�ЭW9 �@��&���rV�'l�'�D-B��Dk&��0�&_1
 �'��H �<R��P�%�5+(�Y�'����3ʈW��rE%�(s�1�'dS��N\�If��) $x��
�'��t�ǝ �r���ƹt϶�`
�'�L�J6._�^�^�BO�=}}�|3
�'�JM0�V�x���jBGB�_��	���D͂3̺m��RMB���3!�d؂,�����C�M�����)�"A!�d݄J�ȱ�P���0~HA�H³=<!�1�����$$�98��^)-)!�$ܭ��p���z�C��̙X�!�O�|^���l܅_�2t����2$�!�Č=I#أXh)9 �q"i�O6�� *!�1kښ'b�`G�JE8¨�6"O0���I��H� �o zJp� "O��)2NC��bM�, 0��[�"Of�rK	K9��,�.9�M1��'��	`y��O�H��j�l����{ �!�y��iV�\(�?
��kE��5�y�,ʧ:Kr�JJH9ze�p����ybM�""B�Є�1~���3iѝ�yN=h���ON�i�t����_�y��	�R�6��tk��Z�4 @3i��y��&X(�pF�*� =s�%S��y��_F�Ru�d�\62؅���y2K�nԊ��5.A#�7�߹
_!�$��<���7�G7(Bp��K؇\!򤗳m��I�&̅4$�aj�=\M�C��@h��0���}�h����5��B�	<C�H�z����/,�S%�IX <C�ɳJ�h20��}���R�ݒ1�*C�I�x�^ċAE�+v��&��U�LB�	�J��D��曙!5d��U�E�h�B�ɖD	�XA��cN]�ª��(U�B��\Q�1Qsj��@>��yA!ڎG��D���{�	Oe��+;��n7D�Hw����c5���'�T� 3
6D����D�B�P9@qi\��͐2o0D�|
C#@GH�����,�I E0D�D!���L�h�A�(^4��Z��.D���� �#e�6�)cn�<ޠh���'D�P�e��Q���8r.��G��	7�0��<I�V�F�}�j��$i{���]�<�p��.S���Ch�S�$1�T��@�<y���(?�$9��
` ���@C�Q�<�0�SQM��9�P�y�LH�G�N�<���ƍ��G�=�����d�r�<����*2���� �))��Tz5�Ip�<��*�l��T�ī\)��X�ǌSm̓��=��j#]����VX�$���Mf�<	^��Ts0/�8R��� �U�I:b���ɂi��H�֋�3Y"�`��@�B�	�(��]ATM^ �D��ȓ5<�B�	1}� 㐀X�m�Xʂc^�3R^C�I %YJ��T�!�����-u��B�	�͸�˜aC>�͕�~�c����	�vAْ'*1zt��ţӔH������?E�d�'rb�`Eh�'/�A����Dﴉ��'�Z|4���$cnX�D�8;\X���O�u��
�+4�Ĩ�*�+~u��B%"O������xhLI�)v�4��t"O����G��i֠,*$(�cj���"O������"`r��Ǩ��V^&�k�"O4�(VE�`"�Lʥ���f�騀��TE{����i�.`���\>��a׫�$S��2��hO\���E� jB���Z�V��T;C"O�9��ND�&$���i��m��{""O�h2���W`s�\�9q,<*U"O�1��ȑ�bk���� �A���0w"Oڌ��H^�2�"Ȥ�؏~�1G"OX��㒁d$����I �:O��%A�
�C�Qt�TT�&/�!2���%���IM��:.�h�e�Ŏ%%P���W3reC�ɔj8��s��˖K(�hG�T�9x�B�	�c9�Y���^���L{Q�ǖǢC�I%p)�0���ʑk��A����Pg�C�ɬa7<�
��]B�U��"�=�!�� �Q(�d��U?���Xg��D��"O|�ؔ@E��� ���S��&�Xr�'��'�t�:&LmS,�*v%� p����'،���¾ @1�¡�d�pɛ�'`���ǀ��3�лr͜	d��'c 8B�/��V�ⱂ���P�[�'d��1*z�ʊ>,����'��p�A-L[	@pC�2�Υ�'l	� Q(:H�GÃ?o��Q���%�'03�=Ss��}� ҧåVPF`*O��O?�	�U
b0@��8q�2�� `�0B䉾n��\z$��Rݨ%
�yI�B��u�#tA��
�z}+F�޸NM�B�I�	
��5�P�4J�0��I��B�	�"+l�@��_�.�#h��?�B�I/�t�QǍP{IB!��	�B��䓎hO�D�7�N�0�(^���
S4]�!�DJ�}ʵ򱢝qג〉�<,�!�޼ba ���J���iQ3Ԁo$!�$�����Q-��!��{���2!�ĝ�}�z=��C�?H�ޘ#V�l�!�֛:6&Yq�fS�@�BŘb��2D1O��=�|j5烩d����(ΞE�P;'�[O���=y�'_���\gK�7O��0<���DU/�4X`V,��HE �p2k;}�!�d%oJ|Kr�N>��P
�?U!�Ѥ]v��b�!G� �U�D�A�!�d'$��:G*L�������ے�!����,�c�0{c@�q�Æ
5!��I%�u�#V5NQę ��/	a~�S�|@��X9<�C���>kS�����>D���]�P���)$2ٲT{��9D���A�̳b|��S&���l�jt�+D�pss`@2�FZC�z����o�o�����䉉�>���D+JҝA'��]@a~�V���1 �<���%�ma���do$D��Ȕ�Y�w�ba��œ �ƽ�c #D�l�E�/�T���6`�1��6����8z�����ـmv�y�#$�soNC�	��|���LL(�]����1�B䉪c�0�'L�7�z���1\����hO>�r��Y͐��Ǘ�hlR4�EF&D�|��ʜ"h�1�c�@,'�ԒW�)D�|�1�[�o�aS�l�t��貵�,D�H	1cP�M=��c��LH���My��'��D �	��Lx�k�""��'��u�R%��4��;�n�	..�[�'u�y�ܽc8�,ʡ�@�"��D��'����T~��x�! $Jf����9� ��D(�	���eP�����-:˘A��"<D�� "e�#y�p���B/o2����;�d���5O4�3WL��.� &�ԅrTx���>	U{�̤�f-w?
�JG��j�<Y�-�$��D��t��T�U��i�<��ह��������V-�I�<vm�1w��$C%��.��@�}~��)�')4<��q��D刧��hk2��<���ap�,4j�BE\=SD�ȅ�X�II�F��bj�K�e"ǴO=�B䉴%�x��	*3�@p	�톀ZbB�I[�69@1c+\�:��L%F�vB�Ɍ²TS��E�b4d�ޒ.�VB䉣E>�ؓ3�J�Xd�@ڹs�@�q������s�끝X���KA�
ΈI�++���<E���� �T¤i��L�$kw�	%$�Jt� "Ovͪ��6DD���9A����"O�	�t(�O���V ��T[j��"O��$V$U�2�AB�2I�2�"Oj�ё8�x���;6v	G"O�i3I�y��B�n	:h'^��Ā<�S��yR�N
If~8b���3hJ���$	�0=	����/ h�挍�X��p��}��'C�e�'�2���w����
C�?�� �S��y�C� �	2-��9G0�3P�.�y"�2V�&,q�Q�[��dH����y��VF��!뙴^H8��F�	3�y�(�*L�p��u(Z/mg$Ɋ6���y�e_q8)Za )g����ֆW�y��C�U�D���m�]��\��fҍ�Oz��DU��^�B�ً8d���2�!�DO�Y��U�=���技�'4!�Y�4���a�/�j.�$�EDP5(!��ֹ�B��mM~�\����Q d!���*]�V����_.}���ɱi^�!�EOa^����S-c�.]�B\>X�!�" 
����&RI���s�v�!�$ʚ/��� �40.p�oՉB�!� 7"�������C��:N�7iZ!�8L5��Q�AO}� 9Wl�5}�!���	Ipr=x*�$I�4�[/!�ŻF�XhӇJϕk��y�`�s�!�,��͛|WV��A��%Y!�D^G�]ˆ`�q>���.J.<S!�$J7Z��m�t�K�IBX�k�+�D!򄉪m�z1p �\�),�+љ !��枈CBa�8 ���ēoy!�$�� <���
�.D��,��s!�J$1�\����(PQ�7r!�SJf8��܀p��C� �!�d��!i����͜<x�𑓢�Z�K!�$G)Vڐ��s�V���r+\r�!�dI<%;����B�$r�����T��!�d�2J.U�$H@�ffl3���M�!�d��8�&x����/tN ) p.Ðj�a|2�|r�� +�Fљ�m�:#��T�v�T�y�-U*��TJ�%#	N11���0>	���ф8҆H�ק��q����B�ƕJ:�=E��' �Q��*L�\>�����#���"	�'n"�� �\�7,ư��CX*G�
�'�b�j�ǝ�@�&�
�h0v��	�'^����A3�h-�t��!n~D`	�'7��CF�?z)��
�aG�f��tH	�'��"�cΎ%
� ��׾4 �	���h�(��W��zm�!��#7�!�$��S-��
UΨI���YH!�(A���s���L|�*�Z;&!�� 5h��!�%ddE�%:.z�!���(SU��a �2]�04��pp!�D �o�e:,@
fJN$��7qX!�D�`Ӛ���ʅ�A5Tq�0�K<P�!���OFX3@Ą.o]e�Q�;N+h���5��Nx�$;b+�+pR@�`a)�(|2`�%D�`�Í*�6� w���,r"�0D��y�ĳS�f-C6��=��@�ģ-D�d�q�G�Oj����@�j�lp��,D��qc��N�v����o�n��q()D���OW#;π�Rw�<yd���(%D�Dѷ���-���P_� �k�A6D�� �|¦)��'@fYy���+���Z�"On�B�ݨE �а&ŏ�Te���"O(��6
�6��5��xP�!B�"O~p�VgU=M{�՚A-�B!	�"O�83uf��$�4t)�o(�-s�"OH�;!�C�I��q�ɉ�}�|t��"O�A�,JP|�j��l�i2"Oʍ�r 3}��2�\?m���06"ODxrpL�:p)����OX;��L*�"O�Ѐ̆;"�^�T/��$�er�"OZ�eoW�J o5<��"O�ݣ��7�$Q��N��,Ш��"Oh�i�Z�(�KE���_�h�`U"OƝ����A�p�� c�-z��93�"O
m�tE[�%�vD�TO���j,��"O�%kЎ�5'�N�07oֲT��"O	��B�`Ii�$� ?�	��"O�Hj�h�����x�B���z���"O(�P��*o<����PoPd"O�i#�D�i=�6��>9ի�"O�����O�~��`)v�Y�^�\�V"O�(�G3#��q��G c�ii�"O���)�<A���ćM&'�,m �"O��pl�r��qK�%���@P�"O���lR��V)�G$��.s�X�"O��)b�l" ԩs%P!)W(ՉP"O�t��>%F��R%܎��4R�"O���I�xdb'T��p1v"O��0���.�f�hT��8�h�"ODi ��3m����ǰG���"O�8�CD�v���c6�ؘ8Ժtڲ"OF5�$��)��A�oP�/��X��"O����I )	���퓼Z�x�@"O��'�M;���!����%_�A�P"O�q䨍�_�|�(#�d@L���"OV��B^B!R�xS,��NzR"O��k�ʒ�H �U��<Zm�� �"Ob��F������&�k�!Ӆ"Ox�#�ϋ�N���#��S�@�|�RE"O��!#�3j�+ץ]�c�|x�t"Ob��/	�0ƌ��7�S�&-c0*O�P'��($�#&�9N4���'�,T�S���Dp�FF�rb�
�'v��ph�R)VI�զ�m��M��'�1���#6���ի:T�,��'0^]��
�nbX4��BK�t �'yb�5(Ib6��t�Al�'a|0&�� ']>�Q��?��@�'�|�:���A�0Q'���I�N�B�'\|.��=z��@]̒pce��y���1�r��`b��@���d��)�y£��=%�L�'�ζ2�pّ��Ǆ�y2$�5l�0�2�OWq|d��R��y�mә!�<�۶�]�K�R���!G��y��/8�A8�KOGx�4⇠S�yBC�z�4Ц�R�=����b��y��4g��ܲD�ު8&��Ä�Ǝ�y��z�L��`! �6P���Ѧ�yb,'�|R�k�A�|���V��ybl�gǆ�J�j���nX���˱�y�+ƾHʜ;&�U-���S����y"&F�熸�W�
�j�90�L���y��P�+��|����5N, ��
]7�yr�;~�j��4"R�0&}y����y
� �:q�O�h�%��׾|�z�c�"O�D���
:�Hs �I�B��"O��C�ã+OD��v��k��p#�"OT��S���7�VБr�:[���Z�"O$�+���}|p���۹1���S"Oj�n��h�Ћ �)�"�*"O�u)�L�?/n��!A��|��0{�"OҀ�dY���UA��\�)��K�<��MX@����!�́Ɔ[D�<�a��5��N�D�i1/PG�<A��I :5� �a+�J��B��B�<��)P#(P���)�;<|F< �b�z�<i�	��:��y5Hմ#&8зH�y�<ɱgч!P����O�w=�K7\p�<�,�0@�K bͶT }+1��a�<�f�Q�B��e�/���C�_�<)� 0j����]��Rԛ���t�<����u�ƥu��B焐C�hSp�<�r�@3�hɃGH�<(S���d�g�<YÇ �$�ґ�Fȟ'�`�����a�<��az�� ���^�:��T�<�R�Uu�t}h!��1"�B�� O{�<)QjKr=,xh�������Dz�<�QF�R�8�a]w���ը�v�<q���{O�|2�-X�P�4%FW�<I�&�]Ɯ�D!өav:�j��V�<I2,�!Z25���>�vl��(�J�<ɖ�ͳ��ɺ&�����qY�<�
�n��]!#�[郎	vo�b�<!�n�>8�r0��X
����Q�Z�<���p��0ء��|Z� ����U�<)��� �B��FC� �~)�V�R�<��K�5[O�5��iR�kr�͠s��M�<�D��)��Iɇ�2nVYh���N�<�������U�V��/`2��g�_M�<!2N�}�ܡ���GL:�
��P�<�+�<�.8�ЌC!j�� EgEt�<Q�� �?�6Qs�fM�	�c@�K�<Q��]yAQ �!BP��E�<��O}xqx���B��Y� ,~�<��FW>v�4��V,�T�nQ*�
|�<�����nO��0GC�6�����#Is�<)�iP�hM��x�4"L<@BWn�<q�Y	���á�&B�R�`eO^i�<��C��LX0�C��r�%��a�<�S� =^��! '3pGt(D�S�<Y`杠 w6�� �;V�*u1 �j�<��aψ^�@M���̴Uܔju�k�<�p���/f���\�1z����P�<�Ӎ�[lQ�D�<1�� �O�<I@Ň �����%�a�'\H�<I��Ս �ɡ��9P�T��A�<Q�B©2�$�ڷ�,�j�I�@{�<a��9_��p�D,I��U�!�x�<� kʾL���r!F����iV'�|�<a�Aƒ<?�i�E�p~�@���N|�<�ph���T�����MU�4��O|�<!�@Bq���AnƀX�-�6��w�<�vN�m��u���M?u�Ep�/�s�<9B�
+��q�!�I�%H��p�X�<�4'Բ+� �c*�'��<�F��^�<��ԕ	���3W#^)�e�v�F�<�W�˙�|8����a�c�UD�<iP�/2��9r��� !d���K�<� ���h[,b��va[���4"O���ᇖH� �hB �?u�f�"O��JbNԶg����ԎN�mn�"Op�*F���!����m��񢤚�"O��"�]���pB�S�H8��"O��#qJ�^��5� aВ�l���"O@�!
^� �``
7oҘ��� C"O+ nܽc\�H�B���3"OH�a�I� d��m��&���"O�t� `'n�nY@+��hn"P��"O<�H��� z��t'��<a��D"O�a�f��'d�#7�/9T��"O�R�t��� rK� NDQJ�"O  �BE��{���>J���1"O�(�[|fm�B,<.H|�B"OB�z-A�}�reԏ$\�9+�"O�=�@�/):(uۗ�ɅFA�	�F"Op��R��"1�ڡA@�/΁Y�"OP0��A�H����@�܆>!4�Ɂ"Op@�p��	Y��7O@7<��u"O�����ϭm��Xr��4�d��"O�]����(<�C�C� l�|��"O-)�KD;L����#Λ5����"O�tCŬ5�Xhq�6���"O�#U%F�r�Ip�'�8�2�s�"O0�$�
P0`∏����	�"O�i�E�<0�^ɵgB�\٘,y1"O,����-�^�8�N�B��!�"O��s����}҅�-_�<�۷"O�����_�-̚�#���V�l���"O��#�Bct���&�}\b�+"O�%ZB	|H���D��@s&"OXɐ��֯.-�1aj�8�5"OX�R1�.y"T�2�MR����"OxI���ݟrr�!C���X��́e"O�`�#]�f��zӃQ�C9F��6"O68ADٞ>�ܒt��
�l��f"On�	GiR��&w�Pc"O���������tۑ��I<P�ȓ;��d��Ov��Uӎ��cb�ȓ	@⽱���9J�V�jʁ'"a�ȓe�Jꂡ�%k��T2"O
�B^��ȓ-�T�h�!���A�b�6U�Ї�B���t+X�:lT���ӵ{QH���1R t�3l�Gܰ�𪁮2l�=��Uq,)��M�}�jJa�J'�� ��UK���2#�C�`��� t���NX�V��Bp���'Q	V��ȓUD(سp�'�e�6|bf}�ȓt�X�4lA3m� ��HF����ȓh��4�T��=��4�P	[�~r���ȓT���&�n3"��֣*�)�ȓ25��Q�������B�N��RŅ�$E�� G	H�4���1N˗J�T��F>yڇ,F�*ϸq�0��':���CV$:!�UB�褫4�֥ �i��S�lq �%C8(d�
ş2�8��ȓ����K��Xw�?`��]2�k5D� 8C�Q�u����o�F1���/D��`6�0WF�=��R;.:w"+D�d�eFʝ
ʄ����*H(����d'D��K鉙r0h�+�7����#D�,�'H�m`�Iդ� ��I�cn7D�d��'I��mܛ'i"Q���4D�� \K`L�'�BqaBM�
�r�rt"O~����+�Rq�P?p[>�X7"O��娎��"��J�nq�	��"ON$b�@\���fj��BU( �Q"O@�������͐`��	 =���"O8��3_&s�:1�P�C�;*v���"O��"�n�?F�`�;`ϕTl���"O��7���=r�ER��
g�Tt��"O����ؤ!�BP�SOύ��;�"O�E��o�g����OӇ���B3"O�Sūד-��a��̒���u"OP�rC��?R�x)!���*$4$@"O���A!��|���#! ��n�-ڣ"O�P��C�t�b�ˀY�m�b�*�"O�a�쀌�b��2e�?)X%"O��1bٿi�b�C���w3��a$"O�'��Q{��!�e!���"O���֩ûrJ�IQ�(��S�"O\���n\�1�D�h����B�@@(�"O��95��(6�X(��8G��"O���@��ܮl �k�6e:0V"O���i�#2�
� �K�~7f�P�"O@01S�ҝA���ڕ/�,fͲS�,�S�����m,C��9G%x�\C�	)7㠨F'	�z0L2 �:	d�<�	˓mc�a��"6L�-�6'�6`����3����kT3($A����,��P�ȓ
oڰ8�G�/T��!�`۬I�|�ȓs�҅�M�J��đ@�
�H���#�������cnl�P�j��m�<�U�/�S�'nQ  ��ןd��0��O�KJR@�ȓ\���G�;he�E�"pEy��'0
ec��ښx�P���H�*��x
�'�&��`�d���`M8*'P�Z	�'m<��D;����G^�8�T���'>���aKɛx�&4�u��/��D�'�N����<
��a5�P.v��:�'�@�'N�+x�� P�ÉiiH���'���hVeC/�(
Q��"��Q�'ڴ���(8h����l�8	�'�0���� 
��:dǍy�T����D)<O�)rvG��Zv�6ȁ˂k�,n!�$��}kE�6C_����6e!��?J�U��C�2�j��C��SY!򄃦z�`�HDV�n�6��D�*E!���B�@�/�2U�n|�0.ȑ 
!�D�	Q�0�2��B�������,.�!�DD�~����N���O_2�!�dǃ[�T���KL�I��8�S���t&!�$�<&��ks܋%C�u�u.܇M�!�dB7r�Q�d��+Y^T� �O�Eh!�DI����@�+ة<h�)�W�֚QQ!�dZ8sy�(�*3]Mµg��X6!��T��PXi �Ae���U@$��ȓ���T+W�NǂD� �[k}�q��|��Yh! ��F&&}3��ڱx�X��VN� �Ն 5<��h���{�"u��'d�Pg@E/~r�� ��17�M	�'D���'�-C�b�0�"��}% 5��'��]Ӧ��;f�0�ҏ5o�d���'G�Ļ�C�{0�)iG!�
�4y�'~ၠd*@����V����6u��'��<s��R�:V�t
��1y�z���'h�UI��߆D����%D�(9��� � �T��r'��9��[G#h<y�"O�� Pi�u�##L+�}c"O.<�E��#0@����!	(����"O����(͠K��QIB��93����"O���w��m᠅��6��`J�*O��� �K�6 ��MP5]�ڔ��'�m�0oP2��y����X�0�
�'@v��P%�M�Õ�P@!�
�'
�H���[�D�R|���:w�|�;	�'0�q���B�2X���#�v�h��'����t�(=6�B�����`1�
�'04��BO
�t�#D.J�o�.e�'�(�@uc�:l0�����6m�΄1�'�T���Y9 �p#c���n��p�
�'>j%�
ĝS�ܓ��F�c��
�'hĄ�1��(@k�=;��_�^�x�'�j}�S��n�=��Z���'�r�����_<0B0��{��(�'c�4��݃[j��B�R�b�d8��'�pt����7N���6!�Z�r�H�'`�85�zl��f�Y�B�[
�'�^�u�͠-q�p�YC�D��	�'%(���C�<c�~�{R���L����'(6�
A�[������0�X��'[�Ғ��S�\��gX&j���'�"��	C��Q`#Ƅj��#�'�bL�lЌ~�����%ex����'�
A�����,�C�NX�8 	�'��<���X2w��Yӳ�R�V�"Dz�'��	�+�}n>A3Vl�GpL4h�'�.�ig�A�V ���U-��<.����'è�QG_�8_���f :ˬ�
�'Ԝ=i��X,%b虊���wa�M�'Ȏ��a.�?� ��V�l�r��'ؒ�ȅ��v��AJC'�#i,>i0�'ª�1�`H�Un<P�[�N��'�4qȶ�{�@3v+�C�\�
�'������\Xc5l�:
�'�l�hq��Mqp\�e&[3��iY	�'�N�cW�ٺ6���;U�V�-r�ġ	�'�Ld2 '׊QS�)�QcW�=DD$��'J8x�1��o�yPJ����HG�<�A�_�c�,�e��`����7 �Y�<���I�C@)yU'	�h8�SA�M�<�����`�	 %%��!P�hEF�<ar�_�1�r$��nB*AG"�9�F�<����.����MD��q��[i�<��BA�8IP��V͘���0��h�a�<Id��v��At�L���8��]�<�2� D@ϖ5n�T0��H�U�<�U+�u̞0�FĖ쮀����h�<it
,l���0o�r�n�b�/AZ�<i�g_3�J�2 ��7ᖀZ"J�X�<�G(A�l����-Y>dRz��+�{�<�ˌ!&La�g�:=�`:0(�K�<�� �C�D�t,K�6Ț�)u��G�<Q��C2;��qI@�0�j@��J�<!�E��3�-��:�jVD�<�a�׈Y�� �@�����I�ah�<��F�lY��A�l�{���e�<�7���@X��FO�$�Zei�{�<�mp&MbF��Ym�m����L�<��m�9Ԭӧl��V�f!�&A�~�<�B�P��t�dK���@$�e�<� l����J�4z`к�\+�����"O��ԭ���	��	)���p�"OV�	�c�'F �W��h�h�"O�=q���?��`�y�F���"O�Q$��:,lHė�;�����"O�|X����a"!�aT++��-�g"OX�bDʄ87݀�(�"Y
�Ԁ"Oty�o�P��Dܙ�p�R"O��P�	Ү�C� ��N�~MX�"O�TP: _�J�ZM�K�bv!��On�2|3�$�o�X�����bh!�$B�0@B�%��~��!�6ğ�kV!��ϗ/���C�#�C�Dq01`4!�DK�{�TA���E��J���AY�"!��u�$daˈ;Ĉy�qjԻV!�d\�t��3�o��?Ӗѹt(Է�!�Dϱ]P~mڥ��*����#��
'!��&[R�z�J؆`!DU�!K�1!�,C�t]q��^
B�w�O�H�!�I�h��M�꒯5�l�q�ճ�!�$�:y��d�X�wʮ�Y�`û|�!���)�����!:� =PD/ӯo�!�d�� ⒜*!�@���I�	�M!��.�Z4���͓Dd�܂p���'�!�d�&L3�E�
���>	2��΂g�!��W����a�	�9��d�c��I�!򤊧pE
Ic�iñe��%�w��6�!�R�Xmf�hQ�@�'I���#Ȯ2U!��AD�q�k�W(p����A!��9�F\)��hK���!�"P'!�dH-8P4���fi`���7!��YR5�v�T�;Sʰ�S�^�!�d
�E������0s>�y�/
�!򄇟O���� �Lɮ��Q�]e�!��$i�lM�!B����m+�l�I�!�䄦�� $+�5c��ݠtb�8ag!�dπK�(��k�H,Fd����~]!�F�E'rep㉩;�8���`��\!����\�1T慴�4� ⯞�I�!�$I@�|��0��W���"R��,!��*���q��ݠt����ia!�Dؙ<cD!QQ�ֵWf��MV�jL!�$C�"��)BTe�(4PqyC5M-!�D�o^����
4f4 P8aAҎsvў��;�ʈ�EA"4[Z������C�I�J�����5��ٙ�'�)2���+�I�p|�H˖E��}�s�G�fKB�	�x��xI�Q$Va��#�҈��b�E{J|2����'��`���_�L�&DO�<���]�A�y��+�d��Y���L�<9Q(� y�zQ��2��	q�^�<q�ŦQ.�]K`�>/�]q@"OW�<��#rD]C#�%)5jx���V�<���]������'%ͺ1�Ii�<!� Y����˗�؟P�����@���<%>y��ۓ-J�P�f�L�۲�9�-#D��a!�v~|
C��n2�إ�9ړ�0<�QG�0=}X� #�t$�䀥�U~�'�?a��[�N\�$�gU�LKo<D�����{	nq�F풿 H�D��$��@��ڸ'��aҴk�.XfI3G��>!l�q	�'.Α8Wb
�u��WK�|J�'*f(�P`��#?���!L�'\�,����)�d)�f�������N�	RbS��y
� �)��P"#`���%��)6#����x��)�S�Bm,�І�<�0�t�܃S7�B�	/Q�伺�+�;Oq�a"n_3]� B�IEsvp:��^��>9J�B�X�C�ɟR�ޭɅ�ʥc70� �g^�,<B�ɗX%�|9`�@YJuY���*CJB�I4q`:�
�҇7.�Ȕ�5l�TC�	<r���FF�� A�88�<���y��)�&�A̽�f�	�V�L�vF3D�`B�Gf���UE���5D��b�
�&��-�3��<��*5D�|k�cǙv��9b�8E>�!�M2}b�)�> ��4�����Sx�r��t�N�;����Oְ�6�˻R||��V���Fl�%���$7lO�� Ao�5�r4�JڈoUB�q6�O���I�/	~�yJ�	_*�!�&�,!��mt\���j�?��蛳Gۀe!�Ą;4�"9�4ț.���$�*	 !�ą�-�⩣b�ˍo�h��iB'�!�O���a)Di��&(��o�!�䂿a썢�`F�]am��W�&�!��p�Fh�(O3$��ʆ��>,@!�d��yo~S�LM��ԁ��	&�U�ȓ�`���̉M��1���hq�ȓz��PЪ4��(��m�%vɇ�\��l�lپo��hb	H(�(�� �h:���[,�[�� $�Y��kI���`mܐQ�9K��ۤlR���Pֺ8�̅!D|b!�gE�L@��Ɠ_*t�.V�6���j�͟9$6�J
�'~I���=�H�g�!'�
�'}4��F$Wl"@C��!��l�	�'�:q��I�p�r��Q �4=�l�1�}Ӓ7�1���<E��N��p��|+�aKC�� j�Q�<��_�ȱ�P�P1$��f-�S�<�C%X�"�ry&X�O�����Lċ!�$�2���#���<iJ��	�wu(����'k�����ָ.q|�+rڜ;�`��'��E(�*vֺY񁆏64���C�}"�*�
��ѱ��� i�Fԋ�<dPB�I�6����EфK.2�A*!�"b�F{��d��7z�뇁C$R�I�SH�~��'��L�q+�(ò	��N�6.�p��M����i>�&�@�c�X����{�bӫ&Ѐ��E7D��	O�wc�Q��ăh�t�0�I}��3��=K^��U��g���a"��0| ��00T^��耿s��P���AܓE���D^�O8�SulݧM�n�R�	2#�B�>IO���'%�$$LM�n�;6Ks	x%���xR��:�c�m��UJb��f��$�yri�,W��Ь~xv�1�Q!�y"
�f�t�1eB� t+� ��i���y�����>���`�p�� ����y�AϚ}�:��a��:�F�B�Eڑ�y�B��ly�i�"^�h�H�ْ��y2Ƌ�t��e`$�Sh��Tqeh�y�^V����#
�̕f	�y��E Zve���w�8�b����p<���D.~�@ ؄	Љ�����Ư����Ps.|�`�ťq�L��S	R�q6�d��&f]['�Z*	+F�BH�+B�,qD|b��rw��S�"��
��I��C�I
zX�|Y�O9K&��7��0�C�I7ph@��P�Z�5�e��2��C�)� NYPc�Rf��t��A�f8�S"O��0b(:G�\	d�Y�
|��kq"OXsĥ�;w�a�f$�[y"= �"O �`ņ!����%�� 4���"OH��G^(NA�� U�.y�$�'ֲ��I����'K9b�ZH�F�&���A-8Q�#�Ϥx�h�b#�*)BJ����k?Q���Iv*�w�H�^ܼ�ғ��l�<�f+�3&԰�$�,k8�S��_�'DQ?��6e�'w	\�2���4� z��)D���gHJ@~Tv��4��$£f'D���1ɞ(��i2*P�+c��r�O&����>�C���O(��+�3�$���"D����*�:bƂ�x�AV/��� "D�d�'�Q�uȢ}-���P��}���p?	b� [� Z#�MK�|a���Pa�<�e+B����q��O%T��䲆��[�<ҡ�$?'���G���$;j�R��~�<A�i�* bT1tǝf���j�Je�'��'�>��4kH�uHP%a���\t��`+,D�[LKe���C6�Sh�j|�Fd����z~B�xJ?牮wХ��)
%W
I�#.�%V�>���Or�>��}2�\� ��R�ܣD��{�aX�hO6��dL/�����A-I|4����6
�!�䐈nXy��V3c�����B�?����>�n
�8�F�ڥ��%i��hr�+D�H��([�Y�Jջ�`�nҠ���*�P��$pN�>�ࡘ׀��v�X%�E6�	U��ϓ7��7��X�|�3�VK�Z}��l�"��QR��H6��Q"0���'�ў��.��)�x���=_�Np��e/D�8q�,Ah�{� d�>����?D����ަE�"�Cdk(�!��!D��Zu�8im<�H�lRE��	K5!2D����`�<\&2MȒ,P�gr��b�.u����I,Hp�����31��ؒ�Q->C���M*B@�U�I��ɒ��C�I��r]�g�\��*y�Tf^�#FC�	%z;x����� � fn8~<���>�E�E4k�rQ�֎�48�@��G�
I����p6O���$�Y�Q\*����3�b�I'"O`Z�#R���+�%�8��]r"O&��4�T��P;e�\6i��0"O�L!�݋T�%
�!�"M�=�f"O�ܘc��H|:�!��	�I �"OX`��!�qMr��&� DuZaX�"O�$�����ydc^#	�qx�"OF���)[zN����#�ƠR�"O��q��H19�t�A�G�w�Vy'"Or�J��(�@���JӾx�Tв�"Ol�a㭆0n�L��d��])Hy�d"OBpx`o@��\��Ӆ�:t ZI�p"O�qeJߛ=�(�C�#B;Y��ӓ"O8�H��ԡ2N�1�-�����"O0}6%�C�lq%��	�!��"O����ᐭbW&H�k�r�乲"O,� �X�BDU3��E�ӠP��"O����75�\	�@�
�p�d"O4�Y4���+�V�B�mZnHXX��"OФ;�����88��+P+���"O��5��<�tMba,��`��"OlZR甉^Rp��*o�pAb�"O�����7ה����Y
u�2��"O�������\�~��v�?c�Z���"O� p1@��P�P�.YB�X�p!R6"O�鸡c��QTqI ���v� ,Å"O�h�ANM�(�*F�O�F�^�"O�E����h��  C��|a\!�"O0�����]����B��c��;�"O��JF�W�q����@�����	S"O\X �Hx�)�!S|m�"O�}ӷ�)'"v8��;,�AB6"O���Ӛ_�F�`�L	()��\��"O�Td\�}����� QК%%"O���-א>��r�KY�.�pa��"O�t#��;4��B�
0�N��"O�D2֣F�~��]�'(��0"OH%�u�����e�J�y�H=�6"O�:�E�6'<���,99p؋�"OحQRQ�b4�� ��-)�a0Ff�"�P�#�
/n��DԞv��)2� �|Jy	a#Ծ@n!�	(�z��4�z�Ic��Q!����0-Ќ6�ڌ���B�
M!�H _�|E�ס�AĆE��a>>5!���
�ܒ�*�P�*��fA�Q!��.�V���
��pʡ,�!��X�����C'��$��Ab�K<+3!�W!,��\��*������D6�!�� b��,bQ&�?N��h�$�2z!�@� h���8s�x<s�M�*Oh!�P�*���"��=Ǽ�r���m�!�dZ�
���K*�d�b�lV�!򄃞3���b��N�zFơ��E�8�!򤝔r� "�B�Q0�ň�C�!���O(�`'d�(R?�q�A�FZ!�dŞb�2�Z %0R;*e*��]�X!��
Ҋ��F�7.2�I%�[!�!hiBҁM,_����GR�/4!�䕤{Ur!"k��{��y�ǅ �!�D�e6�KP�8s���F�>�!�D�8-,�"�Jie����%)�!�ʿi�J`P���5ZJ�З���p�!�d�;k=���W66zL���]M�!�F!Z.U!q�O�8k��3��S�l�!���/_dMcu��(!H2��'(�6E<!���)Mi
U)W�Q0��@��B�!�Q�d�d\�g���p9x�c@܆�!�DC�3��ٓ3�3!�P�"���w�!�d@�TR�(fB��� c4�� c!��&!;�*aK�I���s��O��!��&�&q �Хv|ғ��q�!�Gv���{��_'nR���K�'�!�	u�,�e�,�X|P�i�$3!򤈟��M2�O�I�8��Ǖ�:!�Q9����e��>�ޔs�Y�!�DB$FqBQX��L)�nɘ�ʏ!{�!�DQ�xA�E�d\�K�T��U�̒:�!��:2��eqѣGQ���!B�)H�!�$�3P"F|��RC�^�����!��&MBP�����G� �3��V�!��էU������2�@H���%�!��\�ؓ�M�^@�m����S�!�$O&b���B����n!�)�^U�F��'ҠM�!�Q."i!�gL�0���2m�	ʮ+H!���0�!��쌽s�|("��Q;!����$���p%�=7��;V$�35!�Ĕ�+�.����H.�\�&�E�*!�� �<��Ń�`j��:���4/XP��"O� ��"�� �F�U&h:c"Or�Z��U�#�� ��
���@"O���g]%`�pɐ���DLS�"O�|
uIN�Kྵ��뛺(��H2�"Op���>{6����0�&��"O���0X�
����8Qr���"O��D��3f�뤁ͬ1n�yp`"O�|:l�?K̈ ���o#.-�"Ov�Ҁ�)uo�4`��I!��j�"O"�b�*'N+ ��l_�>L� !"O�бWㅧ@��`J�*K�Q�"O�h0�锵L�v�hAJXn~� �O`�^��I�d$�5� 'J�>���ӂ=�'ð}/X9�w�ƹEKJ���w��0��3`��P"�	��^)��uJ���mS�Z���Q�&E�P��bJ�*��N�W��P`�W���p��{�}�����pRE���]�؆�<���'ل���8 ��4��ܔ�Z<�&(��!�a"�)pFA�򫝵a�~�a��W��l+��Ҕ+��]���!�Aש�6=r�{MʧN�<#>�b�i�2e��ǀ�q��O������)E�� �	�0'�8��'_�<
6H�?S܀+����X��`����`M9 �����5�蟂yRƢ	�U^����	o��єA+�	n�����'��	cpkФ9���w.M4E�����X��?�kN�|��X�!������>c�4BS��7��e����D����"6����dU�Bw	yD�׹i2��[#�Ɯ]��xS�&��v��Ц��97vh���'�H���6�ȭ�3�N/ft��h#�O�xl��/_�6���M�b������5�B"=�$b�.M����uf	3R�H�eB}>���	@�7k4#�"cJ�0�E��U"
�Q�FS� �b�X �Lxu 4n0G��U6n�ѱٽ=�9BnF:,/Pac�A֚���`C�p�h���B�����G�g�,��(�~��	MҪ�r/H�"">4�ҋ[f���TM��"�DR�"+��51V,�~�7*���#�4A���l�&����:A֙�`B�4)r�ضI��*L��kd@�?�mZ�o�4 �B��@Б��"H�{x���㇂Y�l	��5D��%K�'��k0j �u`JV�'��M����8a%���ÃBC�`��J���p�䋗�95:�p��1_���A�+�dɊ6GǄ�J�B&kP< -��	׭hv`|؁J,˚�˔�Z!DO2��!lB��(O$�k֪)����t(�#AG<��Lbݩ:2GJ>M�hk�n�$̶��B�P64DիtA�6�H|Ba,�(-�y��U�O�|C���0�Vc����Th^��jBztX�	Ӻ�i0�LO�°�ߜyĴR��$�J��dު���w��8Ã�+p���%7�=����50��a�h]�\IS��2���U���'D��
Y�c�<�f�ν3��x���L��lZ�¬؉7F��)��a�0�PƅO�7��`�D�9L��T�ȗ}ը��[!J �BL���T	q�ЌX��x�d[�����Z3sj�Ye.E0@�������uղs�A�W�Tk@d[=�Pk-[0t�t���V�O6��E�v�݆h��p���jOv16�.}^�GzҊ_��]�q��7#3� ��g��<��H�k��|������!z覹�V�׵{R �G�K�}�2��n;o�tA�W�A|�����O��K�<(��Ct��QKLV���՚e闦Y��ΐ7h�ժ��ڽ^� ����E�V`Y-\!���'Y:lx7�2V�2����!t�F��b��� �1[H	\^,R+D��~��Y�A����䔼.�j��@ۑvA���Gi~�7ʞ�V�LP�I9'���B�&G�u��,^L[��x��i��R�_�xS�T����DA�
;�O�LY���/*@����3_�$YAG<4�DQ�p�V�}D)��|�s�U�U�I�4K\L�я6TS��	P\��)g���l�г��"�j#>1��?�D�3`A{T�R�������><�C��@�R�h��*_u˓�p`R�F)�x�?٦�߀f��X�A�E�|�T���g}b���s.��s�J�ΟhC���2Yp��0�R>����B0J��Y#J9�":q`e�6�'�xh��H�8N�B�B5(��Cl���'c�a�G*+@�(r��O��z��%|�d7"?��	���#��3=4~��Γ�P��&!2� ��i�X�"h�M�^��'��\s�b�CLɧ�Ԃ@Izl�'���j���3jԃ�����'� �0
A56��5�"�Z�A��Q�O>�oC��Y�Ó@�b�9����G�,��eeN�X`D}��@�f��o"J�J@*��a�0M�Ro��/�TB�I�F��Y0N�j	�`ybh� �B��vc���J�!q���8;�B�ɵe���U)S
 ���Љ�?L3DB�I�PZXX��H^+Z�@F�r�<B�)� ���G�0XT��A�8]s�up�P�<Ђj\S���ɣ������4x�(]*�nO�X������?�<t���3���(�@�0��)7gÎ0!�`��'�j�@��8��".ҩ����X�[@� �a7r"�?�z��X�g*p�j2+T�D� 4!Ũ,D�DIb�(Q�P�W��U�4EC�`ה&0p��-h<���<E��'v��t*�w(J(�GF�W���y�'2�yJ�E�<;�ja�`�\�E*j��'X���3)�z��q��'6�=�7�ˈY�҅p�b�5	�Yy�F�)�O(��/�i	do.DN��q��]�D��W�T�r1g�8)��"�,i41Gx��M'c���
%"sP>!�A�;,��P�E��[��P�"OJ�=�(H"*.�=e'ԓt�����ӂ!8`���W�"~�3t� g��5%�
���D��u��$�&U���#Q�4x��Mj���L�z%*aE��l��n�<�g��*�k���)����G&�\bf$�/�.��ʟ_w�y��R ���(Q�B�H����{��9O4x�ׄސ#wh�0�,R�c`�IJ��{b/�Q�OgQ�6�أ�,� ����J��k�)��.K�0>1�L���p �r@��BQg؞0n���T<�t�'�IY(�w�Z�ȑ�C�sjx<��'�� �S���J�>1[��ĵu�Vt �}R�ݣ��R� �q�O�4���/k�l�a l5�����'
��3E�X4�*��7+�e�����X=U؞Y[��>���>	V�B�e3��)��3V]�l8���c�<i�DŌ	��;e�E�z쾅	�,�ᦡ�A�~����v�'ۨ-ysŇ\�����y+4i��1T����Nu���@)*���Ң���ř�N�Mq!��PD�{��#���
­Y�c{�O�`[֡YRP��I.ff��m��52`lF?Cz!��T������؄w�2I�K�mz*XpU�8n.��'��"}�'��X�1��w���4̖�&�8���'r���kF�2)��l�	��	�n ا���0>1�e��L9�x�[Q M�G̋u���")�>c_���!tf�+�jH�e&�!!B��@�!�$�L�Τqv��cr*�*e�ӭ;��ɳ��s�i�����Έ�;�(�MN9C���b�.7�O���+;^%|�;���]���5.�*.y3�a?�y��Ҋ0�,m�t�V,!�5C3)�/�O$��%
Q$f�A��4�S
R���ÆN	x��ĩ�E�6m��B�	1���UG�;yq��c�.��~t�1A�_@��w�y��9O�3f��	O>�Lb��S�l�l"O��c�C�|�xH�!##Iz��w:O8�����8j
��7<O�9B
,&�L�R�aO	6N$p��'y@�!�a��Sx� ����#CȰh�GKs�2��a��%H:��2a�.�8aN�Vռ��q!T���"�!.c��m�bv�' -ړ�Z&0���c"�DE���ȓN�AI�h<)�y���_$���D�A���������s��4KE\�*\������!�t*8D�0ʣ.M�g�!8Pi@%�I�B�x� kƁ� ��`�`�Tx���� L�B���s�L��V	@���#7�OX- �F�^�z8 s��`�^@ץ��k� 8�Ї�"�yC~����=e���)���HO�'͂� �ң|ڲbO��4��۟	���r@�s�<��(В�lU�	�T�5�GT`�<	������8t0���f�\�<1��a��pɋ5N6K��T�<��nG&��Ma�3DQ�z��WS�<�t [0�� i`�ê(�|i¤��`�<��ؾQ��d�G*��!��Âa�<6dE�i~
���e�pt�(Rrf�b�<����x�^([�ǜ(~ʜQe"^�<�.X�N�9�A�� u�c��_�<��⑮Dp´�� {��ݬ�S!�� ��&#I�G�Tx0�C�`$��X�"OB�q��\���0	�H�h�(�"O�q#G%{ߨDX���%<ľl�D"O
٩�N�c��@���U��C�"O����h[�]vb���@F58��8z�"O�����NG�Ժ�hڅ@�*4�6"O����H%C\ g�G�Jqq�"O�Qr%�t{r�Vi�rV��ӄ"O�ɚ���ku@M�VH�3sE�qU"O�����.WB ��U�FUf�p�"O�Y���B�!m,�!r�W  ^zh�"O4)i�I�@�Ly�bA,5�{�"O��F�TY���+�%O���!"O ���Qax�k�KQ����"O:��1�%:�]����|��s#"Ohٺ�J�"@[�2�"O�1���ֵY.��#I��a��"O���G��w=@EH���ν�f"O�T0@��E���(3J���>I�`"O|,҂lZ�x0��AȆ)2ݔ��"O\p`(؀ %��1P%�� � "O>���iD�_`�0B���FG��"O�U�����l����j	�1���yb(�
	�H¶�P�+F�mc�-ݧ�y�W?���P.Ph$�+��y�&�V�}�d״_Z��ٲ�Մ�y���xڒe��܃S�2�a"��y�G_�7'����8\�^�����y�J	dv�a��
�z�"Ux��G�ybF(�z���U�IK2���y���(v�Pd��nѺ��^��y��DL5���e�jT��E�y2�!m��*2I�x�h��ѫկ�y� L	\`���~�N�;��@��y"$��D��ys҂K:p���I +�:�y�@4 lZ�w�Խut}��H
�y2�Qc�:a�*B�p���M�y��"\�yA	�(���A�$���y��V�!:���vHIңS�y��JO�D�;6�-V���Ĥ�yB�.7�z웳�� �`�5���y©V�W��1�NO����D N�yR+�!8�a{�'��t�Y��X��y"F6D��z���2���eAҨ�y�W�`�<0HR�^9|.���
̿�yB�7f�Td��:li%_�y�)];�4�6j���|g	� �y��As��S� �
+Mԕ�Vl1�y2j�	i�����O�$�� 	���y���9/���E�+��qx�y2��G �	`��;,�<��*�y�Eϫ�2�X���..��b`���y2��`�n�9�K�*7O��r _��y2`P�$a{$�]s_U�w�G��y���`8�x:�웳s��=sG ��y�iY�e�0]c��C�:V���aT��y�J�%�2 �a�?��1�4��y���_��d"��޸+�D�tʁ�y��ߕ�&�
T%$-�.�tŗ��yBA�J��|�á�VH� �Å��y��H�Y�z�x �T z��3��
�yR����"y�7���>EƜ(RC��y2`C�i�n�c�S6&��A	��y��� o��H.o�W(U��y
� ��Qh�4a�!	G��u� i�D"O\U���]K���C��&rf�1�"O��2��L+
L蘒�a��k��x"O�!sj2:8�	[ª+}�h�"O���֍��.w���\i�у$"ODٻ3K�>y��j�E*� |��"OXPHD/ў:��@��S��I�"O@E�G˃& �"dA �y�r��7"O���oӪ@�(4��
m���"Oδ�V!á	�`0{q��!OY�H0�"O�l�d��1�`�0aW=18���"O��iZm�Xl[�Ϟ>D�BUS�"OjX��C�7l�7D[�ṷY��4D�p�*�>S�dܛ��+����5D�89ǏJr��$O�.-��Qئ3D� KЂZ%��Z�_,Y�T��u�7D��ZF� �D���Kԥ[7�l!�0�7D�t���X l�z"�WM�>���5D�4#�N�<��-17*U�.�AKF &D����iL4p F�1D�du��&D�xy���pG���6A�l�V���#$D��[`fB9c9܁�u��:v ����&D��0�&��y�^��,���,��T'D����޳*�	�C�e��iv�8D��B��ƺ��a6cܼ!�7D�����!]f�1��)Iw����8D��z�@иzlx3�)A:_����=D�DIb��g��C���u�htP�*9D�pȵ�В~tN�#m��C����!4�ɀB�����'"Bq"-�g��6.�����bA�'�@��d$X*V�R���c�*Lp� ���T��reOF�3p�T�q�(�Xbd�	3�n�)RO$��R���'"�
�ޑ�7��"H�����y�bȼ�b�bu�B=�qHrh��Px"$^�-ǈ��gm�d�|y�[�Zz��",ة|��txƉ�EF������-Ɔ��w�)]N%2#b�Y�`�F��x'�������ڐƋ4����M��_;j� �ć$�t����\���c���Nv� bJf���]C�� 5[���&z����
�^�D�'N��y�-�h�ʁ�O��n�ҡp!'a�꼃Diͩ%26 ���-H$h����J�ƴ
�c�J��{���!��)P�dV��EO �D��O̸b�.��-T���31	���")p��Q���Tj_�{<�Ybf��
��p�O��;�Y'B
P��ubK�,�p)�G<��IRT ũ^(�,��@��t��p��GZ������):�bl�F
_9uJPI;U� e��#?�5#��Q�ҙ3"������0}�4E��K�#�X�����ڰ���R�_�4ui��).����~���+�I<RB��	�;(0RH�OܶK�B�	0Y��U��=x�MZ�	��n���Ǌ:��C�!�05�:��3'�;@��q�3�Q='&$�j����=q��M�!����Ӭ]�9�A��U~�ʓM�|���ƈ�V�I#���d�Ƽ�t+W?B�d�h ���Ll���)'X�9�J�'�:��' ��"�t���
�a]�J�:���{���r�-�A�T����j� D3�HZf���d�'� 1���O%�`k�k˵*6��P!��$��Y˖�ɐn�j]ٖ�G(�E�lk�xS�KS2nx��&��;E�����͊T�85ۆg��hr8�Ck�,�~��Y6=����$�)T��B�D]9�f�3�hv���ͯE�9�c��8��D��5�D�����'y���pE�2n�����FE�=��v��e��G�`N���� =>��'`Z8xê�'M����Q��]�2�bL���_Iy�hɉ"��4�@�Y�iH�X�G���0?�c�K@AZ4	WJ�"f�1��kA48��JEG��r� ʓ�VȨ2���rΣ?���+M4�<���G�}�@��G~�'�^HB�iƜd3���'=�a;�I�G�NUy7��zl��pweDl��)$M�U��\;�2�8�ѥJ�-\��A3Aʳ�����̯W�j��'��9S���Y��N~*���I����Ĝ/�\ Ð)�c�<��] o�2�Gɶuh���S}R�Ј?L��3�|�OK���c#�@yҭ  Ԍ�o˺nI��a�!��y�
\٦mr���[��uȲ��;��[��a��ET��0<�P�����D����e�[P<�pH�2�9�d��}�`�[5(�r�8��1�� �£��'�<xQr'��[fB��"O�)��ߥc��1�f�sn�5*e"O2̳��Z�\P6�J��:k��5��"O��Wʗ
.(H�B�7<�"a�"O�������@�k���x�H�.O���
'���d^�`�EK�D��!h*j��|�!;����WkXWbB��P;#����
�8T�ȓTX,��/�SB
�k�*�!��Fx�`]��D2�	"��N@P���(j���+q'�*1� b"O����*+�<YԧU�h�H���f� <�l���̑Fy^�S��y�M��y1�43P41�5�3���yob����蘈4���S`�	�y�_l���(3�O�<�y�I+lB����?!���b&�7�0>I7�5��]cD�6�|Q&.�9�X԰� K�v ��C	�'���R��>�16gҷ	�%c��d�?g�(%Yv%˳A�"�?�b(�]� ��u�5?�x܈�2D��$K݅>��dCWgR,$�&�N��B��u�S��4ps.͖�����i溰:w����"��G��wj!���>n�� �A�H�(�GO�nA��F�6貔�
�~�f���T���ŧ(:���*׭�:8�|��\6\��|�@`��#q���V�Y%?�����,��02gJ�ow��"~Γ̾���a�<?ϒE+���B�0Dz�!�g�FP� 哺p�p�#BƏ)H��`��S���$G >'n踢�;�OV���*�)�p�[�^x�!���'jm����;g��ɯ>�y���'r�n�0 �M*�8C�	�n(Cp��#(��p��뉒{d8c��Z��K<���ө^��,�"ܭ?\~�B&k^�C�I�	>�c@�j���� �d.��� #O;���OX0G��Oj��C��#iuE�N�2�Q�"O|L{�+�<i|��jtcS�=���)G�imvy��mν_�dd�j�x�[�#�q$<x�7 �o�J���Ć��U�(�?�QIĬ�0����VR��N�<�F��c��x��#�y����!�s�?�2DXQ��]&��}�FDOV^HȫV�Ə*��e`q�Lh�<��"�(�"����?sࠥ"$](=+|�
@����	��H��IF�w�_L<�`	��Y�EVC䉐,0=�S)$�rl�c�T�2\$�$S�:��UB�'�O ��&� r�� ;E"W/"1V���'�~���N?�A�	;R]X���/T�L�W�J�<9Pjޭ�t��'�'Y��[TUx}"���<�:��%�'"-�H ���VJJc�qR�)O�!B�靃JI�%̚y�@��։�s_PE�:D�<�0cbm)�'�4U��)#��G�����v���fr��l|�P�`�lx�;���/X�b���B�8M�@I�@��SF1�2�L�	��qQdA[9���s���򇊄P#�2�A��\hz$�?D��p㘣E�F�A5MC*������f�0r4.R�,d�"_nx�xp�k�"}ْ�B���% MέQ"�O*P�D$��e��te��b�a|���A�r�B�I;�f���˻l?h��4|��#<�֯W�z2�z�����O��p����Ey�` �pp4��'���h��[Dr�T�G��k3�Zm��r����4}��)��<y�X!K�Q��B�9ot�y"e�Z�<	�_3p9Z���Y�cl
���U�<	�Ejޞ���.��<�Ť�50^|�4j�+u�f ��l�H8���A�_2['l!yЈS0SY�Pj�(Vr�ڨK��,!��*6jdjf�|x@u�҉'
��8A��401G�4�ʶ}$D�BdL�r�qʞ��y�)i�	a��B�1��!�y�BM�`�zC����� ���yR���L��qL��U��7�O8�y�m�5z4	n�\�{�nd�lF�yB	Z�M�@�f+�3 �~H��G%�y2Ș n��5˲H�KiҤ3֭Ā�y
� v1�!%1*�>Qv���a���(1"O �! ,�6	
<�Dg�|E�-�a"O��`D��V	��b%d�,59r�+q"Ox�"Fϒ�6��VdK� Z�+&"OڵR$��y�^�q�DO/��'"O���b��j��U�b�D�H0��"O�i���ĝrBzXr�Y,��q&"O��J��M��NYH$��4��"O*D�����Q	��3�H��1"Ov�#Ì12��x�W�F����"O��Aǈ4@�Z���,�@`�"O��
H�1a�H<j#G�,
Ɋ�D"O���D� >&�hH�/9H�ͳ�"O����D�B��0K�+7�!s�"O41I@�ߙ!$�
�+ �hH��"Oz�f�O�R%�+��l���"Oz���-Ә]�&�W
5w���"O㖤׆g	n�+��T�P�=��"OC�@T�9q��TC\��"ONU�a� C��uk���=6\I�"O�@Q�S�`,:�(��68E����"O,��֯΁����`\�d;���"ON)��#��U���e��E��e�c"O2}�酜͂�z��Էx�:L���i�@�1!̉.p�V���	`�`r�H �4q��	!��m䝡`�=v�4��W�X?'!���0�� %h�M�t����ȭ,:!�$��h��ٹ��)!5ģ��\�!�d�^�����Z1jQ�b�!�D�)c7(8�u�4|Gdc��E�uW!�$��Kj��%�#M+L2F 4SS!�D��j4��`ݻFdtd�ȧ->d(��XޭK���O�l���fݹ�T�'�|,�PEt3胢E)Z�l��gⰈ�yX��`�CJ�����O�$4��BB	\���L��C?
8h��B-,4��E��š(��iIa���שG�.MT��1a��e�cʞ�j�t�Zm҅CQ"	3��];�䉋ç'�pXA�ʕ�Li ��ߚ � }[R��V�TI�� ����)���v>��WB�.lt�u�Â?��D���Y{!��nڹLtP�b��є*�X,�'�h�RI
A��9:�1�62;��f9O��s�;��p�8��퓚/�"EH,V�N�R0�Z�[���q� ١�����S�O�y��%�F�81bٛm�J$�e�'X �	��y<�-�uN_>���MUa�00�ȓ1E���Q�G�F�
lZ@�q�ɅȓsU�d�u�Ȓ,Vx|;��/�"��� �Д��
J�v#KU�.z����W  y�(�T֮9�$�x�t��0D֠8�+E5[8r�2��ɂ,#0���nV��Zw�ѓq�n��ܼal\E�ȓ=���D�>'P��%�Rh�R�ȓ��z��^�o���jCI94Hd$����H��BC�r���@ֵW&��ȓ=(�@��F=U|pr��E16��ȓ|τ��咖_�ܐ��n�y0�=�ȓ5�nJc$˸2��-�5I�12��l��x�����^<R����lֵi�(�ȓ+"X�X�.F��
4'k�}r��ȓOj���K�#F)��/��]��o���� �QY��j���DJ����m�(���%D�j�T��2� ��@�h���dO
%Fn^��XG�E�adB.|*�1�A�}BT��F74�صD�,#�hq�5�C:��,��8��fa�8��06m�=w�B䉐c�9s%$è���Y֯
.j�C�	� �� �U�>˲,�'�ȤC�)� (��b��+q�� %���S "O�x�p�d�|i#5��"2��@�"O4�)V�S(+���*�.��"Op��� ��PN²o���f"OJ�Y0��]�T(q,ñ"�$!r�"O>�` +Ř|CP;4�ƣc�T�Ȃ"On��Gh�`�諢`ȗ�H;�"O���K�*�~%�↊0�B�8`"O�|SA"'.�Ah��В�ΈP"O(�:B�^��� ���8�z��"Ot���<Y��@���*5���"O2,Y��4P�[e��B�UY�"Od�&g¬s�Vl�Q`ϒf0�]j�"O�b�F*{���zW���,�T��"O�Re��b���^�V�UC"O���A��$��,�7Z�c�ЀI�"O�����בB�t YQl��֮�W"O��@�a�s��-��J�?)��A&"O��դ�<�Ѕ���Γ �p��"O���Z�z��TY�f��O�TpH"O����\4X��8���K�x|�]�"O#��>?�� ʔUf٣�"OB��'˔�0P��/7S&,�#"O`\Yt��F$A !ĢP[���E"O����nf����1eO�і"O�Q�ѫ�n%z�!�RZ�Ժ!"O���glU�LWԁ�F ��o:��"O<����<���I��ZN �;�"O�-�2�XTf1�"	�Q@���"OB�RhÍ7Q谀3%��p�Ʃ F"Ojd��&�<Eh���`8s+��it"O���r�͝)P4� �@}�p"O�qpVǋ�Z� ��WB�>@	�M�"O&p��x�QckR�#��<�"O<-���ZA1�tZ
�;+����"Oά�A!��)��y�Ƀ>�~)�"O P��?oOv�aIC2l�J�"OrI�P�ƑYH*EHW-�T�"1"Or�P�� j�L�A�B�_��B�'[�ݠ�kո.@r$�"��N���
�'\V�X0�3�Bu�E��NT�{	�'0f��既r�~j%��w�^�z	�'eH07�K���[� 8h!�M��'yd�2)<�����=[JNU��'D01@iA7�p�7��b��8�'�ʄ3�&�����Ĝo'2��'��@[�ǛN�x�A�I�k����'�]a���N��p�Ŗg���Q�'f�(e$R1�����d��JئY
�'�reI�,��QڀY��J=E��A
�'ˬQ�sk��{�4�1W��@�'�<�%�'��@H�*NlR h��'"� b�X�Ԛ��T�2kܵ�
�'��)j#m�-84 �(N���-��'q&U�G��5>@H vk�B!rYQ�'�tU�$F�,XR�b�h�N��$:�'��m��� S����턣T��	�'߾�j A��y��SJ��s9Z��'��j󣒐4��\��!�/x�N@��'/���T$  r�ݨr��<b�	�'�2=����#��x��ϼ?z���'~Z�Z!#�4Z&��1�F9B(�"�'���֦�ˤŁ�倍]��  �'��<�`$��t���)S��H���� :��aA��k8�@5�]�>�r�C�"Ox��BL`<xtbvg�S�j@:d"Ohٱ3��yG�
cvp%"O�i�Q2|#�앇v��M��"O<���mR+i
��`ܺ3vQ�"O�Y��MQC���(JYCT<J"OV8 �h "		U�;(W�Ex"O�6�V>gJ���v�Oؑz�"O.��3m��Dؚ����$2�0e"O���F��ͤ�	��í��Qل"O��ұ"V5S�@d�gI�O�
q[w"O��C�j֓t�`e��t�P�A�"O�D�� �o#^A���N�,��!��"O:a�
5[;x�I��V�.z�w"O@��%a[aq�0أaɕBUt�Z�"OƩ�b�
4�Ru5��s> ���"Ov�A�W�"ɼ���&ԥp��ѣ"OrM��M8�p�hS̙�y��HJv"O���k�H��H�0��w"Oh�IaG�᜼"���h�U*O��S�O�2^��y&�H�c(��' ���Mr�&u��Ӷ\���'e6a���+�R���J]T�l}I�'��	�-ݨF��!�J�b�T0K�'uRXx���Z�.��,�^�TC�'giR3�#1d@y�.��!�H���'�v-��MY��D�D�Þ�jd��'$D�"���&5-��j�!$b����'�2��'�ӜTt�"��V�"@���
�'��!qr̉�5���X��9d�d��'&4�a���uOtT;C�I& �x�'�b�!�d����b�9/J���'m��h�N�/Yg���ď{J���'��(AI��m.-�,��"OΑ�bo؋$e���˘o����t"O�=q�JB!���C�/�"Y�n4�"OF!aʛ
]j���K�����"O��Bm!dD���M
�8���"Oz	�eh�t"h�p��<�6ey�"OJy��Ϙ!j�.0c ^�mr�&"Òb $Q��0�@ ���X�p"O��AЁ�w�����B"��9�"O�����8�� ��Nԯ@�\9"Ox9j7�چK���#[7�D2q"O��(�Y{b�+BG�U$a "OjQ�Bd�"�(Yw ��3���T"O�4�`�,xs� "���
)�H��"OX-s��)9�p��τ?��-�'"O�Ԓ&LWPfN� ?�"O�Q���(r�x+�,U�K+�Z"O��I��J3u*nI��ׯiT9��"O����H�e
�IA��Z#���"Ozi� Du�ܢ�闱?�T�`"Of�@ ��"�n�Cq�<o�q;�"O�j���P��!8���=V�%�u"O,b�O|/������H�q#c"O����	���KvL�%^J�Q�e"Oi�gC�#R�#���7-�C�"O��Q&E]9lU� 1cȶ�Z5"O��0��-(�b��&�ۊ�1�"O*�	0�(C��M[V�X�{���W"Ol�"&$NW:���F�/vs|̓�"OL	c�]���`�>m,au"O��j�M�%q�J�s��:S��j "O� \l(��=���׋/H��cg"O��R�"���IF�C�0��Q�q"O.(���G*.9��@��Y�n�S�"O�|P��I�a䪑{T	 w���PG"O������(E�ڬ.B�c$"OJ� �o�t�a�lQ8 9��"O���CĀb�VY@��N����"Ov���[Dg ��&	%D�f���"O8-R�B٨hI��0��9�`1!"O0Y!"���v��b6�R'n�R��"O�-[vC�4#�Є��%	{��"�"O��#Κ]%&\�3�ƀ���k"O���a�q����J� .�����"O*l@�ą��Aϒi���1#"O�,��'F�-<hm��#׫9�켲�"O~A(�ҝ$c�{1X�p����"Ov��� J7����=-�P��d"O�(9UG^�DR��#��M
���"O��f �11�����6M��,�yR���ߊ����xH���J�1�y�%��;�Qۂ*�[zm��T>�yR�FU3�ڱ�˕x��2W�΋�y���BkD�(^���V�۶B�p8��rKx�.%��y#v3��a�<�$d�����g�O|ABqk�\�<���>0��Ҁ�2Y�P�d�m�<yp"ą'P����T1`�N$��#@g�<Q䎊�2	J��f(0y<�Q
�c�<	���de�hӵ�V-{�ƍ!��ZI�<1��@�Z�����,N���n�H�<�3�7�d� �_̼`!�D�D�<	��mxU���,#6D���K�<����cB"���ӳ�ҵ���^r�<I�ᐴB��e����+_b�5�j�m�<�T�L�%V�ȣ���l����l�<Q��A2_htq� E�D�X�����h�<y5&N�������].Z�����LI�<��f�B�:��[�9S�9��`@�<Q�f��.%��C$����r��}�<YQN��'��DC���q��x���D�<A��"�f�� �?A��꒩C�<If��s��9{v�Y0��H{�<)��]�/���$HǗ
fq�mEv�<)I��_>Yp�`P�/
���h�o�<a" ]:��|�2�F/>}1��[i�<)�ˇ {���k ��	dpa$��d�<����_X웱'�o�<�h��^�<y���a��H L@t���Z�<٠)Cr����!�ds���U�<)F�8P�����?�Ev �P�<��.�M�0h%%��T}Px�v��F�<	$C�8�\�y�+N<*�&���E�k�<��2N<�`N�L�c��S�P�tyw�r����?�}j��?y�46�2a ���搉t��+;�4Z�_M���O
y3��L>)�f�3 xE����O��V��!u��#��=}Z�l���U�U��Ybw�;�ө�y�/�"�lTP�� Ѥ�bd`�=�d�D�O�|m���\��>���cj^����������+ׂ!��W�����1.i�!'e�!T��e[�θmq*�'���^�m�ן0�ڴ��I��|6�ؾ����Ê�Zt� �+){����0)t�<l�Ο����%������C�P:1����!ݦa/d��֮�
?W�e:��<Xj�@Ō��z����$�Z�nڼ&�h)!�v8�\�l	�����Œ ��B��^rb����d'�����T'��P�Q�h��Pb�#8<�"ƌ�
ېx"FעY��5b����#��b��$=�DS����Iwy��) ���)� p��Oφ�j�j��bf�j�������o�i>i���da�՗��2�� �L���(v�v��Z�G4lO����A@�<�6��	ĶL
T%j7��J�N�T2tj"j�8t0�p��e6�Y�ҥ�	ڟ��3��f��`�"|����2�*faJ�	wyB�'��w�O&�
ҏK�̉se�D�v�%�
�'�FlR�Re�c�S�O�bmR� ږ�M�۴�?���,��&&?U��6��O:˓���Td|��4�[�w 4i�lݹ��O`����W��Ob��+�	_I�P����)���[ܱO������,O5���'3�'�+�,Ob�y�b�%���)&��.{�2�'��O|��LZ�h;�&�+B�$���i�1ڼ����'�ў�NR�M��<��ɰK��
��؟`N�z�Cp�����>���/P��0���(m����I��@��2�MaӜ��<�O�b�'���i�<�A�BI�8� ��}�kbj/��O�b��L>i�nR`v��
��W t���Rɂ�n�fy0e�ĴV���i�'U#}�'U��
��[5*�r�L��1�,-�S��O���W`y�����R�r�3掀�U~q�� 0N��`��c�"�'����"`��ICx�9$��6WH���{|�8�oZU���
�4�J�``�1C�����;v�<��0�X��i���'��|�O��vgG"(�������u$�mq��Rwwt(��J2�O�1J!+H	U�"Vˈ �pH�`�ij�� "CǌP���X��'X�80a��/Q�́�@:&"(��4&X��ٟ8�J<���?H<9��@�n.� �f�XF���B�X��-�O杓p<dqC�G�EQN���dޱ�M�O>��i��d�|��c�6 :  �   y  /  D  U  '   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=��J�E�TM�P������PŌP_`��7ju�r�d�O���<�'�?!�Ov�%ʢ���)�-#�E��-�����L9B8��	�}xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�z (PЩH��ɢ(�Zc���a&,O�$
�-ڼ1V�pU猤IV�u����B�ayR�BNj$����n ����ϻ%���OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O�����KO���O�<Fz�O�r]�pc�A�,�̨B��;W��)�1��jm4���?y���?)N>��T���GN��fg�h]$S�E�'*!���><`D��E|B|�f]�p�&��OnTh@�Ƀ ���S��;��L�Q����bi,�Oڤ��E?:���Aץ>k\�s�"O�����E�"��ƀ5h��×����'���e���M����M�@$S���ī�턙ZPyç	hBY�|�Iܟ �'����bĜ�$!DѦ@{u�@��G�Z��1DG�=�2��,�=��E|ҍ��NƤI��ןa�N��A��>(Ҹ���1(n�Q'�X� �	�i2��O�����'�@7�O�6��<��3�! �kUPub$�R�?k  ���,��䟨��\�b��&Z���T+h#�8���;n��B��@���P�h\�>ϐ	��$��>�RE�OD�G=���i'>��'Q��C�I�*�P��N�9��te�'����}����;��)��G#�e�R��-��`�)���HOJ��3g]�DF�YS��)
xѮ�3�ޏ;M�Y�'O^��'v�P����?����?ɉ��DT�p>�M��m���4	߂��'A��'�������(fZ�`�ʊ�u����ǓY\Q��rQ�:������/:j4�����	˟(�ɶW�t��ޟh��ϟ,ק� X����z5�|� , E(5۱矖n"��XSZ���d���g� ��)bH�/MªL��ЫFⴳO��2�X|R�
F�,��*##*�S�v��	$D�Bm���(w����t�@����&�'� Y[������dp�Ȕ��X�������aQ�LH<I�+�E��,����O�p����K?	�K웖fg���|��'�B�O��A�)��mIR��1�T��Ek�0�&p�ڴ�?!��?A*O�)�O��$�U\��
�F�t�q�1�W�Q\��5#װPm����'��Q�p�L�N�<M�&�J0��uv��'	��(Q׍�-~b����ҫR�4�3퉼"��h��X���Gwȕ��H�O����ɦ���xy��'�O�1`�5xq��h��Ձ����"OB��1�P�	cl����M ^V�<B+TI�	��MS����?�p������TG%R���
4.��B�$��?�M>I�S��򤙻G�4Z�'�� �ؔD�8!��ik�=�P��R�qЉ'e�!�d��U$pS'b۱'�If�w�!�X�x�-˗�V�_V$S�GE�Rѡ�D9<	ra��8=��,*�g� 5�H}`���Ȯi��>m���H� ^�4��c�0#6�d	���6�?	�°>����Z?VУ�MrcM���y"N��@5%�! �8�<��IR�yr$�@匰hGN2�~X���Q��yr� }_0:P�H�.�.0X��p<�7�	��R���q1� �F�*pd6�IK��#<ͧ�?�����kP���!�4Ӳ%s$��15!�d� ��أ9�:���`A!�D]�A��e"�-�+���C��G5d`!�	-q]��G�(�#� ��l)!��N�k�^IK#���$Y�f��(�����?U2�	�2�Н�3`e!���$}b��]�B�'Rɧ�'U�0a���@�r�I %c�Qv����d�E`Y���@��$�@L���.���H�*v�=�B�O1���M2V]�2�Uej�a�fIX��5��s���u��bt���1�]�i�=��ɽ%2���'W��eP��W�a�Z�pI�f6���IB��"|�'C�\t씙�eٖH���'�����ٚ���.�?�
�'.�TK���9���J�(L/��LY	�'p���̩A��nB�<��z�'G*�b��)��e���D�	B���q�~�'��Tc��i�#@�H��$�#��5Sd��9D�<���x��I-� s0�Ǘ(xX�2c�#�C䉗'�Nu�1��>�(����I#i�C�	���a�s@`�@�	�y�2B䉏=l��S�H,M�X5��� Q����ĐB�'J&qHt�X���b
*�ƨ��'O^9���4��d�O���h�[�D?PL$Xz2.¸2��Bڀň��K��幒�����ȓA�XSX7`d�1&�Q9p�@цȓ�8��g��*�� �Ƽ	A��ȓ,:TE�����ּ��LBR��p�OXPFz��D��$�Dq�E�A')1�@�È��	<1����ɟ�&���Z(qCD�gg͹ F0+�"Ox�[�&��Xb�uc��'5��0"O��Ѯ�4�t�hO�Np�0"O����G�N&��&*@!Y�T�"O�l!�OTe���N�i�d)w�DK�'�4���o#���v�D#)�D�86�� m��6�'�'l��Y��Ɂ�U8v� ���pf���Ш:D�p@'��(,S��s�#�z����4D�x�B�ң9M�mI'��=w_l� �1D�(xrN�T򔄁1`�*g����a1�� F�/�F�����k\r$�M4=�Q��F�;ڧ�(��"!�
m�z}������)��'r�֧� ���D�һ`JN8a'BA@"z�h0"O1
b���.3��K7@2C0|��"Ob}S���#V;�xQuOþz(�ŉ�"O84�M�!�Ti�##
V�1��'x�<�d��r\2e�1���n�Cw�O|?e�Tp���$�'�rX��:��*��˟,7��Z'�;D�di�lN�9���݉|�T!�
<D����
�Bgn.�Nb4D'D�h�ю�q9�܀0�x���g&D�,����W2�<�" Z��`"�*7}"�?�S��-$�H�Q�ݟ@��x�� �13����O*$
���OL��&�����H�F��'A�R0Y����y���1a�8���O�ay@�yReS�6��1�D.�E� �胅ܽ�y�J�%��pv��=>�R���@W:�y�^�Rĩ�b��/�r|s4�W���'�@"?"@�ß�1�)o>D�`FgK\��4�W�?qN>��S����U�3(H�ID��-p��eƚ7�!�_�yfh���6t'���d�k�!��^�2�� bSd@�x����i��	�!�ЀIЀ��!"�����$�!����h��`h�`�# $:�`TnH �d����9y��>a��㇧Y���BK#
6��u���?�����>�!��E��ى�V�2��� K�<����J�`�b�� �_�<���Ɔ!U}�X�$X&.�MG��r���YB<m��S�u:�p�㉧�(O�h�w��/�<��T�=k@-�"�O���Q�i>9�Il�'Gx���SU���#a�4R��j�'+lx��MA4.�RԐ�@H����'x.ЊvΈ��t��G�K8���'�R��I�
E�H`��Õ?C%��
�'����#�� -M8|�3�!SU�5�N�������3��� ���v�����( )���X���?aN>%?�!�C�}�� �h�3}�*��c�,D�aP��+r ���LǪh$�@�I,D��І�]�_4� B�)�v��|F�)D��0�B�z��/�aX�A�-*D�p��۴�<�Ui\�O`H���'�<��OV\6�' Ƚ��`����4#�)��a��O��O���<�`ac`Tyag��P������h�<��+�B9� �:@ht(�d�<Aң��� 〮L�v�֫D_�<1��H�t�Ќ���ސ:�<����Z(<���߂IA�|z���,u�*��K�'{��>a�X�O�I���a��a��� ~�L��@�O(��?�OH)4H�31�E
ìL�Y�m2"Or`����0^O�Q��Z�G����"O�]tcA	+ :=q�B�z4aG"O���,�h��E����.�>X�`�'�\�<��H�pO �hD�%?��Չ�A?��G�\���T�'_�X��0�׽p���j�DD9TZ92�+D�8�1�� ��A d��1�N��0G/D�@a׬A�@�eQ@|��Dg8D�lp��^_��`�u_�sT�H�k6D����٧s:(�%�O�ya���d�4}��-�S�'dX��h�^vRT" ӑD���OYS��O ��"�����1[�B����z�jL�1N��y�*PW�ƁV�"x�l��j� �y����#��q6k>:j��ֳ�y��;xI��`�#A��&�Z���'�y�+H"	�-p4�˳s�8�����'��"?���П p��^e��P��'//D)ȑ��?iM>��S���D�8�ƙ�1�!����W!�� ��)�Da㨼i�)�:���%"O�@��M&\��a�H,c�Bm;"OR�P	�<!Ш-��F�
!�p
O:�4	Q˞L��� H��mL���O�+G�Ӄ$YH��F��I���t|�=@���?��xt�	��'r <
����Q�������U9�n�qTeF�BXm�ȓ�Ρ	H�~;� ��[�PtdE�ȓu��E�F�	8 q$��s4z���	��(O��8�+�/.rP��E��y�h(�O��jt�i>��	ߟ(�'�ݰ��Z����Sc��'|\xpQ�'����׏�?.���U��3lk�i�
�'��=��O�/2&iCa�+jRT��'v�d�Iڸ
���6��f�" 	�'��а2*�T@.��L�32��PHH�����	H<��X[.ƣI* R��v��8l��K��?IK>%?��2���b�@"�Zq�����!�Q?V�*��Di5�=���5<R!���8�q���Al!�h�+�
.8!���G�@�SÐ�#X4�7�!�Dݐ9=�Yw
ܡCZl�ْZ��qO<�F~b�Y��?I��ς`�#�
��b]5�_�d��|"����	�7jެ�1*��`����m� e��C�W8��䅞3���؃+[/��C�I0����č�'`���G�;m�bC�I9���S�U"hohY�Ձ�W�B�I�5q
�����f�\R��(T6a@����a�@�}��[�c�"��D;4��B�i�~�2�'a}�AR�*_�D�R��D���B4���y�G���)�O}��w�O��yB)�97%L�2
��E�%r����yr�N�>�t�s�F7;x��Uϒ�p<)��	=܌�A��M�F�z8�s %@2��Z��#<�'�?����$^4V	�eJ��DU#�H����F�!�dȻd�TM0���8V�:�0T!�D�G2l�`#��'F��1G�iO!��.P�0(��0@����s@!�	����	Nx�Ɛ���R*�E���?���$¶"�& Xׂ��6d�`*"}BA�L'r�'$ɧ�'^-��j&*
�|�h� LWEy��ȓODP(��ݢ%���l�,���7��yIg�H�"��S ��4Wu,�ȓC���8��[�(�# .\�ȓ<*��%���;T ��r�֓.:���=A��I1W��DK$S�hq����7Fx�{��0ZӴ��	S���"|�'ɸ�`��:a4�X���C
�A��'0dl �!ZB;>���*�`y�
�'� PåG����
oE<�	�'6�5{Qo�!#T%	�L�/1�,��'d���"�`��5�Ć䳢�~�'�����i��y^$������K�P�GA[E�L�	៸��I�\�2���I�$�u�%�T�#*VC�;?*��{C�[u��cj�L�C�	�o7�=af׾c�H��b �/ �C�I"�r$d�#^� � ��ś<����$No�'t&L����O� А�`Ќ{���+�'{B�ي�4�"�d�O��#�����5!e�|$)��bЂ9��Gd�����El�� F'�)^	�@��-l�e�1�8ErL�e�-����
�� ģ͔a�(�=_��ȓe"%(À��uI���A�&Ѐ̤Ol�Dz�����9����1��~�D�v����R����şp'���
HR���l�tl����r4�tB�"O���%�V<"\Y� ��B����"O� 0��&F����a/�5|$t�"O�Uqcg	/S��qU�[�hnD��"O\0+S/�&(�q�o�M^H����PY�'��ɋ�7m.ly�l��j��]��$Qc�ds��'��'��Y�t�W���q����!�zԩWb<D�Ԙ�mB�nҔ�.�EnJ��7%:D��� 
��C&��S�U�F�R�3D����Ҿeꄡ����2�4�iS� 7����<WԨe�?X�Q����'�'G�Rٶ��3�������yub�qT�'�"�'oƔ��ط/ �0�s��*� ��'�n��pG�4�"���0u�(���'B�,ȵO�sG���$C��s�<E��'�αK"�JY�Ҩ��K)r���(ǓT�Q�,�ӬW;M\k� ӯi��f��@�'gE���d�O��2�2W�@��� LN�g h �O&W�Ȥ���OD����Z�g≥U�N�)���72z5e�N�yGF�"��P
P���	P�'4�ф�)�3��^��+E擹f�n,["5*�p��I|~�$(�?�'�HO �� ٨V.H�7DE=\�h�U"Oޱ�C�G�ZU£��f�� ���>Qs�i>U�	d}���2n��+�k���K7	^4j��ᢟ�8�	�P&��O%f�!v�6��Ҏ��l���+��V� �rk
�p���'��T{�
��?f�%R��[1A}��y�
[(c���  Y�G{f�b��'����D�l*�	Jce�#�b��aD��?Q��hO�b�x�C��Z����G�)��c�"D��Цo�$# �ɗ$B�e��!`�"�	��M+���d16�lx�O웦��h�����_
	�H�C�铧 �����<����?1�O�~��d�ϣm��US��� 4x4Q��O
v�ؤ���jW̉c�=,O�� C<�b��A� ���9���4��r&�hWo蒥a),O��� �'��\�(�e�X��Yh��H�R�%��H؞��-]���)sCG^t��� $��;���A�����������䌛nnu��Xy�T�X��i�'�?�J~b�4S��<�5͐6
��aJ�X.�0�'���+ �J���w�p���-�O��K�Te�[�Q�d�ѷX�B��U�3�ēGނ!`�Tt:X�!Dƨ�(�:�(�R!7O�8�TꐺD|l�;$�xB��!�?)���h�X6m�-G$��.�g��8���QC!�d�vNr�� �ʏF"Ĺ�7Ŗ'�xR�<ʓSi^��R��5|���QV�R.!��}���u����Ob��S���D�'�R�'��I���%Q�L�Ę������B(��&�H�!��L�g�I�O�R1ۄc�W��X�v㖲y��$��.Q }Vt�3�|i���xr��o�t��O�#.�(hEn��N�\�$/?i����SS�'y\m� `:}���dށU�ؤ��'v��R��/KP�T���;a��XQM�,R��4�L��>��%S ~��:��Պ&S���gh
'{� ��n�:���Od�ĵ<a��?��OP�x�Gl
Wv"�S�lM�!(Ta҂뛚M�
 !�w�`k��'�԰q!�
?7���5CӊoJQId��#�vp��mR�	���'�pؘ�A�f�� V��<r�2
���?����hO�c�8"L�W�đ���[�>�*�p�?D�XY`��&��X��{�V��qO
@nşL�'�l�C �~��4-Xᑀ��=�z��N�/)V@�"�'��	��(���|rq�A0)� Ib��Ú"��$��B�ʃ�T4�^�q@���way��4\[�=Ѐ�V�GE,��3c}Q����+�,���ܑ	���$]�5q��'!�	�m@�d��l�*e� ��¤Zs�t�p��I�]���#h�3V2ൂF3�HC�	��Zܺ�I<G�ԅ���3���V���ܖ'����[ir�����M��@-.�舘�D���)@G\�z�b�'���)�j�/u}*���4�r�-�@����C_�Z�$����˥O�r�!��
戟��z�k޷i��ӱ����TŞx����?9��h�x7-Qd����Ÿ]��%�1�с3G!�dC(��XC��
1�b8	Ta�+D�x��6ʓp�Nl�_*bn�C	I6:�!��?A	�&�$�  @�?�   �	  �  �     �(  ?2  =  %H  :S  _^  ti  �t  �  ˊ  ��   �  s�  ˰  ��  ݾ  ��  m�  ��  ��  8�  ~�  ��  �  O�  �  ' � � V �  '' �- 24 u: �@ �F SM �S �Y �` ,g m �w � �  ֖ ڝ � _� _� �  x�y�C˸��%�RhO5d��p��'l��ɶBy��@0�'�F��L��|�t���pd��46b�Z�4?NNqhs��|`I4jE�M�6��"-_�7RN�wk��uGjY�7���
/Y���F�6=b�l��wm�u5�@%=,ĥ�t�X*v�"@�#�0 ��'��O���]37�,����M3����U�̳��A#['�QrDM[Q��=�2�I5'�lÚ8+J��E�Ql�6�\<9I��d�O����O����.~� "G�zʤU ug�%w�����O�RP޺/�pʓ�y������?1e��RfL��篅�t@���ɮ�?������?)����'��$��fe��"�[�AߜXJ��[ !򄟤Y?P�����{ʠ�z��+K�J�"~d�CP��(e2LIcP?���=O9�)�7(X��yr�Є:���1h��(w�HBĭC��?���?���?����?y��?i̟����Q�T����H6&c�hz�'w87����M�ڴQe�I��M�i�6�|���WW&`�sK-n�h��AfىzN��Ї��j�4�rt&��,`�O��f���d-�.���Q0ϕv�Dʃ*��p���I\����҈iB�R�x�4uqNN�I�1�aD�<��2��h{�_�b�u9�1l>$F�\�L�|��� 10C`x���Ȋ�9�"�G{��	����D�ǢյO�t�t!ʌ��=	������oX!VW�=������<��)�?�M>�������`������j0����*U�<B䉵1x@YA���X#N(a��ԃ{/�C䉉"p�]6�ψ���e���0��C�I�_[.}"���̲̲�-�3t��ğ�B$�#����V��Ir��#;��N�F���^	�^T��↸6D�z�@�5���'>a~¥ܯp�xd�5k��9l	 `#3�y"����a咻�xc�&0N�C�I�C�L)�a�Q�Fr��2��FtTB�ɫ�E�P�	�$���J�?����x�����n�˳H�	���d�4���S蟈��d~��K�}�ɋ�l�H=T�0�y�藻g4^x���P�Lɰܪ���,�yRM�P��*�ꉅtİe3�b�*�yrF۲���(bJ�q�4��y$C�c��A".
�jdԂ������VG��(���:D퉲? |��ń�72f�1WV�|��֟H�I]�)�S� �Q�	Z����җグ �B�?e�P#яG�-��)�`��M�B䉬D3ĥp6��30*��9&葭��B��-P���KG��"ОѺ�+N�32�B䉆a~�AX4�T�H
s%�E���OV��>�� ^�Tl��'fR���[�~��S�C��l�8�ʹ]%[�����ͧ<C$����Ie�LK�Y���HH�[��¢;xH��I4=\X��0�	�Q���P Թt
�qq���!U����Dֆ��'���'\F��Ua��^LAPT'g:� �\���I|�S�O�p⢚�/5`�I��B��x��.�"�]�r�6�x&CK22F�q����3�?	,O.T����O�?�����˧l]
�$�d��P���lVޟ��I� =���3I+�)�'<�0�A.ǌ7|�|���Z�p����'-ܠ1��i�S�Oņ�u��
�.�q2��!.Py�OTU���'pr����� ��ݐ�%+Ntt����.[��'D"�'ݾX�AnŔe̐hq�(�m��$�F�O�8C��M��xQ,0}��Ի�{���ʌ��O���'���/
n��6��?!�>�Ӓ�ѻϸC�I�s�4�c"S-LzE�47��C�	�@�0��hS"�ᯚ�K3PB�I�7�
�� �&o�D҂ϓ�l�B�ɲ3Ӏl�P×	!Q�D���R���˓ ّ�"|�s�l�Ԅ��&T:a�#b��l���?y���?H>��Vi�����<������b��z�	�f�!�ݔ&��!���A+^���k��\�,���9�O�%��H�,N�`C�g�iK�U��mz��'l��'��)�<�,�<[,����`�"I����yb���+Q�	�a%��tV*5�6�X ����&�'m�	�1��	v���A
�Y��EL�ߎ-��$��?�L>����Ԥ���O� ~�{"Y�@o�IB��'$\)���'�4�[����O(�,8C#�<er�ѣ%F
2ax���?)��|�"��X��X����y�$�&��;�y�J�s�^���L�r���g�4��?���'����a!%0T���6��O��L>qAN���'���'<� �lQ�r9RU��K�7�xE�5�'��B_*̜a���o�8��\N	�鹢�O��S�M�䈙�	�<i��[�]�B�;n�s5H*&��pЯ���Π3���z�'�}J��Ѝbrp�(Â˧<�&�'�����~{�V�'�2��4�'�\��bH�}���Kr!�S��L��'���'��'���bF���g!�%7��Ę��d�g�O�TaBD�	A>�z�E�70w�(xf�iMP��b2!d����<�	k~�"I&H �� �ƅ+� ���XCvD�O���b��	:�1�1O���/�_�V1y�mO?=�f�z����	�J0a�)�3�e�` ��
-(�H%(�H��{,�D�O��Db�d��4�<���p��ױ����E�
?�ܐ��'#ҩ+���k�Z���a��-��`�,OP�EzR�O^�U�pI1O�/:�Ęi��`��}�t���\���4�?���?Y+O���O��Dϛz��U34 �*z+0�����38�x�	ċ@(SP˅��p>���;{�<��$��ޠ;�N�d:���Y�y�Ђ��	&g� E�&�A��uHu��EeRP���PG�)��������	��M�����O�㟜�)�e���j�^s,ѣ�Wx�<�6L�'����M �ޕ"�oJsyr�'�r6������'��)��>��D x�卢m�Ҵ[ei+� ��������Ov���O88P.շ$��勅��<PǕ�4`%h�"�N���i�z�`��mO:��{�뜼~�2y"�͖;�ԕ�k.u��HVZ}��,�e�'�&���?�Եi��i�OR�q���WT��$�7bn�	ٟ��?E�l̘<�z�H��H"9'�� ��M����?x��$���>z�Ƒ�q��N��|R�'�x����U�� M�hX�4
��lN���b�O��'�O$�p��o�0�F�L&~��Q�"O�1FA������d-;�|"O�0@��/Mx���,W�6>̼"O�љ��3p8��b��4�e*�����h�U��#1(<��ƭȺYY��'/���4�R�d�O��8�e��D�:hD�z���t@����<p�&��c��jѫ%]D���z!�a��+����}���!y$��ȓS�RI˲oD
%����C�!G��ȓ7�I��� �'�bt���U*+�≖'�`#=E��B��*^��8wF����Q3�+���g~,�D�O�Oq�<�B���.��Ze��2ffԅ@�"OH9�W�;�h�����*T�Mj"O���tnX��ҍ'=FVܻ�"O�=�wC��M�Y�D܌}&��k�"Otx ��MT��&�՟uxh� �|�K*�E�J���=��`#yZEs����0fj,��W��֟���O�����>Jh�Z$Ky�uc"O�]T�_�T�b8�Ã�{��!Zr"O�h*�e�!"F�T�Q�dw�4�u"O�LgIB�wa�Q���-][�L��'� �$��+Q�%�2(K~M@!�=Uuў(rP5�'(P�\ۧd�:[#�c��Z�S���A���?1�pj �ST�m�fp��h�!K$樄ȓ"k4ɐ���&6rx�@��H!���ȓA�vݪ��Y�4�H`�S�Vf�m�ȓ/֬�텶,�.xР(*�PD�/4�'q�J�k2�e��B��r%�O��+B�i>%�Iޟ0�'Y��{��w�B�PCh� BhD(0�'��ase�&H�>)᢯GK28S�'�~x�3�
C<d�7�T-� �p
�'����nȁ^t��F���J��	�'��s�43'
IR���iV�*O2aGz��	�{��d�ͺ|u���M
z;�I�I��Iԟ�$��>5D��S�^��D� 7�8,�T�$D�� $��l�8�0���^�ur�"Oxh �
fڅ�.O dct�i�"O$�@Ch�%\�H���MD,jP���t"O��`�/D��u8veX"/dd��|��'�h�L���g^��s'�*,HNZR��^����~�Iğ���O�PyfCKB�h@�3l�%����"O��Z���HR��,|g���"O��	w�N�I� A���įwg�0 �"Ot,�
-s����Շ�jTHH"��'���Dφt�������uTX�J��L�A�ўD)D�"�'r��RJV���ɀ̓3�@DR��?��C؂P!e�B�xl������.׈8�ȓ2"����͐"?�R�x�����ȓ�T� B� �x���e�#b|�Q�ȓ|�i0t��__�����ʥ{���ER./ڧ`/nM@ ��9�9(@
�Jo�8�	�{=�"<�'�?q���Y)i��r�V�0��2צ͏y.!�{�>��(�!�80!6&O85-!���h4����[�]�\<��.�)'!�L�C�H�B�K
,�t�b�O��n!�d�8�@y1�Z�<�6�`��Xs.�	�HOQ>�j���Q��`s�(^	Kԭ���<�t"�?Q���S�'"��Պ��H85�@����`ppC�)��	��b��>��`[�*[:��B�I�F+^Q�5b�n^��z�����
C䉒4�k����jf�,h�ņ�C� ?�5�p�4�dE���7�1O��F~"ĵ�~�D��D�(M�e�ý$�sc%�?�L>y�����IJ���B��5l1�G/K�B)�B�Ɉq��g酌U�}!��^G�B�IV�����-�����	�A�~B�	�<�Z�#��͟LF
��t��o� ����ş�Iu!ȃ#ü��D� *V�2V�1ړ9���G�$ڥ2{&)����k���b� �6k���'Na~r.ȧIc Y���A5�a��&���yr*Z�����:Ѱ�X$*�yR�S�hi#��o)`�k "e�ڼ�ȓ*��`
2���[��`��Z !OJ�Fr�7ڧw6\z�n_���0�Ȁ 5�r��	("<�'�?1�����$K�h�T�ʒ:��&iM'7!�ġq��!��?���mՌ:!�$G�p�f `� �� �+v0e�!���U�P�ր� Z��A���4nN!�Dˁo�p]�c���nt�(�W	ύP�I��HOQ>�i��<b�e+ro�k?��b�<a`B�?�����Sܧ\�e�F�J�\��E 2'�����ȓu�Z���M�Q,����!��J2V����<���B�>ĸi{� �U��m�ȓq�j�`��?)������*G�Ԇ�7/R�1���-<E�D
SzA%�����Z?VB��݋wߢ�������iu��~��|b�'���O.8 ��Ä<���+ba=zN�@�ȓ��Z%��$=���-������m>��y�"
�+�.�괢�5h/�ȓ`�j�i��� ��阮@��]��	*�?����1m�}ؗ$ ��T�0��J�'Վ[��ɘeۺl�c�̃0��(y�f\�@N$���O�����'����H7[��#�mER!�S݆x��܅Sy�m+�I�j�!�3���26OS(��H�!/�!�D��Jm�a�U�D�c+�4
�џ$Њ�I�[���iD�P,4�Z-��J�_�"�&�O��O��d7?q��Wq���&dM(O�m�F�Cl�<�.
5]^�	cѪݬq6���a�<� D�r �M �)H�i'Rv6��S"OT-I����y���ϢM[P�P�"OJ0q��	&n֥k䍁�5KH��Z�������G�$s!�Q(@k��W�K=:˓9^�P
��?iL>�}C�N9Q� �,�ڜ2CkP ~�j=���� �oª��H�F�l:�t��\Ҝm�"[�"�|�pWL=+�Y�ȓ=��XJ_�P�BE	�7bzpPQ� =D��Mc)�p� �dd��荹G��'�#?�)\?�ņ�3vuBo��B�t���x'����w�g���/���&!�ҀTb0C/�!���_�p�x5$�DD\���%3�!��=�đTg�h��D��+|�!�M�K���0U+��#�����`�8\����OZ�7C������W�M�A�8��v�	iz"~�Q��V(�4C��g�FH�+��?i��0?�e`��- �����E�L\jؑҢWc�<��B�2Uۥ��0SF X���]�<�T,ۻ~�.�R�Q1h2���\�<�`dA$g^�R���*.��("�X�'nb�}�D&^t��ץ�RZfx�Țٟ�7��|��?��O:M�����NQ����"\�4"O�0Z*�Wc�8xsK"O���#�"O��R�V-D~�tf昰p��R�"O�uJg�^�qo��٥nQ�X���"O���O?1����F��\x�R��+����/a>���c�CN�֨(5��4@�p��4Q���?�I>�}��`Vd1�@�6���'�x�<)b�
 8�x�r��v,R#LN�<��%A-.�l!�ܰo1h9	��_�<YfԢ`�lE��n�#x@�X�k�S�<�0��j]�d� G���4��1C�M�I��Oc��O��	�	�^ʈ�F$�j}�{$�'��'|"��>I�`^1<R>����P$�l�"�K�<�-<y�����BI�l���C�<yE�D��]
�E�$-e���U�<1�׮VM���h� ,�05qգM��,��<��DPdiʐc�p8��@2r@�E{b�� ƈ� ���C˼KKP�!(��W�N �r��Ot�'�OL�H7��I��	!j"��"O�m��Gt�`H��FN�k;��*�"OJ���6
U��dR�O�N�W"OD`ڢ��Ʈ�!$$S+g�[�I��h�<ԀeL�j0X���Bړ(^ْ�'�8�S��4�b�$�O��7hdAL�6A�����:�b���)6�Ke��Z�� 
�"SZ�ȓ��%��o,�V<Z�F2)�j��R��U�3�ʁg��ةL�Z�6a��Yʺ��p�Y��ԙ%ǄJ����'��#=E�D�!R�i"0�ޯ]�����T���d�@t���OƓOq�6X��"��AifHN%Ѧ!��"O��7l��p&��[`�AS�"O:�s�'�ly�@�����*C�sP"O*x3�˴'3n�R�j�w�f\ d"O�öd�xs��q$H%O(q�|��7�k��0�-�ĩC� �U�h�Y���=8�h��~������O�X�a��|>�Bf�)qX�S�"O� 0vP>Px��C��:M�$,�P"O>�##L�!�����Q�_���"O�����\�HcL|D�	1&��r��'�n�$��:h�5�7#��3d�Awo�3�ўh�TD1�4&�!�)K�9D�q�R<������?�i�&�0�@@�6z~�8E&�
���-���O~ ��@� TG�Ti��S�? "�٤,V{ �)vG$����"O~�{2i�-!�
�ħH��ta���	�h�̸
�e
R�B�1Х�0Ē���'�x\ۊ�4�����O��G���yg�L�Y��ʒ�)j7f-�ȓ_w}���'�I"�$��8�H��bO08�p�\�q_4�6+Bs�^�ȓa� �r�k�nl��I�mw~���E�y0�m�.WY�]zs��?����'D�"=E��-�':���1D�?I'���RK]�����v&�$�O�Oq�����- g�\F��t4@-�2"OLRsG��hP@Pl����q�2"O�EY���2�ƌ�MC�ei:$	3"O"�*Ղ�zLtseKN�b6�y�1"O�� ��+�l P�d�x���R�|2�2�=���:h���/\�yЪ�H�[�ԝ�	X�	ݟ��O s��|`aXCލ/5:9"Oj�y֠��%��l��"7X��I�&"O:,p�-_'=�.mxB�AH0�!�U"Ot8uj�8q�V�9��:?�]�V�'*��$K�;r!�4�֓.��1@��r�ўh1�=�'|�І�A�f&��U�lU
��?��z�>�RD�38v�x�U!�4܇�~_��e�a�Ѹ��q��هȓO����Ƈ�}S�X�(ԇE���ȓ(A|����j;ll E�ą[���G
-ڧm��u*P�U+����M?Bg����/X�"<�'�?q����� `� $M��0��,����e0!�DJ<h����cC�w��ȑLl�!�<��mJF��2G���(M�!���bni۱�A4-`�у#�@!�D�?�d�;Cf��x��� ���D��&�HO>���&��]Z�,S3�ML<�r�f�0*�%S�y�n�,R|��	
|�����'��F	�,9�bpn@ �J����;I>)���?����wG�QxD�`�\�+q�����F���`�ƋK=}�r���/E��O�`�c%�������W502˧)ZвC�g,Գ��˫x�(G|�AE�?����ODlQC$��O��!w�UiN�.O0��D_:M
\x%J�(?̕uh��t��}���<y��Z�G��B3#�1�:P����Wy�ڬ�yR�'G����OjeY���[�l�Fe���]X�-�O���&_tX��/��s���)�'Qj\Q(W�Hj5����^�mht9͓Z�f�ٵe�
yx��E`����%�\�
8˗%e��,a�gP��yNC�?���������d�4@��oe�X��M֣`tP4:C�#D��:uNϞ�f�&r,(���;ړR�?�q$
ܿ-�t�h��$
k���K��D�Iܟ�d��?�M;���?������O�����j���p���JN:�8��U�L#�q�I�P뜜��F����g�'�I�C�-CBm�"*�F���h��׮�2���.�ת���ɫRP2�Ɓ<�pس"�"$�<�>{*a�I���F{�:O�(�EGU�s?���ʅ/��i8"O��v�؟Q�j�����?��)8��'Xp"=ͧ�?y/O.�:5��'@�!������ b��rr�xn�� �	ԟ��'��'0�ɋ"⹫΍4Bi~I��)�-t!`a���;3��c����L��� 	��pb7f]>�Ak㤜:2@��D�b�š��/ ��D�b����d.ڸ#d��DI�I
������	G�'�d���D�!*D}� !^�_#����'�lb J� K`y3��R�L��,O��n����'h������~������F6#����'���71�m�vnZ���d�O����O�����&�c1�×��4�܉8���8���QƬы�r�a�&s.J �ج+�Z�sJ|
ӧ��d8 �Qȓ�,-�8Fc�s�'f�4i��?A��Dhݔa���"�^�C��%�"��(��*�O�m�c�(H��䒢 !i<H4c��'ö˓Hm����O�8ZE5	��	~��'Z���h����O蒟<�$�O��â Y*:��K6��R���	]���[���:5'�8u���6o��'��OZ��ks��"yVb���i��GH��'���۔�K�<�VYcc�V=�?�0�O[��!R%̩u�!�F�s����/�O���;?%?�秀 � ���H�c�������
�(Q"O������$e{2�B�x��08B�ɮ�ȟ�hhr�Ϥ{"�`Ɂb�c�]3� �O��$�O�aC!������ݟ���^y��'f`Őr��&#ހ�� ����u�T}i�
2L� �c�<���I�q���@�e�&��=Ӊ��>�@��O�-��^ÐtA�?#<qF��&�R�P2/�Q�^���o~�^��?I��hO��(�FU����1;"����Իb��B�I2.������u�Bt��FQb�h��Oc�����'g�I�p*�Z�
���I9ǯϔqBx則�U�M[���?9����D�O���`>�:��Ha �4��,ߵ��U�W�/�Ԃ�?�0�
ۓr��!�Խ
;ޜ(��GZ�8��%$�,��К�A��eia{����?�S�¨#�Ұ�#F�dlh�Sg�4�?����.�8��C�J�F$�*@.Z<e ,��L�1�gB�2�M�"��EQ^����iR\�@8�'}��R��"�����c~�!�d�˃�H� �Q����?���^KŪ�`�r�Z��O�C��YrQ�՜Q0�qÀ'��6��8	1G*[}$p�i�.�<P���ʉs¶��6g�?Vb�����O���O���l>��/�c���d�;n<j�S���O��$9�)� r��\�9���薁* � 
�i��	�@=����E��L�F��'��S�X��?����?iI~����D?Y��L{�υ6}\�qϖ�Tax��'|�Ov=!��Z����dL5k���P��|��O6�{��d���b�`^�0�$u���I�����\?���`�T>�I�,�E��L���ƉwZ~�IDJNK~�!}Rb���I;�ħI�.<�hT _��H���d�\=�=}�̭�G��'@�-���O�]i�u� N�>�TM���ܲ��I��	<���'���.�Ը���Z ��gU9��<��a�'=hy���M�u��e���M�M������^����_�*��FP�5�6��O�lڕV�h؄���I��<�rF]��v�o&��O��G�T�G?��l���"�A�eh�W���	���ҧ�9O~X����0���C �D�"#��}/�,��&	2X�'@콠�Ox):��Ҩ����d��n4.�
@$��^"�J?��!�@~ʟ�d�#-�����N��C#�&6�1�
�bD��Q؟��Q�W&I�$�4j�"k� ���'D�L�ED4I� MX#,V4��q���dӂ�D0��I��O��禵��m�m�5��8���*Gp���$ ��`��y��M�ë	�>@��B�˅#(Hs7c�^��W���OZN�ч%�!>">x�(Oa)�р�'�v(� ,΍=�|����N<W�,0�
�'cjU�Q{��q�K�H#�'[�eC��ţ,�<JUܡKHx 
�'���as�)l(�ZQ7R�	�'�N�8R��q�TXqI0��	�'�<��g�-��mk �͢F����'z(�����~И{RK�D���S�'�����#��&��G�;C��,��'Q�D��-_�8��3�B�5)U4�X���ON�D�O���O.́�̋C�8(�t̞-@��p�U��柜�Iɟ��	ҟ�������͟H�SB�� �(��B�O6G�<Q���M���?���?����?����?���?!@�2��+S�Q~kȨ�A
%M����'`��'D�'s��'���'�Bg0
ݎ��ʈ�s<�`1%�
6K 6��OX�d�ON��OV�d�O����Oj��Ց;�l��R�j�<BG�I3YqqlZϟ4�	؟ �I矀�������ԟ`�ɉ���MK�\�td�C��\%:���4�?���?q��?����?���?	�i�t�"�"Z�X�Bp8Äѡ���f�i�B�'`��'�"�'���'r�'�^�(�lC�Hj��#*�K&h=�W�oӂ���OJ�d�O<���Od��O��d�Ovl0P��P�d+C��`D ����玲�IП|���d��؟X����p�	ן���I�:}mp�ѳ����كa��M���?���?����?��?����?Ѧ�ζQmdM��I�	.���Z&՛��'Z��'_r�'�R�'FB�'R"��	Q�b�(�lK#|h*��2�M%Et�7��O����O����O����O$���O��^m��t� YYt�#@ $Z�=oZP~��'M�h�O�d�����r"���6A��6lcZ���'��i�Ħ9�_�fd"�$G�?��ݛDټ{�F��I�� Γ��$�)�(��7m��8��c� m�	۵0wi�t/�O���?s�1��|B�'>yR�G��IXѣQ�rZ�ā����D%�$M`�'�?a
� ,��-!8��Zq��[��p����B}��'x"6O��/5+hEb��#q|,Ԛ�G>r�T��?��(�'���������ӱ2O�j�ϭB�s�Y�"M&�H"R���'L2���I̎'��D��ԋ]xN�bK�O�,�'��	��M�"�O@`�Y��Ok3��yBM�"{Դ@d�'I2�'4r�Z�|������̧4,�Ķ�(}����r��؛�LͽC\6}���	ߟ��'�1��(KE�~��8�,0✕��U��O���?	��$�C}�Z�T_6���T/V8ꓪ?���y��i�+ٚ��i��Z͖�@���%M�&�`��'�j��Ăǔ|"Z�41�Q%:�P�FI�"l�f����R���B�O��	���`c��N�}JqPC�W,6�`�$�����?9�]�t�	��0�.X�(���E��`���#.:]9ҤAĦ���?���!N_����3�������.;R���P�G<U��
��ߞN��d�O��D�Oz���O6��,�'t~8��πT�\�����R���O�D�O�'�B�'UV7�,�ɘ_� ���W-wҒ����Dy��O����O��$αwH6M.?��h�> �e�ʠc�(��	�V�4Ic!CD �~ґ|rR�pDx¨���
P�썊��1g���'����?A��?!ϟvH�h��W�r��PD,�t� �\�ڭO��d�O�O�'V�VS�H��*�\�Q+��t-ʱbkũK��]mZ������VY��'V�'�*�B:À	KaE݉������'�J�ă49Y�<�����2��'���U���ܴ��'�2�:��-Q�t��R$d[�l��	���\;M�7������]���'��P���?��?E!��4�����w���� J�Oʓ�?)��?���?i�����PfzA�٣u,Y�E�^�^�8��?����?IO~�Q���>O����C�K VP�@���q�N|�D�'M2�|B���
��N{�v�O�	�HR�H�x�*�]c`��B�'�$=`�K?QK>�,O����O��8Q�Y$k���1����0�Hĺ���O���O��į<aZ��Iߟ��	#q��9�!��Ja&�pb�\�y�@a�?y_���ԟ�$�!���=1�f�Q��k:ڴ!�ddy�F��7��@�Q�i�0�����'���^,_��YY0�Z�N� X��'��'���S�<��ec�A�e���
����A�̟İ�OH�4��f���l J�̌���fs�B�I�����̦��۴L��H�'؛���t2W�V���ߋe_��Nݼ|�vq� �X�&�֠&�d�'���'��'|�'�D�&��{�lu��J00*� �Y�2�Oh��O��$5�i�OHM�Nu@�KT@ԥ��ʓ�OD}�'��|��4��+O,	0��8uT� P)_5A�MB��i���I�v	r(��H'���'��H��N-m�"�����2tk4�'�R�'���'U�Z��®O��d�LJ�	��kT����)�L�/�b�ভ�?q&X�H�����Γ>��<���
P�k� �$@��u��&ŦU�'� YK'�O~�O���(d��4C��X�`�0���^�x�2�'��'���'���n��Y�`L4F�4�� E�X�����Or�dWW}"^>���4ܘ')��'E��&
�L�'�.N�K>����?Q�J�05�ڴ�y2�'jR��1o߮����z��I���".Z�������4����O���Q!~��R�JU�S��<�D�t�s�'P�X�2�O����O���4Ҡ�Q�X�>q�.�Zr(}�B�ny��<����M+�|ʟ|-�E
D�Xl��iQ,��[�hT��W]D�4!�I�����Q�5���O��C��X��go�S�%�¹��'���'�B�'��O�剭�?�0�O>�xQW@P�}�S�Ժ�?����?�7�iw�OH��'�E��8�������ʚa���p�'|��C:?l�6���:��'��ɛ0[����N�T��X�vH����P���	�`��Ɵ��	��X�O�P��N���x!��M
o���Z������H�	_�s� 
�4�y+�J����Y]n`3&AX�/��i�&�O�OD�]���i��$�.��U�Ů�7j���
�.M�)"hܓ]�`�	�@��'��������4(PV\R�Y*��psf���D:�,�Iџ���󟤔'g���?y���?y"ĒȽR�K,e"<9B�����'~��
���wӐ�$�Ѐ�M-"zʬZ0eH�l��ǃ���ɻɆ(
��o||і'��tI�՟���;Oح�֋�4s�,�[�ƭLbz$��'��'q�S�<)P�I<��8��#)��9�G$I��l��O˓Y�6�����ͻ�o
:��8�����S�R�
0��O��oZ��M{�ixj�`G�i_��=�݀e�OR�e{wa�^��M�e��@����@�IKy2�'R��'�'1���f�t4cd�?w�nա��(��	)��d�O����O
����D3J�r���E�j^�19�	�|9�'o��'Lɧ��'"��$N�M��%�KT�kuFW>�:�F�i���]'�8���O��O�˓,,ɱ�E˨� �.Gd]h���?����?���?q(O��'=�� P`Y�� )�&����&�^�rD�'�:7�6�I����O���g��C׌ % d�X �<$��{��64?��Y8�֣|��w���C�qzl�&��o+�h��?����?Q��?�����.��$i�i���׎��>�f|cQ�'��'ʘ��?���Fr����x�����`�q��!�5I�	'q�'�2�'y�ℕu+�6���~�8ŉ��˄q�ɰa��2�~b�|V��Sٟ<��֟\AU�4g �����,�������ߟ��	my�L�>y/O��D=������X*Л��K�uy�>��?9I>��ܽ�@�@2JY�x���(�ؕ��]0	�px"5�iO�ʓ�ڕ��� %��
��.2x8)�t̓ r�3"�ݟ��	ܟ����8%?��'l"���;D�t�A�Y5 ��1j4RQ� ��4��' ��?�$��2�`:��Q9
` t����?���s�@ܴ����B毱?)�O%R��P�O$i
�e@#7�l����d�O��d�OP�$�O~��&� ,'A
.]b"�]=~.�l!�kC��d�O��D�Oܒ�����͓5Dѫ��)�q�F��
(+p�	ݟ�&�p%?xP�즥��b�@���$x�\����)ۜز ���&�t�'��'c
�r���,���ЖᑊO�����'4�'R�Z�X8�O����OX�DF^��uKi�P��틅�\j㟤©O,�d�O��'��k� B�w*`R�jZ�6� ���Cfy�I�i3T4#����4�L�P�2�	7_
�2L^5\Ҁa#V�u<��O����OP�D7ڧ�y2IX����@��.
ًÏ �?�0Y�x��ܟĈܴ��'g�4W]�� ���Z$)����#62�q�Z�nZ�Mې�G��MӘ'rR9gj|��Ѻ;ŋӐ/�*�X���E��r��FH��Sy�'Yb�'U��':�瘚x�H�)��Sd<1`e���)Or%�'U��'�����'��@��l�&$h$z&#�N��� �>�e�i�&6�HC�)��;�n���[�DC�q�QYC�`��c�f�O��hJ>i*O�(ۂ��(O蹚5��7.�`����O�d�O����O����<i�^�x�ɯ|��ݓ�Ri>$�q�C�GU��*�M���O�>I'�i)7����HX��.c��{�N�&,����F�7m!?1���24��9��ݼk�OO�����0閷;����5��0���P�I� �I���F��n��0�9R��F�`噗P��?9��?y�]���Iٟ���4ט'�h��ᬖd(�
�DηC�e���x�'Gr�O�xl:�i�	�l�n�xtxxj kƫ���0��J�F0��g��_y�O�B�'6R�αuQ�X�#ZS��MAP��h���'v����d�O����O\�'}\h�A'�P����'I���'0D��?��4<�ɧ��ɼ3�~�2�Cɉ$Hƫ�6��:��-����O:�����?9�$����rb\M{4$�	���'Z�Z���O���O4��,���<1b�'�v���V�4ji�6���J*B���?A�B��&�D�`}�}�*�A��j�،.��Q�GÐ5,G�nZ;�M����M��O�xr����O|������:$x���N���@`_����'���'���'r�'d�
����(*{-��2��ʹ^U�1�'x��'_���' �7�{��@  #���jJ\�@�g�O��D+�/�	CR;�6͸�\�AK�CQ�!a�͙�\Љ���O� �X�~�|R\��|ᄣʧ ��,;ա�:(68r*�ʟ(�I����	My�.�>����?1��d����ɍ�A�x�*�.[|8Mяbį>���i��7�{�	=fhF�B��������h�>T�P�'�:ܐo�I�PYp���KƟLpW9O�X�̋�<�>�{�+�:ia&Q��'��'���'f�>��taB��&�,v<d@��hm,��	%���<ѡ�i��O�����a�I�!��(\ <c�˅9"d�d�O��d�OD��S``�v���jpN�~R ���a�R�:qL+�� F��'�l�'���'���'1��'��[t�E1Q��QAqO�+10���[�x��O��O<��7�9O�i���9^�N�]/v�aEV}r�'hr�|�O���'.��S�M\ lN�+RNY���=�r/A������,;�J�4��D!���<Y�k�
��X�'UcCF��g�O��?Y��?)���?������\}�'6�)��A�q�����MI�O����u�'N6�3�	��$�O���k�@i�E�=` ��" �ٚft85o�/@60?�q ؼ:Q�|��w-ι�P�K]����=Jq���?���?A���?�����@s�;����H��(̈ڂ�'���'�T����զ��<��6l�N��#���f�:��E�Pd�ß����8s�eM����'��YÑ�M�:|v�@tʽ^f-4胰��������4���d�OX���=��-��-ڝ$s�Ƃ��TE����O��S������	��O���9�f�x��D.ɔb�p�*O4��'�2�'�ɧ��]gT��ׯ��b��DF�4)�tFOF�07�!?���;�	l�I�$q��a�ndK�)�-<����	՟��	��L��L�Sqy!�O� �-�(d)F��7���T�����'��'�N6M0�	�����O�`�D0�c�s_�p	5�O�����Bml7�??���I�c�c?���l9����N�-���B@��O8��?���?A��?����';����d�=.�\ˇ��2*o<들?����?aJ~�_Λ�4OfU3&8Z8�<����2A�N�� �'�2�|����D����O�M���J�el�I�#Α�o��X��'��[��u?	L>y*O��O�-��]�*��a�.[��j���O����O����<�Q�4��ޟ��I��ژs�HQ+�����g�?�bP��Iݟ�&��3b��f\�P�I\}�"��ǈZ]y"B�>q�<-�f�it�i>)���O��I�W�D�B+F !�.��0���J����OH��Op�$<�'�y�ڃ
�6�0DNK<~<>L���?�Q]���'�Z6�&���?݀a\7r �ڀHǧ��qchKџt�	ϟP��sɊ�m�P~r�	�����"LQm�'{�������V�n �Ɣ|�X�4�	��������	ǟx*�D=d�*,Y)��G2h��Sy�f�>����?������<5!�>2"hp�h��F�<(Q C�>!���4��C�)�S�q4��f� 
��qQ��� 4|��$ٖfv�:���`o�O��L>�(O	�j
�X*�8���	N����O����O���O���<QBQ�<���B� ]R�K't�4Ui��о3f>e�	"�Mی�M�>����?ў'��z�C�7l�X�*�+z"���<�M��O�m�G*����4���1�^�[���{g����ʂy��Ղ��'���'���'�'v>�f`�>SS���ߠ3#��/�O����O���'���Mӎy�E�T��t�.W)w�Z]�2������?���?�ĕ+�M+�O뎜�Sj��Asb�&J��{���=o����f��t&�T�'���'�B�'<iv�O� G\��/�V�\��'V"Q��O��d�O���<�Ǎ	WE��7�#O��Ӈ��cy2��>���?yI>���!Z�&�'���A��8 ��A�ǜ�e��lJb�i���?�2��OГO^aʳ��>��	�b^�xN������O^�$�O�d�O����S�rQ���l�^��0��-�?�)OƝn�Q��Z��	Ɵ\�6l�0���@%�z6�P���ݟl��e >9n~~�%L*M$H�~��D�M&�����&[��h`�a�P�'�R�'	r�'���'d��>\��s�̚H�`L0�������'fr�'����'¸6Ml�Li �B)T6�l��FI|��ҵ��Oj��(��+�� @�6m���Y0�T�]���I���&vr�-��ON�����~b�|�V��Ɵ�Zǁ��Ԉs���mq�G����T����D��eyr�>���?��)��,"��:B���jA�T�@�z�#�r�>!��iDN7��u�	�1m��!��:3E���5�C62���'��x�-+��4c�O�阞�?9��o��R���	5��!�K�S%�Z�2�'���'*"���<� �4OX h+�$�C��L���Z���s�O��D�ON�lZ|������ןm��+%g"(Qv1�Q��?����?� �i!>�ói���O�@	Dʳ��]w�@L3#�T�e�"�\�E�m�O>�*O��D�OF���O<�$�O��*�����Xy0R�ۡ&.� �<q�R��������k���l�vg�m1�� ��K�ZMX�8��dCɦ�ܴʉ��O���S���h+�݋�n�{�<���.��$��O�U��_��?1G%�d�<Y!�C�P��nH�\nv����"�?���?���?�����W}��'���e�����P� ��-�#E�?��i��O���'�2�'��dQ�z J	�#���CLA5z"��ó�i���1��J$�O�q�(��%HFT4ɜt�(�z2 ����D�O��$�O>���O8��/§>�B �ŝ!z�V�rFb�A,ty�	�4�I!����O����1�<QR�]�h��lyw�^zJ
CM�����ll�T���'E>6??y��U;=����ƃJ�Hk�!I�"��	�C�Ot<�L>,O���O��d�O�dؤ�������dA�K�2���.�O����<�X�X��ٟ��	g�ĀD>X/�L���$G;����#�
��$�T}��'<��|�Od��>&�n�jd���D�Y�Mf�Tcb-��������6T��$4�$�!)��㔎��F�_(A|���Oj�d�O���*�	�<�s�'aP��E��T\ah�W
l��ݠ���?q�hr����\}B�'?D�⠅�0U2� ݳ,0��sg�'�)�->H��?O��d
~4�L?牔�� �0KR*F#�5P�k]0@����By��'��'Q��'W2�?�Ц�J�.�̚�^x�x=Rto@E}2�'�r�''��5nZ�<��EEl� ���82PlX������	P�ڟ0�	���H��̓ J`�)�L�-�c��8(�-��A�ẟd$�������'p
=A��E�c�2h����QUJ�B@�'2�'�rP�@�O��d�O~���ip�MI2ύ�p�x�Bsj԰%�P���OFHm���M���x2��-��L��M�����K#@B��'�d�3���D���O&�iЩ�?abh�܁�C��6<��/�}���e��O���O���O6�}Ҟ�� :t��Z+U���QWNКό���'b����d�Ǧ��?���1�,�c��у#kb,�v��dU��b�?�vLmӠUoZ�3lnU~B��9֬`��$zL4��DJ/.h��ֳxU�����|"\���	ߟ��	��H�I�$� �E�-�lsB�2e�
��sy�ϯ>)OB��;��>K|�-�'TMFxc"�F:]�x᢬O�<l���M[��x������J�l�����U��	��B��@t�	�&�X �'��%��'~N�i�q��$�����b�'�"�'���'��Z�b�O���yl\}daI��!�c
9�p��^Ǧ%�?�Q��K�4囦C�Oƍ�#cÓ0L������Nz���^:y���(���Zp$��$�Q�ʼ�HX��蕥Ylڅµ�ȟP�	ޟh�I����	Ɵ�E���ΰR%�(y f��3a��$"]!�?1��?!U��	�d۴��'|����aۮGgZhA�`�&��	�O>A��?��W3v��4����x��b�Y����k_#Y��5�G�{��I\��|y�'���'�r�o3̩���s��9bG�w��'������O��$�O��)�.L��덺.�:���X��'����?����S�)F4��b ���7XҼ*1fΤ`�b�A#��ݛ��<�'O�d�IV�I����Ѣ���,��������Ο4�	�(�	\�Sxy"��Ox��wG8	���Q�~1�)��'u�I(�M��r�>�ջi5� ��!���3ͅ�1,Naؐ�j�6�oZn�Ftn�p~�a+��Ӫ1&��=�ݙE�xILmh��7H���<9��?9���?Y���?)˟ƹ�FW�G�t���G`+�m�To�>���?9�����<郾i��D�=\�!j�a�!|����5`T�p��6���a�N<��'�R��1v\}bڴ�y¥Yz�:��W-Y�X�28�e,�X�����ʔ9�i�O���?!�f��ŻP�(3�`��H�[^�x9���?���?/O��'}��y'%�C:%�m%5{,M2�<��O�)�'���is(�O�	���?���XQJ���RtJ'�'�2˘�jJ���,ť���������NI牓bK��[�:��<���������Oj���O ��-ڧ�yR�4 �c��**<�s�H
�?�AP�T�'��6�'���?��ׂΩvb-0�X�`��E柜�	�H���	�� o�<Y�� *����~�T-ذ6~p��.&X!mf�Py��'�R�'[�'�R�Ğ ��PK��9ia��+�Y6*~��:��D�<�����'�?y�dN�o������5����o-"H�	�MS�i��O1�����%aY� ҩ�<<��$K�N�(z�HP.H�	�d�I
5�'���%�L�'z��2BEr|�!JD�M �N����'��'b�'f�S���O��$� n&}`�aI�/Vz�(�fQ>j�X��YǦ	�?��Q��ٴ%��F�O�a7$W�#~B��Q����q ��[.U�v���)vTiD�4�)b��v��g2؉q��3f�ȌCP��O��d�O��d�O��d�O�#|b�l�X���r� \Kf�5%������ퟤ��O��d�OԱn�J̓EJ����@:G%�)� Y�"���IL>�ݴ8F���Ox���лiB�$�O�,��gGZ��1sӃB1	N�B��D����2=*�O��|����?��s� @[ #ԏ.Lhp�l 5�T��?)*O���'Z�����OL���H�V�DT��!_?~��-O���'��'�ɧ�ӀBB�D�UM�(��M�F��1�F�&d��x�.��R�����?��Fy�Ʌy���b��c�]	WHO-�	���'���'�"�'��O��ɷ�?9�E��4���2��@��ğ0�'�X6�"��0���Ot�v�Bc�"�ʅ�,Fv�j�B�O(��!u�7�:?�;T�<���O���5�j���Oq�T��DG�� GZ��<Y���?���?���?aɟ���@�Y�PH�gi�g�ꥒU��>����?�����<u�i���׈Xu 𚔧C;M�I
��Ӕ-�R�'z�'��Os�a���i����(U6��
�$�hNµ�be��Q����������O�d��H�pC��,A��r�U�#����Ov���O�j
�	�������A��b1T�7N�	~j���f��4�����IL�"X|�'�Er)��3Ԃ9�$)�'2�����sS�&C0����~�8O�XJSꜳ nP�rC�ܓ/?�MC�'���'���'��>E�qO\�7ƒ��T�w�Y�$��I�I	����O�������?��� �ٳ������i��kR��ޟl�Iߟt���+6Έl�v~Zw��crߟ&�����L�*e#�)�*l���8���<1���?i��?I��?9Q��iP<�J�" ��n%���'�b��?���?QN~���=I���M	�!�у�FI6=���T���	���%�b>�X��ъ�|�EĈ�,X�b�Eqndm���`�(��'��'W��7|�`Hp�ޚ����&E
Y�"h��՟��I՟��Iҟ�'w�듦?rL��=�����C�'�ze�� ��?!�i1�O���'��'.�D�mL&�)d�/T� �
���[� 8�t�i%�	
N�n9��ݟ<�����Z����l A� N)�.���O@�D�O����O��+�g�? h�%ݸzc�@��S*ʸL���'Q��'r\���ߦ��<)��Ŏ
�ڙ� �6N�@m�SM�j�ޟ8������'�ΦΓ�?U��R�[���� ���@�!���0�饟 $�������'�'_B4��k�*nYK�e�1vD�qiu�'��W��ɮO���?aʟ �&�
k�N��tK�'v���� Z��+�O���O֒O� ���E,�A�h�����Ja��/W���ne~"�O�^����N�j1z!ė�m@�X��P�$t����?���?-�M�M~b*O*-�I�(b`��E��R�|�GH�g�H�$�<	�iK�On�'��$�=P�-�4b�]S$C�,��'��X���i*�ɫGi�A�	D�r�p8����.^c�)r�aE�H��Z���	ɟ����p�Iן<�Oh��3� �~,�I0��P'��9�U���'2�	�禕ϓkD���D�_,i��<�D���86��	���&��'?A�I֦��Cl|s�Z.+�9z��2<���	0G�e���O��O4��|��C�|�	�f
�9�� �)���Hy��?���?�*O�|�']��'cbgJ
G25٤e�
_����C4`�O�t�'�07M��uYH<9RaR��Lh����vd6��������3����L Ȇ�������"Ȑ�I�y�ax�D_p5�ၣ��V���O���O��D.ڧ�y���m!�	��)�PL�yp+���?�Q���'G�6-?�I�?�w�$��K2��3lՋ�A�ԟ@�ٴPH��gc�0sGf�x�?R�Z'��DqҶ��kv�(B�G�0تl��
_������O����O��d�O.�dҕd��hh��~���CTe�I�(ʓ2N�I��\�Iߟ %?�ɉ�h���BΞj_R|a�f̬KR��[�O�Qoڷ�M�U�x�Ot���O��u�(Ӂ)U��y5��Y HƇ�2	�4R��xRnA�r J�	gy��P�\�l��ӃW@�`c+��F�r�'���'���'�������OVm��b�*#hH��8Q��L �G�OȤn�L���	���I�<-U�N(S��>Y�q@K��%k�����h�
����T�i��}y2�Ow󮞨&\ ��nC3���3R&�[Yb�'�2�'M��'.�ᓫ\��A�Pi�^��\�S'/I"���?r^������4�ٴ��'�>�� E�]6�:������M>9��?��K�,q�޴�����ؐ�9NvZ\����'&��0C��

 ��I^�IDy��'s��'.�ͻV��&j��}/@y�$Ş?]�'��	����O����O��''��$8!�C�4u֍�Ы�s�(�'����?Q���S��� IK���c�u`uأ��^����./�����<��'m�t�	E�ɷ.6��:��B�D���X �Gנ5������	ԟ���|�SFyZ���1[0�;�,cQ��K"�'��a�b�dp�O~�D
�>�����-
�*T�F"����D�O:��hn��Ӻ���K���?���ފ'��X�CE�xL�m2���O�˓�?a���?y���?!����ְ16�d��i�?�b ��X���?����?�O~���S���?O�愋�� t@rN��=� ���'��/ �d?�I�t]v7M��:��"-��򂨞*k<�tI N�O����BX��?��-���<ͧ�?Q"���8VX۶��7f�"j���?����?�����DB}2�'Vr�'�m�f��*K��M@夝�h9��YP��MW}b�'_b�=���nМ����MRg([
���wo�`& A�Xu6�����ßP(1<O�E�Ӧ¼F�h��Փ�����'xB�'���'��>�Γxg:L����'A�`�X Ě��8������O��������?����A�&#�� ���1k��&
�9���?	�����3,Y���А�GU�����D1���=sԊ�Ud�n8�D��|bT�x�I�d��ܟ���ʟP+��п(���aOE�V�|P�doWAy2��>����?������<IU�����OV��F��`��27��$�M�ihO1�8�kw��?"�aǊ1{P<x��I�_�҈��i�<�X$4M���'>A&�P�'�f�h���Q�a
�/.kd<ѐ�'��'���'EB\��k�O���x���^7@D�m�%��5�������?�bX����۟0�{�b����L�q���w�����J���'/���f�c�O�� >4ڍp$UJ�鑃S�AR�'\"�'$��'(R�F��t\�M�^�$���w/��$�O���PL}�V��ZٴƘ'Q��"��HJjQ)���6�N>i���?��?%ְ�۴�y��'ˢ�"uH*_��4[�+�iy�I�^L�8��䓤�4�*���O��dA6i��T�f���WkH�!Q�������O�ʓ.��	ܟH�I���OW�ͨEă3\X��T�/>�T��.Obx�'��'�ɧ��m�ཙ@'_�)�f�����w%�Ы�/��{:(7��Ny"�O������O���˴eD:t/:rW��)�e���?����?�������� ��,l%�͒���)�4���O`˓]����W}B�'�"#�q��`	�D�"�>0��'�-�"p/�V>OD���q��h�'��$�N�P�6e��n��'��D�P��<���?I��?���?Iȟ� FiH1�X�ck�a5�޲Dr�(�c�>y��?�����'�?q��i��%1��p�H
3Bp @##�B��'��'8r�'��a "8]�F2Ob��E9?�P�S�ġU�`E���OX��@��.�~��|rZ����͟���x3��W$� ��Kp�DƟD�	蟘�	ny2#�>!+O*�:�4Y�$���~�x�^�[�&⟘z�O�]m��M��x��B�a�@�� _)���S��I�|���r�H��C1�'?�j��'4�ϓ.p9Ҁ*�3NXtj��ݙ"��������	����m�O��@�v\x}�"�܀�\s�J�?�b��>,Ol�_����s�uL����K
kT0ȣ��;�?Q���?��aŬ�{�4��D�=�l��'�b� �.2��,���\�E���2�)�ļ<y���?����?���?�W�W�M��=�(D�@���)�"��n}��'��'��O��LB�5�N���)]�|p��I�EG6b� ��?����S�'B��}ȁ�8�&,�Pf�7��|��6�M3�O���]��~�|�^��YsO��o("a�O��ɄM{���X�	�(������	py���>��bp���kW	2h���r���j��X����D�o}�'[20ODI��MUv�e�ܯ7�X�K���Uy�����c-]RQ>��;r�����/��`$N ��(y�I��P�	۟��Iԟ���R�O����Aa�!Z=�mC|�
����p����ĭ<1�im1OzM $�ɇi�d,�@Ñ�!��|���|B�'���'e~źƸi��I�^C �֭�,6)���%A�_��P�Ͷa�2��n��wy�O��'�¯l������s�E=Ӕ�����?�)Oȑ�'�R�'�?Ys6�?T�[0@�0d*�Φ<��^�0����d$��OnH�T�����ION�:憎���&�[P~R�O3����� ��'7���&M�r6�9ʗ
M��5���'���'���'��O��	%�?)���5D�uR`�ײr�2��U�󟨕'��7�.�ɱ����O�
7��2��X�$��� A��OR��#X�7)?Y��*i ���&�� ��,9k�j�?�X$8�,֥�b_�������I�4������Ow��r��E�pH`h(����p�R�CwT���	���p�s���4�yRa�h� �a� 	m��:W��2�?������}����4�~���2KY�kY0`�zE��?9�D�~����+����4�����'n6�Iq/�O~�8jP�P�Eb�D�O��d�O:�tX�I̟|�Iϟ C�Ɨvv���&׊9�`�����a��0����M���i)�O�@��#ϻv�bV�]�2�@\���<���J���4�r->��'������y�E�s� <���;VTh3�ȃ�?���?����?	���o�pr1(�' �N���兎q�:�kGG�OB��'-�	�M�b�O#��u���
`�wO�����&�''J6-H̦���4*$�[ܴ�yR�'�A��o��?����U8��]F��G�0X��┲r�'��	�������͟��,2!��o�6J"s����R�T�'���?	��?II~�ՄQ@GJE�5��A�Kӧr1�!�w]�,��4d��vn&��IO$�&o˽{��S�Hv��ypKkR�� q�+�!�O�I�J>/O�D�գ�[��j�BC�c��S�o�O���O���O��d�<�^���I�b3	HLP�U�i���1Q��m�I��M�� �>����?��'� $W2J�
G�SU�\P	��)�MK�OR�BB�a�E��2�:�C�L�>tb�Bs��n�=#��'2�'�b�'D��'9>�)�A|3N�;Ê�D�.M2��O`�d�O^M�'�I��Ms�yB��>���s�x�f�����>v�'�7�NϦY����J l�<��tJS��4,��̓�JY0�8��k�u���ͼ�����O���O��DI�2j
�A�S�Kl�,y��="l�D�O˓Z��IΟ8��ӟt�O�l�wi]U|]��mJ-<
��P-O���'8��'�ɧ�S?=��$7H[`�B�æ��f����B�YR�N7M*?A�'aN�	h�	07�8�b���k8��Bd	 �B��	�����	n�Sby���O ua�֌B��P���#KꠌcE�'�B�'D6<�������O�Ճ�Kу]I�A�� �8Lj�Ɔ�O���%[(�6�=?��R�#B�c?q�5��{�.|T� e��� �c�O���?��?Y��?�����I� ����V�ղ<ښ��`I?����?���?�L~�,I�9O�����C�,0���_5p���S�'���|R�����nܛ6�OzD�f��&�����+ИX�
!a��'$�j�]������|�Z��SПx@[�
T"-s2�-7l��¡���@�I�����ey"��>i���?y�.�#�l��������s�]h��>!���?�O>!����\�z�QD^����u��$�O� �D�ޡ?�@1;����S9Cz�
��<!��E�(4�0Ջ�r˶��4)��\�I̟(��͟�G�d=Ot�����zL؛�ꀛm+�	v�'>������?Y���
�Òn��f  � �jѱ^_(D��?i��?���M��O��v,���z\w��M��԰R��F���R�O>�.O��d�Or���On��O
� &1���\��Up lָ����]�8�O���O��d=�9OZ@xTA2r�Y�!�.���P�D}2�'���|���;P��`wON�Frx YE��=��!�iL�ɅV�|�O�O0˓{�E�ł��>��I�FW�f�x��?����?A���?�,O�Q�'N�7{���d�(9 �t��
$WC�o�`�tҫO��d�O�扬� ��G�
���ti�d|jeq�hp���4;\�10k'�'�yW�ϊT�\eQ1l�? \��u�vc��'5�'���'���Ӏ!3 �Ss"�52��
��&SB�d�OP�N`}R�ܡ�4��'ќݰu��y|!��,w�|�bM>���?9��^j�z�4���T4T7*��	��w,$p )̞z��J��O��~2�|�W��Sן���џ�ӆEoh�A���ړϾ����ݟp�I]y�E�>���?1����3$�"�Z��X		:Ti��܆I�I����O�d?��~��1�Ԉ�c낞 q�R�(L�!.��s'�٦ݒ+O�I��~��|���uR�y*��rF�p�O����'Y��'"��P�@��rH�P �H!'^�ӒgY�!�T��IEy"k�:㟐ӪO����=h�L��E�>�t�dbQo�f���O�M±�w��+S�e��F/�S�NVH���Įs�R|�`��b
����<A���?���?i��?�Ο�����'�̉(��Ŋf��HRcJ�>���?������<)V�i���^�|Qp؉�#nVn��(¾[��'2�'q��'t��
*�v1O��H�E. ��I�@f��DȨ[A$�O�2�؄�~R�|"\����X�OJ:G��8S�J�>Bx��A'G ����I�����[yȷ>����?y��S�x���>r�4���7M̕��̣>���?�L>�7c߄B���j�*�V��q�.����Ѫ#`X���.y����|2eN���ϓ0��!č.[ꨅbUO�0C�ru�I۟d��퟈��j�O��D��^f���A�pcd���K'��>9��?i�iD�Ov���u�� ��(5�ԉ�����2�(�$�O��$�OrL��sӆ�Ӻ� Ҽ��� �-�<9��인*�B� oJ �'��I��0����x����l�	�@��Xa�E�: \�Ȣ�[9Q(�8�'�`��?a��?��`I�]X�����=m�hq���8I���?�����O:  &-�B�2�Wa�&bLt�7��^^E �O8�oĵ�?�@">��<���5WD>�A��T&$�6ݚuf���?����?���?�����$Nj}"�'��8AܤH��	���i�p����'��7�?�	>���O��dq��y��a��Y3��L9�y��C~+<7�&?	�A��>dT�)9�Sۼ�EˮX��RtfD�TSD�r ��ӟ����T�I�8�	��G�4OW8<�؄!�-l\ɚB���?����?��U���'�46-/�I�O%&|hG#�E�qwٱ �
�O���O��:7W*76?�Y�,�3����Ex`�i�،��Aa�O<�SL>-O��O.��O��5o�J<L`�!H�l�$�@N�Ov��<)�[���	ϟ(�IA�t�˿q!���a@=l�`G/ ��A} ~���nں��S�i޾�J���"ǀN@a��Lo�<�ӡ�	ktB�HГ�l�S��2�GP�	�94�T-��A����:Q��}�	˟����(�	L�S`y"a�Ov�F�!.jC� :6ǲ��''��'P78�����O���$I�z�S��U�@kӐo�a>�m`~�d�?I�|��ST��+~�j�nD9Gǘ}��%��;��d�<i��?���?)��?yȟ���NQ�Xx໶��2�F]�P��>����?����'�?q�i���
�e�8V��u'6^O�ֵi��6�z��_�Su�N�lZy?ђ�21�� 1�)ߠ>C�Y0$�4SC�B���e�IVy�O���Ҹ#k��u�ۅ^I|A���:|�'�"�'~���$�<���+�0X3dI_�B���[��e�X���)�>1s�ie7mPs�i�u9�ix��yӎL#.��Q2T��aC�|yZX��F=?�'7�����:�y"E�{-ҷ��|EY��?���?���?Y�������w�\��ʣK ����b�'����?Y��5y�V��矊�pc�
�� q�<rԝ���j�������ߴ&mL)0�4��� �Tr���'�uw�_�Uܦ�+c��sw4�JH�&������O ���O���O��D��(����f�d�ڦ��2�f�E<�	�����㟈&?����C�X��!Y�e�-����I��*�O�%oڪ�M��x��$��.F)��P�C�[�<)��
B��r+����$�	������OʓjxJ�B6gߕ_X&@J�a	]0�t@���?����?���?A,O���'��Ȑ��(�[��h�&l-��X��'�,6�/�I#��$�Ħ)����'
����$I�C*����Ʃ?�v����Y��M��O��M���47���ЀW��´i����S�B==��'r�'T��'=b��-7�zX�o��T�nٰ&7U�J�$�O��A}b�'8Rf�*c��y��<ZP�@�a�bCr4�V"�d�O��c�0�w�v�x�4��G�6��T�aF=j���i ͐�p�~��h��xy�O���'��� @�Ҷ��Ms8̂���~�Ӧ�'�"R�(z�O���?a͟�MJ�ٱz�X
���?�n��[��r�OF�$�O��O�')8�e�Ϝ�W�V�{�O�"^Qb��b�X�-n�B~��O{n����?�l�PV�Ӥ��#6'\&�l����?���?������DW��:�Չ-k]��߳6��1�F�OP���OD5o�~�z��	ğ�����Q��U��k�$=�&��Qʈݟ��	���l�l~Zw��i��۟��'`@V%�1G�*}6�-pN���젉&Wg,�2�ߧ�|�h M�rf��E� i����M��Ɯ ɧR!�ꡠD'�6������~��p��ͥbD��� 4}�ى��ȶ��X%e�t���Hvb�Q�s� �#��lR���sĉ�[[*1��)�*"���!�%�{6�)f�$��|�3K�Xn
lѦ!��hvѠb+� 6��y3�,fؓl��=ư�W�=�� �U�7��ɻ���%j�;��6�o��!��B��)�Vx	�柪 S.ꒈM-d����Ͽ:t���rd@�$��d"w�]*�K䚠4k^�*�J#x;�%A2
M;¬�Vc8؅��(�v����Z<1��׈r�`t���Y�����a�+ݲ|�G�E�$z�x��J)[�̘f�0�*c�E���Qc�?���	ŎN6\xB�&�6z`�h`��d�Q T&~}*M b��5�a��Qt(��%�*B(�b��4i��A��ڲ��ԮE2@A����o��=rBx�0���O����Ox�'3���|�<���%	�~�h�q��'s�~��?��h\��?9��?c��A~����i~������?��?��W��'���|2��ۜ�)!�Ú$f��᭐-#��	!^ބ$���	ן���w����>���Qd@��Y�2��L٭�?�Y�ؖ'�b�|��'��H������,�T���lK�C��e�!�'������I͟x'?}�'Co�J"-ʷ���3f%�e��L�	�l�Iޟ�%�h�	ޟ�����[�DA6P\�x����Dv�i��`y��'"��'��O���?��i��W�u"��I�+��Y���<q�����?y�KS�5��y�b�=(0��wNR/(�HL��GR(�?	��?�*O��d�J�T�']B�'[fds�B�U�J� "�T�Tt:آ�]���П����Z6�����{>ٰĮi��\��]����g��O(��?����?����?����򤒧f�"%�f�`�V}�Emġ	�4��O��(2�D��>yكc��^74�R�׀dC0�p%��O��D��i�	ǟ��� �O2�%�ء1X�>g���$r�Ah����Fxr���O���ڵR[d�23gZ*}�ʄ"m�����͟H�I���	�Of��?��'�"rAG	nPhP6皞�F�Q��"E���'���'���,�2���l
T��]/p�p9�'���'7����D�O(�O�q�aGC�^�̫4��1��� �<ɇ���?�+OT���O���/� ��"[^9�⠆+E>�1W��؟)�OV˓�?K>���?yg���$6�H�*<�5`2 ��f����H>���?����������Aq��Elkz��@O_��?))O���&���O���X�ʰ��#H��e�e��I���� �>�ʓ�?q��?�J~u���l:��k3��?}�\`�N�>8B�'��'9�i>��Ip�D�!W 1�u�n���hC�8�?����?�.OD�DU��۟��;����Fƞ<]�$��!|�Ν&� �'�"�'V��y���`qJ!�V����b
�C��^����%�M[/�����O�L�'a����d��A�N�% �e$,x������O��>�	4��J��ҥ�ĝ�x��G[�=�˓�?���?����?!*O�:&�}1hZ=�ܔ�!@�A�V��'
`����Ӻk�8�i�N�x͓U�.�4��՟��	����	CyʟZ�3�ȵ�j͞F��1õ�ύaPf�f#��Oy�6O����ӬF%���A�,M��Y��':b�'��	P�t��0O��q�
bAA\�\����P &���"#]1O����<��'��b�
�[}�)�����Ƶ�������O@��?�Iȟ��P�>��@W�c���SԫA�4p���q��?Q���?�L~�0�Or2t����<1��=���S(g�\1/O���O��O���|B��l8 �w�:�P
���2J�p8O>����D�</���$ޝ���YbA��O[����ѹ(K���%��񟴔'%:��K��r��'S�&�7�[ Y��a���OH�d�<	/O�˧�?����yW$Ϊ,�x��akۻ9D��M ����?�/OL���I�D^�8�mI�^A������!Q��cy��'X6��|Z���?Y�R���랸\Q��2���ۼ52&�O���?����'��{̾��!�	$�l�e�>a�D�s���?Ǽi�2�'OR�'
�O��
1�6���ɯ!��8`4KC�0��'b�'�ɧ����j�(2�& �냸C�0��Ӏ����	Ɵ�����ԗ���4?�6����Ff��oK�5�aoN1<N"<�I~����?���I�<a�F�?e�`M:�J1?�@*���?Q�������!��Q<cb$dx���1@�L�L	]SH�O��$�<���?�����W�~t�D�d�E�{Q��C)?q(�d�Ob��3�D�<�� bhw�ݝM����%��q�R\��'�]�|��ޟ��It�S*��S��*
�HRa��o��'Ly�'�R�|Y��ǟ! 	��Zؒ�k߮<�����O�Ky��'�r�'/�OS��'�?m%O�d��6�F1	���?������OV���Ovh����擿b�,�i��;D�q@)B�(^�4��ȟ��I]yB�'�\맾?���?)��Oa�P��� @2�t�
���O���O � �;O��d�<�;\&��e��-�p%�1�Ԝc�V��I\y2�'̈7��O����O&���q}g��S�ТAo^<:���Ȓ@�8M`��'����6��ģ<Q���nL�J
���%F�������D�?��WX�f�'�r�'tbe�>�/O*��p�B�2J`�1f���u!��@g)�O���45O��<����'Z����B�v�V8R`��{�d�Hׇ~�����O��O
��'��I�X�Ft:���� [r���*�6)���	ɟ�'���Ce��$�'�B�'#t3ǣV�r!W��`�]��'=��'�>ꓻ�$�O���y��B��V�ʥX�`K�e� ���'k�I�'����Ib�'g���Ŋ�$]*(kf��C�L������D�<Q����d�O��d�O@��P��-�VM�f����>����� ��$�<)���?y��� �db\��Z�6IR�DS�Y����?(O���<	��?I��tU� E�ŉq�]������,��!�	ܟ���IBy�OA��g���%D��`2�U)Y��L�k@�����Oy"�'�b�'J�9�Ο�牰4��
�HQ�g)fT;1�mD���Or�D�<��7���ΟD����X*"�W�@���P2ɇg����#Cy�'#r�'���'#�'�C36�3V�T�Ya'�Y�B�rS������M����?���?1�\����@��h0haAj_�G:�d�������֟d�b���IQy��	LS�aR$CE�h��M*.�+�R�'�R6m�O����O��ĆJ}^��h�ΜBv��� ��NI��l���q�.���O�RF�_o�j�E�&l�$MKC_�7m�O��$�O���x}�U���	�<9��x�$�bg.Q4��'G$�'�bˁ
	�O��'0 δJ/x��C���Pi� �8���'d�,���O
�0���vR\V!x ��mU�#˓a���<a���?y���ɔ$Ir�<3�`��!�ԯN����E�'���'��'���'h�"U�)v(�!�x86��w"ɂW$�R���	ğP��J��3���DA���XqQ�G��x�	XFyB�'R�|R�'Lր�~҉K'%�f`���1-(�ʐ逫����O�d�OX��d�$>-�bO��snQ���zV�P����,��U���(�	�-n�e�IL~�+��=��HɣC�#(�
�������?9���?�*O��dRa����H��d���&�р6^�5IB���L$�0�I�� ��E�$�H���̈ .U��BO�<�2aP���O�ʓ�?���i�����\��1��d��O�Te�����M.r4b��ʀo��'�rc��y2�|��ɓzviq7�M7BOI�%3N���'��6-�O����O>���[�I���	1��Ek\��Hʫh�,�$���`��ܟ�&������T��S`�"�p����.#b�LJ��iK��'9b�'�2Ox���O��H�Ra�@B�w^~ƤL���5�ą�S��<���?i�w_�F@+&���8O@�H! ���?a��O�'���'��'��3�	�O���p���,TH$�_���HI�X�'U�'�r�?ہ��?kZ�hr��9Za�4��OH��>������?���1S6R�BD�.Ԕ���L]:�����<�*O>�$�OH��+��B�?ə BR�.<`���ƚ� �<����?�H>���?��,��<�����3��y�3J��N2>�+��;����ON���O���$>�����C@֤*��ޤ�����d���	n����		���{~R#ڽ9��
M�Ggf��&�ո�?��?q,O��d�v�����ɘ �Bd�2�hH�E�Z9OW�e'�L�	������<'�`�'$��PBPCó]"B5�b�Z2
q�Iey��'1.6��|r��?�FQ��6C3��@k�'��=��"�<�+O��<�)��@""�T
��"�V\Y�V�?������'
��'1/1�4����A��O�6����\�q�6��<�������O��M�,�J�����pp���P�^���'��	�`�	���'��8O4�l[.1�<�z�%I��<�b���O�������O4�$�%�f,�VA��pG� +n���O��D�A}����'�I�
�nm1½�EN�$p��@#�<9�ʦ���?���?����D[c��"�a,*�6,�XN��	uy�'B�'��'R6O���QhH/�N�C�	n"��'zx	��O ���OF���Ob�'��ĭs*�{a�Չ%���-��?A��?Q��䓖?Y)O��4�R�2UyѦU�#1��b���ʓ�?���?�K~r'Z?��I%Q�5��În�6�K'$[.��H�Iӟ`�I��6��y
� ԙa���hBAN�8${�l�5�'���'���'�B�'��'y��'���E�9vK�MA�B�\m(MK��|��'l�ɺ_&"<��GV1��Sr �4�x�ɷ� (|hٰ���=#
�t����vbP`�
,��C�'�u�g�����(.�8�/k�a@�j�-�ēOV�d~�|�oڋ�?����?�����
T%�%�]�\�R�F;`��?��K�lM��!BT�CDfu�iE���!�6l5X%ۯ*����%�'K*Y;7������JBR��(q"��I��\8�ֵ�8a@��	3ڹz��͂9�H��AD�Da>Hp֡ %eZ!����6	l���g�m	"h�`��2�0ʳڀ�5���S�
_��[fI�	NΕ�f	#9�{*'	�̡;�eQ�]�����	���3�O�56>u{�Q8:�,1%�|���Ȍr:X�VH��yg����BϞ0���X�N�\�n�x��4s]ؐ���:@�ӥN@z@m�ğ�lZ+x��`�VP�1c�HBJn������H��;a��	�b1w*�Z��$�`G�,+����0��hA�!�Y�P�k��]�
SLC�{��E��EK
\�1�TF�=/k����P��dQ�22�'��)���>���>�8�)SČ�!��y�ъY�<Io�>˺0r��JFrp���
W�'��~J1I�5��8"Gΐ�q�<�h��S?���?A�F��$?�6�'�B�'X��	�h�Ia�
�$E���`�&ѳN�r�}o΍��a�����'��) �Eͷ#h|8�����`	������	W��i�Gh�3�I��sdn�\�(G�ˊ"%��Oڵ�!�'-����	��"F}��'@H�n)���$"Od�{G�R9[��]�!�0,�~8z��O4$Ezʟ�˓l���w�� � ��N�S�ҁ�e�I8y���'Wr�'��I�����|���&l��G2u��l�A����hq$cʡbQ��Z��B=��<���;U?���	1cn�A�/�r����Sa+,I�:%  ���<�ca�)���ʂF���Ф��'W2#e/�2�?���7ғ8P�
U��!䒨�&�#a0���aւ�;"�νe����Q,G�̚,�O��'��I*A�Z�ٴ�?����M��!C< iH�ؑ�7H����t��O�I����hX�Iß'��n]91��1�)D�z��ȫe呟�dN��Y��sŭ���鉝mQ�4KQ�� )Ð�b��߯gǑ�`�r��O��$^K���\;��z�(���RשJȾ��I�?E���@5rD�A��$[���8I�V6���ذ�)§'Ǜּi������E0����ᑡA�&�p���<�㡓�e���'�ҟ���'ћ�&UZ��C��]Qv03SB�)Th��
�C���HWb�* 
C�ԗ68|p��O:�O������9Ct�%�K�o�A��Od}0A�I7:+�4�)V&t��I��aQ ت`3�e�����)��d�䝅Y�6y ��F��$�, �	#�M+�i������O����	�t��=�1m3�xu�W�i�N���O���)lO��֭ضw��Q#��������ɒ�M[��ir1��u��dE�u�LU�F@��iq?	���t;�+�7�r�"&�G�}�%�ȓ!��P�����K�.��ҫ]#PZ��a�lΖk���tS<��=!�eZ���ŮH`YP1�'�Gi�<	�홚K%��c�+�;	�h�[�EOa�<Q�ԭL���Iޮt)\�v�GK�<Y�.��Y�T�a�i(D��̸�&�F�<q��F�0D�t��e�*&?�HX2"|�<�����{��,9w� ?=ܑ�f�t�<1e���!���2��5V��x*��j�<�AH������9���\�<9rI��M��Y�n�5��Q� CX�<�$*�+1�x�ʓ�Xk�B���a@W�<GdX�<���c% ;1��I��O�<d���bļQPIY7���I�N�<�J��f�X���1Di�%�Sj�Q�<�"��b�Εa�Ŕ3�6H�̚S�<��]"���C��e�N�+��U�<�S��yRy��@W��qB!
[�<���ҳcm�` 7�
�4T����Iz�<��ꕚ/�|�!�8in2���R�<�æ�=~��j���\
���A+�q�<�S���LY�ћ�hZ75w\�B�#�@�<	tN!P�, (�'	�����H�x�<9D���"�@ 
e�i(�倳	�y�<yr]�co�E+У�.�qp`��q�<���-2H��`�;E�X��5St�<� �I�����rNf�]�P���QB"O�M���4P�>�@W�L���s"O��rB	�(8v���n^y�����"O�壠�}�ZP�Q�H-�B"O�E�`�D5�h�K�d%��"O���dHޞP|l��l��ZG�eJ6"O�6i�
a�@�1�$�E).D�� ㌊]7!���O8f<�%a D�hȧ�A9/��ʳ�=4���!D�XUϖ����а��:w$����(2D�p�"3Cf|�gO29��� ��,D���pd�f2�9��Ɍ2.��h+D�|��+ܠ^ܝ��HF�k��];�m)D�,��f� Ȍ9A&C[�d�ʅ�ǩ-D��(�F�~Gd�q�oL!22(8�	+D�Ĩ#O-os��iK��923�"D�\���Ͷk9Z�	 ��M��j2D�� 4��T(�c���$0}*İ�
3D�83�&@7
�TA��.��`S�գ��2D�@�+�[��(k�)l�h�3D��0��E�S�fp�	}Shp��);D��x�NWxW��b���*�J��l'D��@RAV�t���І��CIV 0�O8D��(S�@6x4����(ѥO]D<�W&4D��bO��]��P�/�N^����2D�,�L'T����)�%�\LH�%?D��L�7
P�K"�ěn#�Q�,/D��S4��#B���s̅��۶1D� ���-<�IQ!@3G頔�
.D��Ib��.�d\��^�w�@5 ��.D���B��KQ�=��G�A8�R�!D�����]�t�5&ɛ�D����%D�����׮�1V��N|NA#v�#D��bÇ,�:�ٖ/����=*� ?D�\��L�;q{��t�AF�M���=D��R�d$F�}##.Y���Y�@ :D�p��A� Aƴq�Ԯ'��hpL<$�h��	�'b&�QC��y)�h�I��y�Gͼ-�<rU/�O�������y�%�63��f��m6d�s����y�$��t�
�� #J�� ����yR�VN�481u�р{�����4�y��$f�RQ���s������ŉ��'������I8���f�#K�b�8����1���x3�*�OXyg�P7*I����'�ȱQ��94�`�E���?�v��YXftZ3c�39��� �`�'��8��ˍLon�j��|�)�Q��5��o�dsA��(�!���2dN�"�n^��`�!�<�R����<U�u�ʀd�T����wlRA
Bg� ܂��f̾b�=�<��&L�`���d�*>�A�$�ٌ;�V}�`�U�h|����'�ݘӬU�TM��W>c��	��dklqA�`ˡ��*A�Ivu�h��VW؞4��.N�����FU�Jd ����L$�����n�~Xa�/�S��$H==�xK׃�+~':�z7`����)�7�r� �T0#G#��g^���M{�'m�)A�$
�F ���%E�-��'L��q�B�r������>X̙Fl[�%�*d�pμQ���E�c���y���6�(�(�ѣ
�	u��XP��'{�tm��dx�������;$8�W�_)Y\F�Q�go�5� '�
B�m��Z?�N�pQ
#�4��A��	�?T^hh�闤2��1x�/�z�X��U?�%��_4W��8˰bÛ_H��85�F�][5�3/8����I�P��=��ԟ�7�C�[A��H���E�m�I&�n̓�'7^訫矇O�LZQ*�>}DPB��.�uv��/[E�|2�*��H_�l�1�I��f�����3S�*\|pºib֐34�U�{8XʒŊ�BL��W&:E�H!�ǂ�*��EI�J�9����v��(=jPH����Ũe2ʅ2>������)?i֝0kV���!�V�V��bمZ�ܜ�&�\�U���[ �u��i�iN�������T��:,8��3�h�!� 6	���C$����v(�W�WHY��J�>@E`x# +�2�f�A%���
�����9;@X9
$س���3:U�J3V�V����@�<N�r�#�ʠ7vj���">�I �$�U'A/\ݚW'�9+��12͒(Qt��E��[��Ti��APe�,N�·'K�*��A�2� ��6��f�jJ�d]�<3t��q��0hצm��Eϖ�G|Bd��d�h�l�@<ᳰ'©9�� 6�I#oo@�xT��}(����K�`֒,ʆ�ċG ������j�0��FċE.��a���q�t���dH$f�q0I\�'�蘥/�:j0B�9�Ă7�0�D^������VX�K���f ���l��$!E>oX	) �P} a0KF/KZ�����C H�?]ʂ�W,3����&��+��[����U؁`l"P$�#y�}[��K�]j�9h�a�#L���:.^r���L�P�Zq�+A�-�|��#�T4�j���7K��˲跟�Pv��?#<��䜔,9X�`���4T�=��G�I�M��c��q�tHs��,�r���rV��0!��+�Hi.OkL@*o� a��x<*���o�}���	n�ڶ>c�Z	&	�0/����@�5��F�U `��4��"�o3�K+O�M�rlG�B���(OP��$@�5_J��f��#6��hZ�I��D��ˉ�Y�j�q�F�O��!I�t#�\����hi2�Y���8���iR����&'I2��r"�	�[�fi�e�I�|u~�2!�%[��[N���U	�B�$L-X������>��)K�3�r�
Gm�;�����Q�N-sWcX�v�x=���	t|}��ȋoL8��P�7e�a�7GVhK�!��B}�-sp�'���8�D5"�F���]
<�A�%�?CVL���u��C�4:���"���*0�ԥ�5_��	�j̨!�%���|�w��/?�˓{��2��KA4�:jP�B�|��א���)=��S�)X��%��CRJ_�Z�����)uӶMbB�3{.v��P�kk�C��)tѲy1�+D�Z���`�j�c�`�)qR����b�$�3膆
�$2�Ѿ*V!�ĝ�#9n䀥�Ȥ+j��Ł=U{!��ˠA�&l�1d`�AB�	!�'괜{w;dfn�c�G�8R!�d��p���X�X��ꊛF��	>�<��b�}��ԫ�� 4`L���բ|�d��o:�Ox��m�>k���c[�?x&��Qe�s M���X��y�#�3@��P{�|��Y���'�O����	d���&(�S�o�����"_,|�!��	^�Su�B�	Y(� @�h^�G�b�r��ݢH�jر���m9T��ny��9O|��+4d��M3bܮߪH�"O� �ԍQ�>�e��	��|S�;ON� �m��W:���))<O~q����cF�5x�Ȑ'�^=q��'D� �7
�a���Z��	���pp�&y�Qx����#���Βw=(�㦃�W�^�ၮX(J?�#5��#�b  g�G��x7P��$g�6`��@2��sV|x��w�:M���&R�1Õ/P�/��`hӦ.%8Ir%�2���s�d!��˿xB�=��� t�ՙ�m!D�42�C0t0H��M�>���q��~�㇀�'I��ڳI	\x�����=�1��3x��s"�<�O��!&o�=q�����A8�����.Rn�:����w=��h�S��yRe�k��e�q+��/$�u��aQ��HO`ͺ�CL5s�0�|J�"��y�NM���ʦ�h|xҎ��<��O�%z^�h���1j��Y�G	�	�I����e���\�k�p�A�,�!�?i�Eѷ/m�p)(��D����X�<��	:$4uj��2����*c�?of��c�%3씢}dg�m�Uf��;�d���{�<QĂ�(?�� �O��HΦ��I�F&P��Ӂ���	��H���	3l���`�G{�q���'j_xC䉖m��x0' D�=��m��a�7����h'���=��jJ�w�LL���D�&�Lx�J\؞������D����'�-)Y�!�z���g��xh����'��x��ʮrB���D�I�I[h0:�}��R�\ Wc�R�O'�T�2�V)
grDx�E�qF�,��'�epR(ܠ.��c��K�Za�,�&@��$����>Q2�>!��.
\��$�*d�X���_�<1ƀG�f�����ϥeRB�zCo�� y��h�X��Ɉq�E�2bF�z]HQc%m�##j����+h�Y�';�H���Զy�Lx
a�@U��i+�'��(����H:A�AR��ၪOLR�I������ܽkrPTi�N��(�phH��0E�|�a�	�� 	7��#G. ��ꂙ%��uy4
	�u�<̈́�8��R�4.�$A��-�$'|EDx��Įw&|�ge"i]�<��w�E,6z�E+t�O�5��}��"O� a�`R"0����;�<��V��o	2�q2A���S��y��?H�0���E��Y}�AHw��y�!��1�Ys�*!X�r9��y2�Q4�� �EkFaC�y�	��E�����ɟ_�ȹ`q��0>�.��5�(̲$��#z��DH�GۋS�
�j!턪G~�Ѱ�'�
���I�7�S�O0ZM���D*
? %Xfi��� �?}�%�R �z=SХ��
��!��$D� $IΘQ�Aڰ�W�tm�g �"C���I����	�p핧�����2vxH�G.����0�ҹ*&!�䛎{�%��NG�)��۰.�/~,�ڢ[�z��2��;����D�?R"6Ih�&̀/�4��(��| ":~�:��Ԉs�Ւe��2<�d8���iɰ��ȓR�`t�G���Z�3�&�����鉲4������BY�O`�0˰$Z; �.��D��*?�0�
�'���C2�M�|66l�ӫ��?���
�'?�� ���Y��)��U���R��yB@�(_�I�F,�?������>�y2B>�2�E�R� �Z1�^��y�c@�2yJc�k��J��PC��y��̱O"��3���sۨ�� ����y�n�[���!`��0c$\�`���y�̌ޞ�;�n��`-p���'�y�.}�*I�p�*��@]�y¡��TH���ܩ�
�9�ʏ�y�Ģ`��u%!�l�~Ib����y���i�l��8~.a�q�͊�y2h��2 �Q���6m�� �q�ۧ�yb�TnX����ԚcJR��Ce\��y2c��*�$j7��!K�h
s����y2�L�d�P����Sl��r��
�yrʒ�^r�ai�"_4��I��yr��2`,0�*���W-n�!�W��y�M�=D`�ժƅ@>I�*Ԣ��ybϻcʦ�sr�_�F-�����#�y�Q8x\b@�6��c���4�y"�=^�eavb��S���s���yr�M�X%�P,�N� ��A���y��W<tO�u�7���2F	:�y��/qM��MQ:��&� �y�Z�L�T�R�O�VР�!ϕ�y"`A�W4l���'�ډP!`J�y�
�L�Ā�Q�cX�p^��ybGV��Y!���=B0��y�dI�0�x����߂�F÷
�""F��p�l�:���P�'[�;T��z��J�J\tR	�'����mW�T8�W�ɼ'�<��'�H�2[�4	ׁ�3 2<x	�'��1)%.Z	?�,���`\��y�'�\=�t�M�5����%JӿF���'Q�|��� 74d���9k��	�'c���ċA�%��s�N�4l �	�'y�P`0�P��	5�ݦ,�Bݣ�''p����7>��XRCcR�x"ld��'�z-b��TA���1%��'�b1p��F9�Q�flϬ)t����'6�L*��7,@�Rfa#Jz±��'"&��A�֙29������Y��'6tq��P�B�!s��Ї6h�		�'��0����d�G�
5��Љ�''<�@` �p�`��f�H�>_"-�
�'厤;s�����VnX�80d�P�'�h�����S�h�k6|S^4#�'�@�Ƥ��;½��/�&T>��'x`@c���5,(��[�1��@q��� ��yg�,$�@z���R�L �"O�-���<U�����MśPO�{�"O>T�Q.��v�|�(���8�1�"O��遬ن\���#�kP��`��"Ox4b7J�Y�4P3�k&�2�[�"OTA�1�<'�|��H�x��	�g"O��R#.[��y�ef%� (	�"O��"~v�y0�F~MF�"O�xGoۡA9��D�]?'����P"O��x�"��1��)0V�ǥ92�B�"O�,�1a$ c�I+�x��"O���e��<nϔ���"�
e���;�"O|ѐ2a]UU�,�9��t�"O>�фA��ꡢP���^�*p("O���g�(>y�g�0�j�:'"O��a�U�e8�$�ʬ{���b"OP=�-�

v]�ы��K[�	ca"Op�I���S��r!V�nA����"OfT��1f۔5Å`\�[5�5�U"O����-ͣY�� Bb��"#�l!�"O``Y����w_�, ē�`p$g"O����SET��:��T#�m��"O�d(���1#}�$��̸r�"Q��"O.]@�`�	e�����2r�@�=D�(����4�.�XФ�tҔ!�*'D��ۀ��"�xr�k@J�X�)&D��S����4�rH�� �*h����M$D�|�J�\�&x�nۯa�V=Pv�"D��B�6P*� `#���P�&F?D�4�aD�j�0�1rK�7K:�ɰ�8D��p��uA�I����32�Q +D�Xz��>"/N���NF4w�.Kd�.D�����"����+Z�.�ܥ��,D����4(����f���M��G,D�0K�fEb2ֵK�B�(ش����4�I�,Ф��˓VXt�b��q��X6��6db&̈́��RPd%�1+\�b�@"��ބ/ĨMq�ۑ��C�	#G$e�E�D,�TMz�DF0�z��$.~.r)P�{B�I�g����K9OTf�8��y��U�p�$aīJ:,!��� ��DÊS�dx�{��	6|����$�D�h� hU!�Dֿ`���`g"߀;خ��T   >TqO�Lj� ]8���P�q?�	�ӎ��rRPԨ��5D��Sb�
-8l}��G�69!�(p��%D����
$�"�"�w����n9D�D*%�32�B��"m�
�6��.9D�{���xSn	�v�[.Z���)�l,D��J��Ɨbt�ga�K��1�W�*D�xbe��w��D�u�;���S׋*D����*A/��A�B ��F]�@�#D����	�V���a��^p$K'D�j�/1�lx8Ĥ[:�1��#D����$�~�ђCؠ5� h�,D�|P��.�9#w�ֿ�C��<!J� ���H�S�$#�^��R�R�=+ZP�W�
��>�Q��>)rh�$VS���e�8*���Gˏ�"�6i ����O�9@���&5�B�c�ؼa�ؓ�鉌O:��Pvn�*?a`����8B�(��xeX+��V|�e�BݕEH�X�S���&Ӡ)c�oO�p=��Y7R��*�mˁg4BQ�mզ5�@��33�4l:��^����IO�(�eۡ'�R4De5H>���.lTI� �$�c�j��y�NL�Gh�3KZ"��|Ű�~����y���9T�(`��.�t��6GBrJ}	݀��T��.)�zt�2Mi� ؑ��D'�p>fKZ�s]�T:�G��]V�+�+�C���IϻS���y�aݜB<�	9��9�g��w����]1O��;wm���R��&��2�%i3�I�V.�8qa��c9��� ��<rj�$k7��3W� �У�a_�CŪ�0r�$W?r��2lZ��$9P��.c��Ap��'���d���j�^-A��
J�<@Ehƛ.v�8����"4 �͢���34Df��`���*^^,C��<J��=BA`n�>|H��֬m��Jc��x�[!"O LZR�P�5Ѡ�,�- ڔE���WnX-����FԒ1@ MXV�ʦi�M�[�؉X6x�a��$��U&e�!�qW��ˤg6�O.2�E�lE�2M��3�
ы���_~�ڗdO���|9Ѯ��?���Ǐ=��e�4AٷSm�Ј���{̓o�jܲ��G�	� ɶ�O�4�-Fz�`�1�����D�d�eX�]3ZK|Q�ƿ-���q�]0|�Â�ի0 �ن� Y���"�Gl�X���I;��"O2]�h���!�'���	�r%�ゞ9)ڒ�st ��z�vWW���pC˔M	l9;��~��Z�G n�fdh�́�+ P�q�
?D�`(�� pmΕQ�Z�x�a��K�j  ��T�1�,�J��(��`*���ON�W�B�d�(`��Gz�E�厏� ��5��ߠ@>��G�9�O>��A�A$9.x��V7]�f4:&�I�2�*|	�� ]>�uҟ'2�E)ǦҷP[� ��N=,f58�}2�;pA�)��ɟ�pK"[?��D|2��(��Ň��ΕA`��]#l�S%P
Zp��!`��?4���J	����9P���G�'p>=���P�2�$ �2��x�'l��֢�C���)�I�'�><��Lm�0�,��y�O,�m��d�-5\�؈�h�&[����'��yY�� i�����8~<;����� ��8O�s察�o2~��'BܵO���{썒EK^-j��f���2���&|�|�#�M�O� mۢ���.V�����d�f.v�ZQb���Hh� [Q��bq8o$�I"kG�>���zr,�(`�d��/��]1���B��p8�e� 9�
�%�>�|�����i�v��+߉0�R!���*%e�P;m�/@p|9�Y'[��˓A? ���L�$lp!�BY�c\�dYt��ʧf���H�?]�4��MW�o�޽�ȓF�5�$��oRQ&��$I$"�i��I3°�t.�3���I֡	HEȟ'�D��W�H�W������

���'uD��I� U��	Y��ۍ�(�8��>�D[�_��ppu�٠H�Q���⌇��q�@D!^�hr
7\O<�'�N���ԻA���"C�H�;/�`���=G�R Y@�rTa2�<� c(J=|�슔���O`l��+ q�����TN�-��	s)�{�Di�0��y$ބr�ҙ��B�P%!�B
��Č ?������+����*�"'��T�v�C;�B�	�iX,��^�(�xBs�L�k�B�I	]72aY�'�d�v@��._�ZC䉚����@�>�Z,�%eڍj�C�I#Ir�d��H �FH&�y֯�t{>����9
i���!Y�����%6_�i��Ꜣ">!�$ݖNMȴ���ӊ"���C��F�"2���R��yj#|֍�#Q
@@��i��/���x��J�<1PhZ�FY���g��-u�0a�����<)%ێy~���<E�$#VE�F 
�d��Me,]!�#к�y�h�"_���`\�@���&G�������H)�w�'z�HZ�i�"3Nd��ۯc%n���b���G�>�X@9r#��AΈ�YrBۖ%c�L�ȓC��8v�ՌH;ry� 
�S�2MD|��C���ډ��	g� K���?5v�U��!�@ Pԛg�[�|W�DsBÇ?�!�dE:0	�Y�R`N�%��,J��gN!�$�+"�UY�"�$5�^A���),>!��O�'$*���l��5�
�tH�%)-!�$Ѻt?Ji��C�9��D�&�P�0�!��<T��#���D"�q��hޯV!�d! �Jt!��#��'H�PQ!��P1f��������̔=����&D��j�ř2޴Y��D�W���"!�%D�T@�,	�)q-�z֐�X� 6D��bEǙn�xi '�L_�$���
3,O�ђ�N[̓a�&ɠ�hPp�6�O�f6�i�ȓ#a�lr�%�,U0���H[@ԕ'�@��)��ا�ONBe�"N��.-B`�?0���x�'����]�p��x�$�A�x��}�CF7���]���%��b�#`�t�2�Q]�!�Ģ;��Y&
^jܻ�fY��CK�\<� |Pq�[�:�F�����*p��%1!�'�V�ˎ{"�+<�(�&�B�iD�qPđ��y�HZ>?�Ё��&x2(��C�yR�FuHI��$ t�Hh����y�eɒJ��Ⱡ�#o��i#�R#�y���
X�ZesfKZ e��Ms���y"�B�n�2!�A�ψ�bՁ�+�y"M	w�P]����5	�Y�����>�G>>'�Iba�_�E�@�r�	6@��Ȇ+Y4!�6�t�T(�p.�ݱ���&(���`�G_2Xj����|��2E��{I�K�戃y�!�PSR�8a �P�H����Boy��JK#+���K��s� 0��&W�C\!�q��+E��'�B��"`��q���-؃i�T���O$���F�l�lSϓ<��]ȃ玫sDL�{eJX�~݇�I�n��C��G����M:k��(;�A"�@0�'�z��U�!��T &�Q��|�Y�'�$���˸g�����3�`b�'�.�k��G�T%�Y Iͮ%h��
�'�	��	^x�,ȓa��#/rY*
�'p���l��c ��L	�&� �'��u
C���hwL����=�@��	�'Z�t�v���~�%�/j@�};	�'(x�j��F��:i�bO�J��j�'�.lbu���;c�}j�Ë�r��
�'��EÇ �,gh����� �	�'%~��-�G�^\���3��H	�'������7H1��GMq,�{�'��lB�$Q�'��i"'���'���8�G>UvHyDO��
8vyQ�'��d$WaD�8��ً�����'��}j7��#x�>��*��tr�0��'֝�5�۪I�M�aꙚo�j�{�'�Y`A��� ����n�@ɇ�z���B�Q>k��p�+�1\��T��#J�U�1�A�;�FY�ǭJd����u\3[P2���0� 
��Єȓ\��ɓ="@08q�>w�F���h�l!�7adM�X钾r0���ȓH��`x��D�����jN91�f���H���Y C���!��;']��ȓ?�=��lɣ\��!) �9H!�x��6z[�Z�hN��F�ڼK1:4��p���T�P&i��!�Sj��M����ȓ.fŻ
5gٴq�t��p�P�ȓeY�!�T'|e�YUDě;>nX�ȓl������S ��d3"E1PE���[+�`��㌬0�H�`�M��1�1�ȓ[���Yӣ[�{Z6��0�;?���ȓ:b|��䈑&d܀aDŜ,�*U�ȓyؔ�����'>�"�;$�]1����ȓi26�A���> ��K�!M�{��ԇȓz�����\�g2�	cc��E���H�VЩ�̨�,0b�j���ȓn�#Ɣ�`��=���E�����t}k"A/�� �ˈ�-{����j,�Yw	 4�u��!D�GL�`��Ӿd���h��$���REB�m�!��?qw j�B��,~Dd�7k�B�!�Ǐ\��}A%�@�Z �)�ȅfj!�$H)yp4�q,� P�:�BGJ:�!�$"w	t��爒�b��m1e�X�!�P�,�FUXsn��h[aKG[�,I!��9q�l�b�3Fp�[�e�4�!�� Hl*�=R1b�т�f�<�C�"O�;E/Oo |��C,	z�,��"O6Xs�j�jc��Bf�Ši���"O���jTq�"x#���/t9�|0�"O�tӖ�|�����;��
�"O��Q�@�$v����f�v�c6"O�Á�Ө<�i�¤�!N,��"O��B�F-	)�=;%��EG6A¦"O��5+�A0Р��э,;��*�"Ot�VZ�6�C��.u[S"O$u�@�������Dn���F"O��j#e�+&L�6�O"T�踪"O�Qf���Cm�=�!۷_�ѹ"OpU�D*^s�� �T��-Ht�R�"O	�g]�T�bH��ơ77�[�"OX��G����s��`) �²"OpY�dES�l(�b�?."�0U"O�h�wd��N��7�*u`:�"O�1[��('J5s��Bpn���"O:s%h�c�D$�d��{P���r"O,<{�EO$@ Mz����=��b "O�Q���Y�u�\C�2x:nx��"O89�Rʜ3&�5Ue��.M�"O4�[��6pr*�T�	�(t!�"O@@"gN8��y�5�T�HB"O�]0 �H�W�С:����a�����"O�X�%`f���=\�(���"O�X0�$څ[�R�:�G\>H�vLq�"O栣�G�41�2�&�4:�\�"O�����څ
9DT�0����!�Ě�X��T[�0aWvU�f�
�!��7~LZ	��+�,W%��J8<[!�SL��AN�VU@�K</P!�?J��h��MލKĤ��rJ��!�B$m�  ,�L��@�`照q�!�P0#�:a�-�>~��r�E0 !��
h�ʈ�T�~����G�l!�S	�4REZ�Y!��Mg!�DI�@̼䡶舤|�^��E%�$Ik!��~��Q� AC&	Ӥ�]!�#��\���M1
 �fC�	L!�D��$�j��]XĲ��%�\�6-!�$�B�\5)AB9�~�"��ʇH!�Ӎm�n��͜JH�q҄ޟ@+!�G�+����)Ý3`�d�,!�dݠbށ�(�E8�CBCE�#Z!��زIT�AegS�J�&I���0P��NU(�%�oD6�Kb�G.ij0����� �s��$SG���$�E�ȓ�r� a (p	�5���NY�ȓ�J��	Q�m}���M�7�4U�ȓuuF �FIO�\G\)
�o\�'��a��n_���	b�L�MY�i��܅�'n<S�υ*��k��S�u$����l�Z����K% #�1�� �;% HІȓmV�Pt�P�@a����I�ȓK�	J��_+E���aKЖg'�0��Vb��G!>1T���>0Nh �ȓ~��9�ҋ�,@��!I��E�ȓ" R!J�ʌ%L��"��� ɇ�m2�( A,<4��\,��T^���FN�f̂`"�e�E��ȓ��5R6���ы�E�z �ń�����y��&�P|6%��S�? $4������)v���];��bG"Oz8@F�)J�h�Dͨ:}�!��"O�sĊ�mҰd2�2v`1�"O�S�j�Y���h����Ҏ���'���3R'Ӿ�uS��/̨ɪ0M9D��jA-R���Q�Q���P���!�b3D��xtAј1��{@+ƼR����A�2D��d��5�=��"Ȱx�^5Jgn-D��0�"ݙ'���ʷƨI�Hi*�*D�@����p���qe�"\�.�)D�lS��%䤙ʁ�b�ʷJ%D�dۂf�(�
�@�OZ*'rؚc�&D��+�B�9��K��9XW�P s�.D�,s��=8ݲA��R�z���j%B7D���M_1k��B3bV&^tb�4D���w�б)I>��qc2(o1D��lD'�J`��? I�%��_�<Ys�'0
f�J􀅾&) $�b��ȓyD�d��?�T�1�	�D�ҕ�ȓ<T�3�֋UZPYb�!R<�
}�ȓu�L����Z`��"Ԅ��$\��ȓV���Hp(B/�q�3��=\4v���24I�q�IlM��/�X�ȓA��b!�
'U4�1�AET=��Cbe	'a�L�� -nV]�ȓ�za�%f�� ڵK�)��|��8��e�\d��On�:D���T�ލ�ȓC�����������S�Q>|�X��+p*\BկB���X"��>}�R\��c�,Hw�L�t"Y`ň�`�@�ʓ}evm�f@^D�@��#���:C�I  ����S&Jv>��%$I�C�	�p�lT����@��-�WA�,��C�	`�q�-��E���vf�>x&B�ɖm)nMp5HΜP~��ұ*ӿt�C��3��)�*t�NIS/���B䉭8�0\i��]�(�
U���-� B�	!>����.�z� ��ID�>�
B䉪'���#�ԡm�����ˁ� %�B�I-/z����	�:6�I���8e��B䉱"��ͩ1�X��m��&ǔ��B�I����:��U+e�M�#�� Q��B�ɽ�R�o�V��t2��N�~K�C�����▫�	R�ܴ��/��*�C�.� ��%,	�^�t!%B�RC�	%Z�: S�3�n(���"4UxC�I�w�K�/�5H�8��-�� ��B�	�i��p���\;8L���6	Y+\�C�	G�(KP甑4.�Aa≃+��C䉺C/�y��ŏ�Da|C�f��}<vB�ɐj��)�1K�5k<1@�/��-B�B�"n�	�f��/����	�0|B�;-�(�%��32�C�ņ�0��B�	�;>�"��ŉW��Y��$��B��, �)�홛E����V�)Y�B䉭?Y��	P瑜-��hQ�ݙw��C�ɔ/��I"c���#��f`݌L��B�I7�2�`��] �9ae,)G�*C�I8<��v� 
!�m;'Z�:B����}����N���`Ù��C�I#qyS`�j�Ы�bZ�ZU�C�ɯXT�Wm�~��Ybv�� C�ɘ;]�r�G�6Nֈ1s!H�3��B䉥ZM@A��+���c"��0�B�)� �vQ0>�3��^�G�>��f"Oԋ���"�9���șK�6�Z�"O����mԖw�D���
o~�U@�"O�аq��!"1sv�<f^�5��"OL�+GËA��Ke,�O�W"O:Pzu����p3,�-���"OҘ��퓾|1@Aa�
ӹm��ś�"OL3�'�Y~�`��_�yz��{Q"O��H�`�1z歑$�g��!"O쵢�@+du��*M�U�q��"O�%�#�Ֆ`dF%�O����"O쐁���I���q� �4o���p�"O~l��Ŕ�8�p��nO�>L�x"O,���K̻e4��rnD*V��Q"Ol,�a&ʗeP�L)�l^��>�!"O���5��lj|,S�K�q���"O��Q�!I��е��"�"ORUÖ��(n�2Ɂa�C
*�:�C"O�=�T�H�x�F��Dd=�$t��"O:�� �R�o�����	B�Ne�t"O~�S��
,/�&	�3ⅵ����w"O���V�A�4|EA޻d����f"O&%A&lA~w^,��O]��t ��"O֠�� W�`L�M ���*J<*��2"O����&� .�q �%#&�]�"O�!��M�#T8~)aD���,��Ա""OP���uv źF��&,Jr"O�%[�y��&V�b�"O�iAk?J̜��^q5��aƞQ�<�6�۠S����aMF��ye�B��/gˆm��*�i�d�"��*K�DB�I�rrDܳP�X�'6Y�G��!F��C�I/�|�`��O�pN*!)&�B C0�C�	�dt|��!$�H#e�ц��"{�C��,EQ|RRLʦa-Jh��"R;{sTB�ɮ`*<Qy���/�HP h�!"��B�I�@�
̻�/8=�T	�b͜~�BB�I�m�Q�T!^+D�IPi
P :B�E��9��j%v���_�\7hB�I�=4�C''��j4��9���0:B�I�C89఍�Li���5LZ�vjjC�I�vT^�Т�W��ܥb��V�� B�	C��e�aR3��љ�MV���C䉶>�|�y�o$j��@�O$C�I�i��e5K�(Eh�O�;��B�	y��싷"Β)p���M��7��B��1b2t�2��*lL�����M|B��< �r�;�m��vp9d.�bVB�I�I�A@c�f��;�̒-ĔC�	8y=0� Bb�&������
}&B䉚k��$HZ�y$��
���?�`B��I�>���J	?����'�@�%��C�I=!�,�
�!P����#��`��C�ɦ+�#ҥ	G8�ȴ-�ʹC�	�>%����N�H�X%���N���C�	�m�� ��2��&PCI�C䉳s����!i-,��`X��+�(C�ɷ;���3h�Z����ڰvN`C�I,�61ԏ��4���X��p;>C�ɖxt��J�)J�k'���X �>B�	�R0�,`�O�F
�$�N՝e�C䉢Bt�Sq��(�p[��GG��C�I1C6���i�_�\ k�>dvC� ¬EXu�8T�`�u脰�C�)� l]�T�� HjU��ᓋK��9�"O
M83f�5D`� S��٥(���T"O�%A��W�`=�X`�݁v�Z�"O
�K�E�k�,@�
L��BY "O�LC�Cӝg��!�L°τ���"O�$��똏pjae�],���R"Ox8�I��2�V��tע}J+�@r�<+�+LvTIrP$�>���7��r�<9⃔�c���ؔ �zl����B�<!�o
��|	ئ��_�`��X�<��B���e#�$��t�D��x�<�c�Hp�|劶[�4�y�Q�Cr�<��fY��&8z�h�Z�f Ѳ��m�<At�8JP� �W����&?T��b��B+v��Be���h�T�3D������S�91�J5[�ʼ�!�1D�0C�M�����Ɲ$L�T`�*.D�� ���;� ���*V>WєpE�+D���MߣRk ���G�.�|���O4D�� 1�7
�P�J��޸d�
y�=D� �b̂)l|%:�꘿Dh�� �I<D�D����	f8!�� 4�V�9D� �f�#N�l��1A�
n� 4�@e%D�1��ުg�2={vHT�m� \�C D��!�P1V�zia��7��平�?D� ���W�/Q�$���6Q��Ѓ��=D���ů�*���3@��W|���n:D��+t���U�B��/D!�֌9D�xH�*ڕPH1u�[�����-D�ZwD2=,��f�ʯ/R��'& D����m%W�:�c�I ,,���4L0D�(*�텥?�򽠲��U����0D�!F�-��J��EKt�z1�+D��s��B�C2��Sk���`�k��*D��6
C�ri�}6�S>T)r�`�%D���DΛQ��E#��о  ��g�'D�p����\g�y	�.�l�W�#D� f]
�j�m}Єٶ'!D�D��#�M���s�'	�,�Ve�%�$D�x3��ȰH�H�1@I ��! �"D��JgB�Q0�0'��p
(��a,?D�\#@H _�"��E�̭	��Rb D�[��/��- �]8��u�7J"��<�w!�x;r��փ_�=�b��c+�B�<���<^�(+LT�o�4�)�j�s�<نmU	H"i����#x��91��o�<)T,��p,�i6,�*4�l����g�<id_#`�)��� @���HHD{�<�,O�s\$��1��I���� ��P�<iD�D�>v�0��狛A�V@#�n�N�<����0���I�O����9s	H�<	�AǫL��X�2f�)2nM
t`�G�<��AA�3�q��E�L�lhc�\�<�!V2P�d�F���)�L��a��V�<��H�K�P󵩛f�z�"�W�<�#G�6AiX9	С��de�"eTV�<)����j�Vn�G}�X�S��N�<��gN�	�4 E�s؎���eI�<qTGd�V��c�XݐQ�ƌ}�<�4�uj����b߆� A�Cw�<�#^�Sޥ�q�ЦaJ��ԤOX�<A�b��f�"�VND7_~]R*M[�<��JN�2���r��!O�1xT-�P�<�0�]B��Q��)9�ڬ"�'P�<� ̱���
�+S ���,]#y��,�3"O>0�dLсG;@3�O�^� �A"O`�d��,���D��ܸy "O-�6)�F�(؁���$���U"O=��.{W2� Vʆ���,�w"O�$�pl�&ϔ�TdP�r��,�v"OHar򌒢����F6�<�"Ot�k�H����y�+D5��l�g"O,�(�HЮ�F(S�M�a�Ѕ��"O.�x����"��<m
&D��"O¤څ�ѽ��AH�L	�S����"O"���P�C� d`#I�D�ȥ�0"Ov�C؂!}B� D�Ѭ@u�$"OhhY&��?�(x�`��3�<z�"Oj  S&��6��a�׋2���
1"O�h(Cʺ*��Ő���,at�Y�"O���RL�"EO�L���50T����"O(M���:����P�ͪgO0�@�"Obb��C�qw��� M�Wk�$y�"O��Xg!Gp�|�9#��>K,�1A"O*�����C�:���J�1m;��"O���4��I������#���W"OF0�g/΀�$�dO:+�x�q�"O���b���3bh�I�+o�|0%"O����?���a�`�!��)�V"Oly懽x�`P9��Z9��ҵ"O��saG���.�+l��`"O��`��ϲ4�l,9����[��	H�"O��p� �jB@����BK�"m�!�Dگ||d�����Т L�!���n�Ǣ�T�����kM)a�!�
7�Q�rCF�jg��0�A�a!�ļf`:�;Q!�YZb��C̝B5!�T )⍣w�R7^���(X'!��@8ֲ<�d�U�$?��a�N۽!��V!�8��Ņ�4>9�9)0+	�"!��U�4��P��#����#Z��!��!#������<ePv��P�$j}!�d�q�¹�)rN�\V��"@y!��,d����%SM��a�螴 y!�$��t���0q�NL����fV�o\!�$M9FbI�F��]�Y���S�<AfRE��5��"��6�ԥ���LJ�<1Ҡ��5�vm�	%Hh|�� E�<�0 �/\����Q�ًl�r8�d�A�<IäHǶ�[�Fؾx�䛦+W�<�$OD�'E�]*7��5�h�ӲF�l�<i�(��>ܒ ��� �9'
��w#e�<Qn^�*� �X�څ ���:T���g�M��b!��߁Q���%l)D�D���2H̘D\%/Q��(D���[���͓O�>E��B3D�x�G��⠬��I<��B�+6D�0r�F�8n�>(��Ŧm����D�3D���&�U�bG 5�v�G���p��1D��1ͳf�&(�u���,��|�H0D�t�!��(A꒤�9"F���$.D�营!?{\�Á@F26�l��*D�����^��	��b�P�����X�<��̩flXcpZ��l*r
�X�<�BO�M|4x���3�1"��GW�<��e�!�ޤˁ���,,DT��FQ�<	�"�&��dP�@�:lb�x��,�L�<�g�=O�Isg��;B�<��C��m�<� �Xb��G�8� ���.\�r(��xr�'���U3[B`4�#�g��x�'&,x�S�V.Ԩ���9	��8ڮO����`\� �AlH�~Kj��2�H>��6�>�M�"~n?N��邬�.0n<�{'�+�.C�Ɍ1/
�uL�-&�r�@���C��=0#6�Išò6���@��@"O�����-*������'�H�R"O��hTb�p~蘂%щN�ܸ�"O����L��fF���ĕ8 ۴���"Oek�.<`Gt����~�:Xq%"O^�ˇ�לT�x5�۠YXp� 7"O�ɓ�덝R��L���\�1OP��"O��FX/+&L"�X0ZX��"O�3�e7����� ��D�(��6"O��Qt%\�zO�š��B�Pй�"O�8c�a*&:��R��HH����0"O>��s�M3
@)�e�f4d!��"OZ �`kA<nT���,|��"O�R�l�aNy��!ӂ0x��ڳ"Oj%�Zh�r�V82e��F�Qb!�ۢi����# Q:��@��f�k�!�$�(k�6��稛9i�<��tO"C!��#;�v4�Sb�/e����O~I��'n�"� � ��x &@�$l2��'�X�`��(	���%L
3- i�	�'z$@�$.|�`� �� �(���	�'W.H����,0疥h�k�&r0$)�'@f���X :0�P� ?L��a	�'˜q�#�3
�
��2��u�|R�'ުI��AтFʦ��b��>pTΉ�
�'�\�P��%dUb+Q!���I	�'	��y�C]�Z�LX�Q��X�X���'�ٚ�Q�H:�1�K5L~R�B�'��,����:4���DMD��X��'�V�zgg��"����r��&0\L5�
�'
�%��ㄲ]�Ps�!�$^{N-�
�'�9I�8�R�x!RWQ��1
�'|~��<u<��9�hXO�
�)
�'�8��7H�-#����oǾM���2	�'�:e,`|$�Z!.ԭG��z�'��Y��\�m8t�×���:U*�0�'Ƽ!�3%��)sPݩ�Mט{���R�'A�w R�EqP�	�Ʈr�n
�'�P��G�.:^({ӊ��n�Z� �'�Șs$�.l�0�2�ȸR��u��'霨0�7��0.�;� ��'���s�Ͷ�t��J���9A�';:x�5���
$�ŬҩD8V]�'2�Ч�]�|,�/��B�~0��'~`E˴f $�������'���kԍ���LB�ƕr�6E��'��SF��o�L��U͐^N��[�'��D�Ш�-�I�a��VFޝ��'tvX�W'W:G*]P!�{�Xp�'�5.U'BA�УX�>��=��.�c�<���1ly��r2�O�u�P�15_�<!��B"��S�܋��\1I�o�<a�"x*u݆!.�s�/R�<Q&`�-�0������h�*}k��c�<��$�	C.�A����4(�\ġ�ND�<9���'L9� Y Ƴ=(�	RC�u�<Y��V/#� �Bɑ-"�ʙ��}�<�7�n������e����a�<� ���ɵRh^t8È	�>n��w"OB�8������	�<���c"O�5�c�;C��H�CЀ�C6"O
ݒ�Ոx�r��g&8���v"O�`邃~X�Ks�Kg��a:�"O*��֠"j���:$(�"O�!ᑋϤn}
�fLZ�G
ʘh�"O:�1�A@�N)��j�	F�M��: "O*y@�X�԰略�l��@"O؈��R�����_���e"O
h1�
�<U�F�s!��;Q"y��"O���ǒ_��kť܊SJ����*O����h�*eDD����<��
�'}6��𧟼�~9��. t��	�'^����43�t���^��bղ�'�a �c�zW8��C�̦��'�
�;ì�	��$	t�M6���R�'R�� ��A�5��!�NL?Pb*�'�J	�GJsv�0� ��KZ�a*
�'��Z�M'o��Q ��4=�^��	�'K<�J�m�� �8X��!�:8*f�C�'~ݐL����9��م7�؁��'�Y�C�ɏW�`��F
*&4A�'�B��e��%�rm��h�(����'�x��>_��A�ٽj6��'���
PM�0d`�e�x��x�'|���0g�>h�5k���$U��'>ą�7d4�ԭ�ħ9/����'�Xi�CB�I7�k!��&���*�'�J�;�ƍ:^�TU�q �� ����g�~(�r��"J��9�aɗ
fH�ȓh�f��whХ1��@�&d�rA���ȓ��!&���v/��l�+F��̅�V��H����� ^*'@��7`�Z����� �*�-�7��M�ȓ�ֹ��/Y�r��P�3�ɞ?^�E��i�6|H���q]�hY�*@�Tݞ��aM4�rr��L�T!鄨�!y�نȓ�2LpW�H+*�z���B��
��ȓE�H����!!�ҁ��C8N��ȓ�<IR� 2H0�,h�h���"O(�b�F�3P����ʅ���"A"O�Er"�Y!D}�)P�K$|����`"O�x���_��J� 
#w�`4�b"O�A�&�8y�̙�W�M:)��u�"O�`)��/R�0��ꎔn�Ґ�1"O�����$�J��zѰ�J�"O�"�f���q(ȾZ���"O����e�� �%Ɏ�v���"O$Mۃ���R�N;��C���"OD��N]	]@�гh�.	��9x�"Odع��5^�p#IȻK~z�+E"O�Ւgꋙ"�UcG	�CM�p��"OFH�ъ�V� I�/�EQ�<H�"O`�H��\�:v}�.�]bD�Ѕ"O�xC* �5AV��ä ��s7"O:I���:N�t��4�2<GЄ�g"O���1Oߓs���veؿs(�! "O�a�eE!\yH�#'(ޡA�"O褒�ʂF�
9@� �N�<�q"O~���,O��D�ҏ�d�Y6"O��&"�!*x �e��W���"O�\b��З$4��.H�P1!"O�����Ș{�Tm���M�V�x�"O� L�0��;S��ݑ��֍-�z��E"O2Ԫ��� �t��sO�*Ǹ��"O�,�c�wD�ha3��I�"Of���B��p�`��#���x%""ON�x��+h ,��W�N9n�0�R"O^t"�� �S�.����'0��a�7"O^Ԃ�l��ZD��f&ϱ^�0 #"O��HL]+t��`2Dԧf���J�"Oؙu�Y�b�VE�T��""O  �	sޚ�ۑo�9�Q�5"O���/��CB~��G�X��x�"O��`u)�*x�|p�,�Zǂ1�"OZ��*z�*()`K�(#��(Y�"O�)�K�W� pDQ+C��j�"O� Y�o��]\��
��,A�`���"OJ�	�����`b܉#��р�"O��ӱ�[����oK&>��y�4"O������Q�4��{���"Od���͒=XHɢ"$AFt��"O�����,R��q��"�a)�"O�b�I�X��t���Ќ���"O��B �>(>�#-��8�z�"O�А�ƥK*�Q��� �2�B"O|����+P����,��'���ʢ"O¸�e�S��{B�2N�v�I�"OTAPr�L�truH ��AY�"O&$�s��00�!�e5}�m`C"O�p����>c%��AjжoA���"O��+���2\�u�5J�"�m��"O�=�f���JXp
�>jْ�)"O�=� $p�T��B�J�M�"O*���ԲU�X���a�H�ٓ"O���p��gjl��f�P%l֤�`"OJ�y��	3�A�v�.P�D�9#"O^5P��U�%Bq�waƠ@�\�H2"O�`S��J�-�.L�C��P�X���"O��0d�7���*�/�35Z��g"O���ׅa@�KN.H�xw"O��0���a� yd�A�"O$0����&�UFݾW�&��"O�Tc�lE t���e�P�65c�"Ob�2�C/�a�NǚC��Q�"Ol1з��$���$K�-e�t�8 "On4)TW�9�����.4�,�"OZ�����d�N(�Pd**6���"O. ����=e���C@�L�x'�H�R"O�ҥ�"`�RQ���4C^�@"O�dh�IľU
Y2%��'�x "O̩�wa�Q?�y�n�#G\�ڰ"O���N,T?a���.QZ)t����	@��<[�%T�9��ʟ��P-���:D�p�S+�`X�#�@[�LAKW�:D���R�C7n�1(�Q=92�"D��ʶោ}��mB����V��2է%D��A0$��f}p�x�GK!���TO>D��h4�T�Z�,�Rb�Rkr%j��:D�Ġ�M�)n��kӎ�vmX��=D���# �/Nl�7��=�0e��&�Iz���x���9���E�&����G�?D����d�� Qd�@��vT��Ao3D�������6��2�(�<,�;`4D� q@J<Q���iF���>G�)9�'���D�|c�-r��KB����
�'s`���Ȅ,AB\ё��!9Gδ���� ı���Z�¢�+v4U���<a��4�p��2�Շx�v�Q�`��Smf#ǘ�8���JN�b���?J�*�cD�� '�B�S��]Y���KB`�P�)2pC�	�d���9$����|�b�i�sOhC�	.?��q��-a��@���;@BC�ɀ@=�a��|5H�iRjX�fY�C�	{��]"D �
s�����?�,O:�=�L�pxe�X:4�b��e�rR�͓��?�%���[�Ni����;7�2Y�6"�T�<Qa!��\G��B�K�5#���-LS�<��!�������= }#YI�<�2͜)u���bG��fB�qC|�<a�%�L�<�C$�1l�^�B�p�<�ǥ_Q�ə���.��=�`�';�yd�oX�	1
֮j�Y�dKgt��Slt A�pe�-.!�aZ3�!�$�����c S�^�ʍs�R2�Py�Ȏv�>t3rAI�M��4��:�0?�)O~���A��Vp^T��6=L.���(�S��y�%6aY�����5,
Ή-W�֍�ȓy��E�8~����P`K n�ȓ��lI�I!Z�� ����\pD��ȓ �Z����K�y5Z�o2
�� �ȓ"��d:�j���U"B�\.Du�ȓl��ȗ��*{��p�`ʕ���}��D�t`���,"��S�/�&&$B��cH��g�[�.��"�;(�C�Ɂ5d���-�>��!��B�-�B�I���5�� �	 NC��hO>�*�%�"�4�`b�N�\�i�N'D��&�ײo��y�- �D��#e$D��C�O�d.X8V���C�\��� (D��@���5�z�Z�Λ�c�Py5�>��T�j��A.ç(��� �aI4,G$M��S4̼XۂQ2p�pR)�.>f���hO?�a�Q���1[���if�6?9��������EL	(5�9Җ�^��@!�"O6�k �\'bfD�X5O��4��"O��@�a�3T�91�͉#{��#"OZ�AEB0�*�#�A0 ���1"O�01�	�Pn�P���wLy04"O"X�3$	�ZXv�9 c·T<-�eN/�S��y����/@��e9�p�V����'�ўb>ѫ��/]T��R&-tI" M;D�8���,f��7'�>���DLx�<��� 2��7�:(���g�I�<�fZ[	>�b�,��� I�J�C�<	(ۚdv���vlX�9�G�A�<�уY�p�=h��;ԁSQ����'F�𙟌�r+�>zO�yI�#T�ՓA�1D�Pq��t�ق'���tҜ�j��2D��{��Wj!�1�PEb=FK1/D�0�$H
o����+���0��,D� ���s0�8�R�fE$�<D�8��!;�$đ��[$D!���:D�\�⦆�k�BS��.{/���`�:D� ��oK�P6@m��2@��1�7LOl�H�E�+� �P����^�yB�s�Dx��mL�'�� ���y�V
T!��c ,H�P�U��y�L@2Kд$���8�d�y��)�'x ���TTH�c�"w��A�����m��QP���8��Ї<tܕ�P"O� ��;V�ɢS�l0�Ԁ�r����"O�`��!�>O���-˖$?2��1"O��V/��f.0�g�M���u"O~��(i�N���k�n�P�Cs"Or���VuD$�!Lڏ^��yI��<�I>E��'Ī�q����r�"��e1X��O���;�)§#���Ȥk< �&m����Td�}��Zz욤I�/J��
���n�J�ȓ<� �cK\��Ij���/V���Q��H��*TD��!���"2=��/,@�sRaQS�e�1�XNK ��ȓ3,><3�O�D�iY����jH��z�^8
7h��+(��1�߄<ܪ܄ȓ9&���%E�!�F�G� ������?ɡE�{�����J[<{Ƶ����L�<!sbߔw6Y���ґ}D��Yfg^�<i3�֊mx@���(R���'n�X�<!���JhI0ύ'�hݩAfZY�<ɐ�G?Qvn���#��:O���wc�Q�<)UA�l#�̣�bƙL�\���K�<�q�Ñ�#�mH�#�h�:A��A<�#TPR�@�N�pȐ��P"T���a��E;֧C�*��İt���^��Q�ȓ\5(�3oҼX[�@(j_�+k���ȓ�
\����.��ˀ���-�~��ȓ.�Zc!�]-�j�%���jU��-.�)�$"�:TvjQ�q�>
��Dx��'��p�e�̘�af��l��	9�Or1QA�ֿs��!tiϥj) ��"O���'P D�vp�`(r�9A"OU��[�R0��N�bE��n��yr�H���<�H�'4Vl��!Y��y�B܄w�ܔ3���1��]� ,��y�gZ�j�Jy���-rs1钧�'��{��_�����H;��@�֩�ykJ�Qٶ���J(2�H���ψ�y�"�b�d��"��,'�B-���ד�yb ̳z|�S�"0!J�*U���yb���$�q[pFX^Sb�
D�"�y�*�:"b�23�)P*�T�����yR���
��ȫ�k؂�F�@S�+�ybh�n��Ʉ�Z�8 
\��yrH�R̐D���|DK����x��'�Z�&̞� 3X؛�Bܳ/���k�'�t�[�o�W�
yx�@Ι,3LtC�'q���o�a��fhL;6��|��'6�LP ��G=Ȱ�7�Q�_�����'��Z�_�+^��N@�l��,��'��cDG�)~0X��̫x�*�B�'��x��) Ii:����o3�5�㓙�D�OdM��L,h����o�#I� �(�"O6��B?玘KWnS%H��Y&"O��f'A w�U��=J	$1��"O��ddH�#��M f���P��Q�D:�S�'qۂ��g�Yj"��Z�ߣvv��(����ێ@鴄�צ�!�4��(>8�ᖩ^�/=4b����
XD��d����օ�W.��y�l� ��%�ȓM�qz�+C&s(&�1C
��Ț��hZ�8'	7ib����4���Y�I5���X��V�&kf�pmi��B�5���Eb�qVfX{�@��..B�I%�X������U�4䂤�S�T�B�ɀU�%��&�4_E<M���
B�)� �lb6����&=��)��|�VU`�"O�UI�O�3�1S�g��X�j�q"Oj@+5��n�f(#A,;W���'e�'�h��fաUU��ۆÅ �ȅ��y��'��y!T?U}����a�v��-3�yR%�`U�#�I�jR���yb�Ɛ:F�墴��
3<`T$F�.��'U�{2�ea��CFB%c^�(BL��y2�ثN�@*w-�.N.E�&A	�yb)@�wՒ���DoG�2�d�7�0<���$ڼ3P��t`X�Fh|��ef�
��X��	#:���a��I��P�	��C�	n�r��̉�-�h����T48ϸC��/����`O+6 ���$_���t��`Tˏ�5!�	�kN�p���c�6D�l�AΟ���=C���ht+ֆ4D��[�'��9���1�L�a���#4D��RǬþ_�ȡ�RN�sS��邤>D�TxB�S���Q,UeX���6�!D���b-ϭ{�r��-
o�ԅ���,D��gd�9Q��`��(�1ҙ�G+?�	�c}��QFG[�U��)fڵx���ȓ.[�xR��Z�#��I;0��2\�ل�$�~�Ȏ�j���o�kM� �ȓ��e�#�D;bS����`=��@�}0c��*!v��*� J�h��ȓt��p	��̑I��l�F*S�%�x�ȓDF"��E�ŚV$b�����1o�����V�9��ū	����f�-f��e�ȓfL!��*�*lb�C�'�&x�(H��PE�� �X%iFY�7J�()���ȓ]�ء�q��>)^��n۫t�1�ȓ#�@]BWc�S��|p�X$J+�Y��P!��c�B�4�� h�B�����g��ܐF/�S38@cb�U<���.��)�?�=�!G�(g�]�ȓK� QD�"J��)���$B:���ȓR�±S��(w�Q�w��"�����z���`��/0uQ���ܗN����ȓ/w� 	@�ɮ_�x�hu r���ȓ\\) rkN�7�@�yЭ� D��a��+�4�,JV�ɰ�N1xP]���!u�߿n`�\�2��de$p�ȓ�n�# �����,��ȓ?�l�BmD�G:N��4���N��ȓH�J�sPM
>TEBSE�'�L�ȓ8�6d{�jS�B���&���-0���E����%�2WVDaG�C32̆ȓM��Q�q�Ӆ:�0Q��2K;�\��m�(�	��\*y�l;$@-s(����[
�4j�*f��c���c/���{FŚ�'`��g'ی/�̈́���P;�F�#�Y���_1��1��_�����	�kBj�z��Ϊ`Յ�j�����5)X���n�k[��ȓ?�:h
�mR�&�:�J��W)u޾$Γ�hO?5�N�D��xh��ъs
�W�<D�h����$ȵ΃� ۶�"P�-D�8 g'L=<���9��#��Q1�,D����Z�m+�)��˫� �1
*D� ˓g��~"����*J���ɥL$D���T�[VPs��05�|��S�.D��`s�N�l�����͐I�E���^�����D�5���b�Wk�( vl�S�!�� �\�d��#(.T�f;�n1Z�"O:��A$�z���#�����1�����i��+��ȁ�+r
 Y��:,!�d���${e� rD��)��Í
!�Ă;2��ӵΗ&_b~apN�!�Ç�<a�0��Mi�|�4��6v���:�S�O&�+��Pdt��tIH<0OFLi�'�TsՋY�b�*��S�C�zt�0[�'��M�#�3&N ��u[ab�y�)�S2:��jP�@(|=���"iqnB䉶PgEX���B/@�s �V8u4B�	0�2U�2�4�lř�(��M��C������S��aȎQ��A�-nx�B!D�pG✃�0u��K���0` ��?D�dIC��,aJ��5Ɩ�H�:�x�+ D��R�ϑl+V�;em�{D�@2�=�hO�� ������-R��ԦͿw��C�ɑI����E+(ČM	�Ÿ�nC�I0BĒ� � l9�U��"f� C��d�,a�Q��B�!P	ґp��C�I~��0YS�Z�
�p:���*+&�B��^-���㝉e�r�h��[YnC�	�y����5�"��e��c[�C�	?H~8�p�O��V-�I�B�WE�C��.n� %�ׇ 9�6$�$³PЬC��)QF,H����3������x�RC䉀�Х�&�� �5yӰ�hC�	�f8lD���C�v��4���Pj�6C�	�`�|� �(�6$Dp2M�,xyC�	'�.��܂E��y㵏L�XS�B�Ʌv}�Ȋ�G1�9J�h޼E6�B�	[���@��6rua2�	
DJ�B�ɲ=N�A@)P��TM�p�/}xTC�ɧ���X"/�m+\���h�C�	�F�l(�ʔW���N T��C�	�N������"iL}�'���"O��@��[��ؗ�E�e�V82B"O�A�2H�Д�2hQ�kz���"O�y���σN��]{�'��X�ۂ"Op�Tb�/M�(��Egޖ��0"OL����ШY���x3�0���4"O䬉b�'6�b��Y \X�i�"O��� �G�%��!��c�.S�D"O4�q��A�z�mA�a�S�<�y��	K�O�����&�hh�7�O!?���x�<��o�&"�Ȩ�ӆ����d�"
l�<������2�-P:��3�L�<I&�ҫ��0ذ�n��1��KN�<�2�ގ	5�<�Q�Չ\A%ӷ�M�<���	�%��hH�&�Sx��b)�t�<�qJ�9Zθ`�2���J��@��Rv�<s�H<���K�O+���lh�<A��K?�y���>xu��3���`�<qp&�}� p��'�(��-D��pr	��^XXb�B�z ��ǧ �hO���Y1�W2a�ҼW@��C�I,;�n�����(�){�$R�C�3`���`�9�x3AŶJ̐C�Q_
9��/�"l�d`�J�G8~C�	����$��{z%�Zhq�a4D��p��9܍!d@�2�����@$D����+�ISR���#S�}i�Up��"D�4;0����qvmO�U�Q�G�3D���C[�?���aSd�9?V:��2D�� ���P4A�hԒ@R�>��y��"O��S�Q��`�ϗ�r4i1"O�i� �˿b v��1��R�t1@�"O��%IH(pR�@�)�<j~�P"O�kc�E�J��@��CI\̰!"O�h���yEr8�Vg؏ g!!�"OzͰ���)��|S�/_�}e@�@�"O� !&�A ̒��F�0�'�'x�Br��*l N�j�+��"�J	�'�䢵��fp+5���^�c�'q�l�� ��k��z�n���(;�'����&�ɿ)i8p��-� �n�I�'g�d��5&R�J$�@�@�$a	�'[,e	� G-\Δ�bS��3�xIX	�'&���J�6�B�[�)�%x/�-:	��?�*OƵ��f�>4?t ƃ�ێ�p�"O�ӵۜn�0�#š��V,�f"O h��JI�N$݋¡�!M�8���"O��x󤆥�z��b	4M�A	"O���*A�X(:��� 1
��g"O��C@^e��8�"��*(B5�`"OLH���'p��d� �2�*=�S�'!�O4H�t�m
`�8Яx��M� �!�Ą�G#F� ���	B�ءRub;|�!�$A0����L91��H��j '�!�I��I��dʼg��(
�jV�Uc!��3�^9���@�0�gQ[O!�DBG�V��s'�a9��P���pK!���]Z�d��� @3Z���Mx!�dG4�l��&��a0А!�l��&�!�$Vv�:��@�
��x��#{�!��ɾ=P�pr��U%��1��+t{!��
p���S0%�-v�VU�(�wd!�D�9*2�� #�4����^51u!��0`�����3�2�z�%�:i�!��ٓ+�pU��E-��#2E�/a|B�|2A��q��Y�.\���(R��T �y�̓0>Fb���Y�MUP-�T��yRo�+n!r�%ƽt�l�b��-�y��T*.�a�Z�:�(�CU,�y���:�f�y���3J��zR ו�y2���rv�"2N�����L��yB��TAܼJS� �}��-��� ��0?�.O"�a &��^R�AP��C�1��Y1"OR��ꙣ_-���"���ꩰU"OĐ��MC�1�d�Shښt�za��"O�Ȓ�� -��*�F��u��Dє"O8������\������1��H��"O,E١n���$@�I�1��q0�"O�@�ЭW9 �@��&���rV�'l�'�D-B��Dk&��0�&_1
 �'��H �<R��P�%�5+(�Y�'����3ʈW��rE%�(s�1�'dS��N\�If��) $x��
�'��t�ǝ �r���ƹt϶�`
�'�L�J6._�^�^�BO�=}}�|3
�'�JM0�V�x���jBGB�_��	���D͂3̺m��RMB���3!�d؂,�����C�M�����)�"A!�d݄J�ȱ�P���0~HA�H³=<!�1�����$$�98��^)-)!�$ܭ��p���z�C��̙X�!�O�|^���l܅_�2t����2$�!�Č=I#أXh)9 �q"i�O6�� *!�1kښ'b�`G�JE8¨�6"O0���I��H� �o zJp� "O��)2NC��bM�, 0��[�"Of�rK	K9��,�.9�M1��'��	`y��O�H��j�l����{ �!�y��iV�\(�?
��kE��5�y�,ʧ:Kr�JJH9ze�p����ybM�""B�Є�1~���3iѝ�yN=h���ON�i�t����_�y��	�R�6��tk��Z�4 @3i��y��&X(�pF�*� =s�%S��y��_F�Ru�d�\62؅���y2K�nԊ��5.A#�7�߹
_!�$��<���7�G7(Bp��K؇\!򤗳m��I�&̅4$�aj�=\M�C��@h��0���}�h����5��B�	<C�H�z����/,�S%�IX <C�ɳJ�h20��}���R�ݒ1�*C�I�x�^ċAE�+v��&��U�LB�	�J��D��曙!5d��U�E�h�B�ɖD	�XA��cN]�ª��(U�B��\Q�1Qsj��@>��yA!ڎG��D���{�	Oe��+;��n7D�Hw����c5���'�T� 3
6D����D�B�P9@qi\��͐2o0D�|
C#@GH�����,�I E0D�D!���L�h�A�(^4��Z��.D���� �#e�6�)cn�<ޠh���'D�P�e��Q���8r.��G��	7�0��<I�V�F�}�j��$i{���]�<�p��.S���Ch�S�$1�T��@�<y���(?�$9��
` ���@C�Q�<�0�SQM��9�P�y�LH�G�N�<���ƍ��G�=�����d�r�<����*2���� �))��Tz5�Ip�<��*�l��T�ī\)��X�ǌSm̓��=��j#]����VX�$���Mf�<	^��Ts0/�8R��� �U�I:b���ɂi��H�֋�3Y"�`��@�B�	�(��]ATM^ �D��ȓ5<�B�	1}� 㐀X�m�Xʂc^�3R^C�I %YJ��T�!�����-u��B�	�͸�˜aC>�͕�~�c����	�vAْ'*1zt��ţӔH������?E�d�'rb�`Eh�'/�A����Dﴉ��'�Z|4���$cnX�D�8;\X���O�u��
�+4�Ĩ�*�+~u��B%"O������xhLI�)v�4��t"O����G��i֠,*$(�cj���"O������"`r��Ǩ��V^&�k�"O4�(VE�`"�Lʥ���f�騀��TE{����i�.`���\>��a׫�$S��2��hO\���E� jB���Z�V��T;C"O�9��ND�&$���i��m��{""O�h2���W`s�\�9q,<*U"O�1��ȑ�bk���� �A���0w"Oڌ��H^�2�"Ȥ�؏~�1G"OX��㒁d$����I �:O��%A�
�C�Qt�TT�&/�!2���%���IM��:.�h�e�Ŏ%%P���W3reC�ɔj8��s��˖K(�hG�T�9x�B�	�c9�Y���^���L{Q�ǖǢC�I%p)�0���ʑk��A����Pg�C�ɬa7<�
��]B�U��"�=�!�� �Q(�d��U?���Xg��D��"O|�ؔ@E��� ���S��&�Xr�'��'�t�:&LmS,�*v%� p����'،���¾ @1�¡�d�pɛ�'`���ǀ��3�лr͜	d��'c 8B�/��V�ⱂ���P�[�'d��1*z�ʊ>,����'��p�A-L[	@pC�2�Υ�'l	� Q(:H�GÃ?o��Q���%�'03�=Ss��}� ҧåVPF`*O��O?�	�U
b0@��8q�2�� `�0B䉾n��\z$��Rݨ%
�yI�B��u�#tA��
�z}+F�޸NM�B�I�	
��5�P�4J�0��I��B�	�"+l�@��_�.�#h��?�B�I/�t�QǍP{IB!��	�B��䓎hO�D�7�N�0�(^���
S4]�!�DJ�}ʵ򱢝qג〉�<,�!�޼ba ���J���iQ3Ԁo$!�$�����Q-��!��{���2!�ĝ�}�z=��C�?H�ޘ#V�l�!�֛:6&Yq�fS�@�BŘb��2D1O��=�|j5烩d����(ΞE�P;'�[O���=y�'_���\gK�7O��0<���DU/�4X`V,��HE �p2k;}�!�d%oJ|Kr�N>��P
�?U!�Ѥ]v��b�!G� �U�D�A�!�d'$��:G*L�������ے�!����,�c�0{c@�q�Æ
5!��I%�u�#V5NQę ��/	a~�S�|@��X9<�C���>kS�����>D���]�P���)$2ٲT{��9D���A�̳b|��S&���l�jt�+D�pss`@2�FZC�z����o�o�����䉉�>���D+JҝA'��]@a~�V���1 �<���%�ma���do$D��Ȕ�Y�w�ba��œ �ƽ�c #D�l�E�/�T���6`�1��6����8z�����ـmv�y�#$�soNC�	��|���LL(�]����1�B䉪c�0�'L�7�z���1\����hO>�r��Y͐��Ǘ�hlR4�EF&D�|��ʜ"h�1�c�@,'�ԒW�)D�|�1�[�o�aS�l�t��貵�,D�H	1cP�M=��c��LH���My��'��D �	��Lx�k�""��'��u�R%��4��;�n�	..�[�'u�y�ܽc8�,ʡ�@�"��D��'����T~��x�! $Jf����9� ��D(�	���eP�����-:˘A��"<D�� "e�#y�p���B/o2����;�d���5O4�3WL��.� &�ԅrTx���>	U{�̤�f-w?
�JG��j�<Y�-�$��D��t��T�U��i�<��ह��������V-�I�<vm�1w��$C%��.��@�}~��)�')4<��q��D刧��hk2��<���ap�,4j�BE\=SD�ȅ�X�II�F��bj�K�e"ǴO=�B䉴%�x��	*3�@p	�톀ZbB�I[�69@1c+\�:��L%F�vB�Ɍ²TS��E�b4d�ޒ.�VB䉣E>�ؓ3�J�Xd�@ڹs�@�q������s�끝X���KA�
ΈI�++���<E���� �T¤i��L�$kw�	%$�Jt� "Ovͪ��6DD���9A����"O�	�t(�O���V ��T[j��"O��$V$U�2�AB�2I�2�"Oj�ё8�x���;6v	G"O�i3I�y��B�n	:h'^��Ā<�S��yR�N
If~8b���3hJ���$	�0=	����/ h�挍�X��p��}��'C�e�'�2���w����
C�?�� �S��y�C� �	2-��9G0�3P�.�y"�2V�&,q�Q�[��dH����y��VF��!뙴^H8��F�	3�y�(�*L�p��u(Z/mg$Ɋ6���y�e_q8)Za )g����ֆW�y��C�U�D���m�]��\��fҍ�Oz��DU��^�B�ً8d���2�!�DO�Y��U�=���技�'4!�Y�4���a�/�j.�$�EDP5(!��ֹ�B��mM~�\����Q d!���*]�V����_.}���ɱi^�!�EOa^����S-c�.]�B\>X�!�" 
����&RI���s�v�!�$ʚ/��� �40.p�oՉB�!� 7"�������C��:N�7iZ!�8L5��Q�AO}� 9Wl�5}�!���	Ipr=x*�$I�4�[/!�ŻF�XhӇJϕk��y�`�s�!�,��͛|WV��A��%Y!�D^G�]ˆ`�q>���.J.<S!�$J7Z��m�t�K�IBX�k�+�D!򄉪m�z1p �\�),�+љ !��枈CBa�8 ���ēoy!�$�� <���
�.D��,��s!�J$1�\����(PQ�7r!�SJf8��܀p��C� �!�d��!i����͜<x�𑓢�Z�K!�$G)Vڐ��s�V���r+\r�!�dI<%;����B�$r�����T��!�d�2J.U�$H@�ffl3���M�!�d��8�&x����/tN ) p.Ðj�a|2�|r�� +�Fљ�m�:#��T�v�T�y�-U*��TJ�%#	N11���0>	���ф8҆H�ק��q����B�ƕJ:�=E��' �Q��*L�\>�����#���"	�'n"�� �\�7,ư��CX*G�
�'�b�j�ǝ�@�&�
�h0v��	�'^����A3�h-�t��!n~D`	�'7��CF�?z)��
�aG�f��tH	�'��"�cΎ%
� ��׾4 �	���h�(��W��zm�!��#7�!�$��S-��
UΨI���YH!�(A���s���L|�*�Z;&!�� 5h��!�%ddE�%:.z�!���(SU��a �2]�04��pp!�D �o�e:,@
fJN$��7qX!�D�`Ӛ���ʅ�A5Tq�0�K<P�!���OFX3@Ą.o]e�Q�;N+h���5��Nx�$;b+�+pR@�`a)�(|2`�%D�`�Í*�6� w���,r"�0D��y�ĳS�f-C6��=��@�ģ-D�d�q�G�Oj����@�j�lp��,D��qc��N�v����o�n��q()D���OW#;π�Rw�<yd���(%D�Dѷ���-���P_� �k�A6D�� �|¦)��'@fYy���+���Z�"On�B�ݨE �а&ŏ�Te���"O(��6
�6��5��xP�!B�"O~p�VgU=M{�՚A-�B!	�"O�83uf��$�4t)�o(�-s�"OH�;!�C�I��q�ɉ�}�|t��"O�A�,JP|�j��l�i2"Oʍ�r 3}��2�\?m���06"ODxrpL�:p)����OX;��L*�"O�Ѐ̆;"�^�T/��$�er�"OZ�eoW�J o5<��"O�ݣ��7�$Q��N��,Ш��"Oh�i�Z�(�KE���_�h�`U"OƝ����A�p�� c�-z��93�"O
m�tE[�%�vD�TO���j,��"O�%kЎ�5'�N�07oֲT��"O	��B�`Ii�$� ?�	��"O�Hj�h�����x�B���z���"O(�P��*o<����PoPd"O�i#�D�i=�6��>9ի�"O�����O�~��`)v�Y�^�\�V"O�(�G3#��q��G c�ii�"O���)�<A���ćM&'�,m �"O��pl�r��qK�%���@P�"O���lR��V)�G$��.s�X�"O��)b�l" ԩs%P!)W(ՉP"O�t��>%F��R%܎��4R�"O���I�xdb'T��p1v"O��0���.�f�hT��8�h�"ODi ��3m����ǰG���"O�8�CD�v���c6�ؘ8Ժtڲ"OF5�$��)��A�oP�/��X��"O����I )	���퓼Z�x�@"O��'�M;���!����%_�A�P"O�q䨍�_�|�(#�d@L���"OV��B^B!R�xS,��NzR"O��k�ʒ�H �U��<Zm�� �"Ob��F������&�k�!Ӆ"Ox�#�ϋ�N���#��S�@�|�RE"O��!#�3j�+ץ]�c�|x�t"Ob��/	�0ƌ��7�S�&-c0*O�P'��($�#&�9N4���'�,T�S���Dp�FF�rb�
�'v��ph�R)VI�զ�m��M��'�1���#6���ի:T�,��'0^]��
�nbX4��BK�t �'yb�5(Ib6��t�Al�'a|0&�� ']>�Q��?��@�'�|�:���A�0Q'���I�N�B�'\|.��=z��@]̒pce��y���1�r��`b��@���d��)�y£��=%�L�'�ζ2�pّ��Ǆ�y2$�5l�0�2�OWq|d��R��y�mә!�<�۶�]�K�R���!G��y��/8�A8�KOGx�4⇠S�yBC�z�4Ц�R�=����b��y��4g��ܲD�ު8&��Ä�Ǝ�y��z�L��`! �6P���Ѧ�yb,'�|R�k�A�|���V��ybl�gǆ�J�j���nX���˱�y�+ƾHʜ;&�U-���S����y"&F�熸�W�
�j�90�L���y��P�+��|����5N, ��
]7�yr�;~�j��4"R�0&}y����y
� �:q�O�h�%��׾|�z�c�"O�D���
:�Hs �I�B��"O��C�ã+OD��v��k��p#�"OT��S���7�VБr�:[���Z�"O$�+���}|p���۹1���S"Oj�n��h�Ћ �)�"�*"O�u)�L�?/n��!A��|��0{�"OҀ�dY���UA��\�)��K�<��MX@����!�́Ɔ[D�<�a��5��N�D�i1/PG�<A��I :5� �a+�J��B��B�<��)P#(P���)�;<|F< �b�z�<i�	��:��y5Hմ#&8зH�y�<ɱgч!P����O�w=�K7\p�<�,�0@�K bͶT }+1��a�<�f�Q�B��e�/���C�_�<)� 0j����]��Rԛ���t�<����u�ƥu��B焐C�hSp�<�r�@3�hɃGH�<(S���d�g�<YÇ �$�ґ�Fȟ'�`�����a�<��az�� ���^�:��T�<�R�Uu�t}h!��1"�B�� O{�<)QjKr=,xh�������Dz�<�QF�R�8�a]w���ը�v�<q���{O�|2�-X�P�4%FW�<I�&�]Ɯ�D!өav:�j��V�<I2,�!Z25���>�vl��(�J�<ɖ�ͳ��ɺ&�����qY�<�
�n��]!#�[郎	vo�b�<!�n�>8�r0��X
����Q�Z�<���p��0ء��|Z� ����U�<)��� �B��FC� �~)�V�R�<��K�5[O�5��iR�kr�͠s��M�<�D��)��Iɇ�2nVYh���N�<�������U�V��/`2��g�_M�<!2N�}�ܡ���GL:�
��P�<�+�<�.8�ЌC!j�� EgEt�<Q�� �?�6Qs�fM�	�c@�K�<Q��]yAQ �!BP��E�<��O}xqx���B��Y� ,~�<��FW>v�4��V,�T�nQ*�
|�<�����nO��0GC�6�����#Is�<)�iP�hM��x�4"L<@BWn�<q�Y	���á�&B�R�`eO^i�<��C��LX0�C��r�%��a�<�S� =^��! '3pGt(D�S�<Y`杠 w6�� �;V�*u1 �j�<��aψ^�@M���̴Uܔju�k�<�p���/f���\�1z����P�<�Ӎ�[lQ�D�<1�� �O�<I@Ň �����%�a�'\H�<I��Ս �ɡ��9P�T��A�<Q�B©2�$�ڷ�,�j�I�@{�<a��9_��p�D,I��U�!�x�<� kʾL���r!F����iV'�|�<a�Aƒ<?�i�E�p~�@���N|�<�ph���T�����MU�4��O|�<!�@Bq���AnƀX�-�6��w�<�vN�m��u���M?u�Ep�/�s�<9B�
+��q�!�I�%H��p�X�<�4'Բ+� �c*�'��<�F��^�<��ԕ	���3W#^)�e�v�F�<�W�˙�|8����a�c�UD�<iP�/2��9r��� !d���K�<� ���h[,b��va[���4"O���ᇖH� �hB �?u�f�"O��JbNԶg����ԎN�mn�"Op�*F���!����m��񢤚�"O��"�]���pB�S�H8��"O��#qJ�^��5� aВ�l���"O@�!
^� �``
7oҘ��� C"O+ nܽc\�H�B���3"OH�a�I� d��m��&���"O�t� `'n�nY@+��hn"P��"O<�H��� z��t'��<a��D"O�a�f��'d�#7�/9T��"O�R�t��� rK� NDQJ�"O  �BE��{���>J���1"O�(�[|fm�B,<.H|�B"OB�z-A�}�reԏ$\�9+�"O�=�@�/):(uۗ�ɅFA�	�F"Op��R��"1�ڡA@�/΁Y�"OP0��A�H����@�܆>!4�Ɂ"Op@�p��	Y��7O@7<��u"O�����ϭm��Xr��4�d��"O�]����(<�C�C� l�|��"O-)�KD;L����#Λ5����"O�tCŬ5�Xhq�6���"O�#U%F�r�Ip�'�8�2�s�"O0�$�
P0`∏����	�"O�i�E�<0�^ɵgB�\٘,y1"O,����-�^�8�N�B��!�"O��s����}҅�-_�<�۷"O�����_�-̚�#���V�l���"O��#�Bct���&�}\b�+"O�%ZB	|H���D��@s&"OXɐ��֯.-�1aj�8�5"OX�R1�.y"T�2�MR����"OxI���ݟrr�!C���X��́e"O�`�#]�f��zӃQ�C9F��6"O68ADٞ>�ܒt��
�l��f"On�	GiR��&w�Pc"O���������tۑ��I<P�ȓ;��d��Ov��Uӎ��cb�ȓ	@⽱���9J�V�jʁ'"a�ȓe�Jꂡ�%k��T2"O
�B^��ȓ-�T�h�!���A�b�6U�Ї�B���t+X�:lT���ӵ{QH���1R t�3l�Gܰ�𪁮2l�=��Uq,)��M�}�jJa�J'�� ��UK���2#�C�`��� t���NX�V��Bp���'Q	V��ȓUD(سp�'�e�6|bf}�ȓt�X�4lA3m� ��HF����ȓh��4�T��=��4�P	[�~r���ȓT���&�n3"��֣*�)�ȓ25��Q�������B�N��RŅ�$E�� G	H�4���1N˗J�T��F>yڇ,F�*ϸq�0��':���CV$:!�UB�褫4�֥ �i��S�lq �%C8(d�
ş2�8��ȓ����K��Xw�?`��]2�k5D� 8C�Q�u����o�F1���/D��`6�0WF�=��R;.:w"+D�d�eFʝ
ʄ����*H(����d'D��K鉙r0h�+�7����#D�,�'H�m`�Iդ� ��I�cn7D�d��'I��mܛ'i"Q���4D�� \K`L�'�BqaBM�
�r�rt"O~����+�Rq�P?p[>�X7"O��娎��"��J�nq�	��"ON$b�@\���fj��BU( �Q"O@�������͐`��	 =���"O8��3_&s�:1�P�C�;*v���"O��"�n�?F�`�;`ϕTl���"O��7���=r�ER��
g�Tt��"O����ؤ!�BP�SOύ��;�"O�E��o�g����OӇ���B3"O�Sūד-��a��̒���u"OP�rC��?R�x)!���*$4$@"O���A!��|���#! ��n�-ڣ"O�P��C�t�b�ˀY�m�b�*�"O�a�쀌�b��2e�?)X%"O��1bٿi�b�C���w3��a$"O�'��Q{��!�e!���"O���֩ûrJ�IQ�(��S�"O\���n\�1�D�h����B�@@(�"O��95��(6�X(��8G��"O���@��ܮl �k�6e:0V"O���i�#2�
� �K�~7f�P�"O@01S�ҝA���ڕ/�,fͲS�,�S�����m,C��9G%x�\C�	)7㠨F'	�z0L2 �:	d�<�	˓mc�a��"6L�-�6'�6`����3����kT3($A����,��P�ȓ
oڰ8�G�/T��!�`۬I�|�ȓs�҅�M�J��đ@�
�H���#�������cnl�P�j��m�<�U�/�S�'nQ  ��ןd��0��O�KJR@�ȓ\���G�;he�E�"pEy��'0
ec��ښx�P���H�*��x
�'�&��`�d���`M8*'P�Z	�'m<��D;����G^�8�T���'>���aKɛx�&4�u��/��D�'�N����<
��a5�P.v��:�'�@�'N�+x�� P�ÉiiH���'���hVeC/�(
Q��"��Q�'ڴ���(8h����l�8	�'�0���� 
��:dǍy�T����D)<O�)rvG��Zv�6ȁ˂k�,n!�$��}kE�6C_����6e!��?J�U��C�2�j��C��SY!򄃦z�`�HDV�n�6��D�*E!���B�@�/�2U�n|�0.ȑ 
!�D�	Q�0�2��B�������,.�!�DD�~����N���O_2�!�dǃ[�T���KL�I��8�S���t&!�$�<&��ks܋%C�u�u.܇M�!�dB7r�Q�d��+Y^T� �O�Eh!�DI����@�+ة<h�)�W�֚QQ!�dZ8sy�(�*3]Mµg��X6!��T��PXi �Ae���U@$��ȓ���T+W�NǂD� �[k}�q��|��Yh! ��F&&}3��ڱx�X��VN� �Ն 5<��h���{�"u��'d�Pg@E/~r�� ��17�M	�'D���'�-C�b�0�"��}% 5��'��]Ӧ��;f�0�ҏ5o�d���'G�Ļ�C�{0�)iG!�
�4y�'~ၠd*@����V����6u��'��<s��R�:V�t
��1y�z���'h�UI��߆D����%D�(9��� � �T��r'��9��[G#h<y�"O�� Pi�u�##L+�}c"O.<�E��#0@����!	(����"O����(͠K��QIB��93����"O���w��m᠅��6��`J�*O��� �K�6 ��MP5]�ڔ��'�m�0oP2��y����X�0�
�'@v��P%�M�Õ�P@!�
�'
�H���[�D�R|���:w�|�;	�'0�q���B�2X���#�v�h��'����t�(=6�B�����`1�
�'04��BO
�t�#D.J�o�.e�'�(�@uc�:l0�����6m�΄1�'�T���Y9 �p#c���n��p�
�'>j%�
ĝS�ܓ��F�c��
�'hĄ�1��(@k�=;��_�^�x�'�j}�S��n�=��Z���'�r�����_<0B0��{��(�'c�4��݃[j��B�R�b�d8��'�pt����7N���6!�Z�r�H�'`�85�zl��f�Y�B�[
�'�^�u�͠-q�p�YC�D��	�'%(���C�<c�~�{R���L����'(6�
A�[������0�X��'[�Ғ��S�\��gX&j���'�"��	C��Q`#Ƅj��#�'�bL�lЌ~�����%ex����'�
A�����,�C�NX�8 	�'��<���X2w��Yӳ�R�V�"Dz�'��	�+�}n>A3Vl�GpL4h�'�.�ig�A�V ���U-��<.����'è�QG_�8_���f :ˬ�
�'Ԝ=i��X,%b虊���wa�M�'Ȏ��a.�?� ��V�l�r��'ؒ�ȅ��v��AJC'�#i,>i0�'ª�1�`H�Un<P�[�N��'�4qȶ�{�@3v+�C�\�
�'������\Xc5l�:
�'�l�hq��Mqp\�e&[3��iY	�'�N�cW�ٺ6���;U�V�-r�ġ	�'�Ld2 '׊QS�)�QcW�=DD$��'J8x�1��o�yPJ����HG�<�A�_�c�,�e��`����7 �Y�<���I�C@)yU'	�h8�SA�M�<�����`�	 %%��!P�hEF�<ar�_�1�r$��nB*AG"�9�F�<����.����MD��q��[i�<��BA�8IP��V͘���0��h�a�<Id��v��At�L���8��]�<�2� D@ϖ5n�T0��H�U�<�U+�u̞0�FĖ쮀����h�<it
,l���0o�r�n�b�/AZ�<i�g_3�J�2 ��7ᖀZ"J�X�<�G(A�l����-Y>dRz��+�{�<�ˌ!&La�g�:=�`:0(�K�<�� �C�D�t,K�6Ț�)u��G�<Q��C2;��qI@�0�j@��J�<!�E��3�-��:�jVD�<�a�׈Y�� �@�����I�ah�<��F�lY��A�l�{���e�<�7���@X��FO�$�Zei�{�<�mp&MbF��Ym�m����L�<��m�9Ԭӧl��V�f!�&A�~�<�B�P��t�dK���@$�e�<� l����J�4z`к�\+�����"O��ԭ���	��	)���p�"OV�	�c�'F �W��h�h�"O�=q���?��`�y�F���"O�Q$��:,lHė�;�����"O�|X����a"!�aT++��-�g"OX�bDʄ87݀�(�"Y
�Ԁ"Oty�o�P��Dܙ�p�R"O��P�	Ү�C� ��N�~MX�"O�TP: _�J�ZM�K�bv!��On�2|3�$�o�X�����bh!�$B�0@B�%��~��!�6ğ�kV!��ϗ/���C�#�C�Dq01`4!�DK�{�TA���E��J���AY�"!��u�$daˈ;Ĉy�qjԻV!�d\�t��3�o��?Ӗѹt(Է�!�Dϱ]P~mڥ��*����#��
'!��&[R�z�J؆`!DU�!K�1!�,C�t]q��^
B�w�O�H�!�I�h��M�꒯5�l�q�ճ�!�$�:y��d�X�wʮ�Y�`û|�!���)�����!:� =PD/ӯo�!�d�� ⒜*!�@���I�	�M!��.�Z4���͓Dd�܂p���'�!�d�&L3�E�
���>	2��΂g�!��W����a�	�9��d�c��I�!򤊧pE
Ic�iñe��%�w��6�!�R�Xmf�hQ�@�'I���#Ȯ2U!��AD�q�k�W(p����A!��9�F\)��hK���!�"P'!�dH-8P4���fi`���7!��YR5�v�T�;Sʰ�S�^�!�d
�E������0s>�y�/
�!򄇟O���� �Lɮ��Q�]e�!��$i�lM�!B����m+�l�I�!�䄦�� $+�5c��ݠtb�8ag!�dπK�(��k�H,Fd����~]!�F�E'rep㉩;�8���`��\!����\�1T慴�4� ⯞�I�!�$I@�|��0��W���"R��,!��*���q��ݠt����ia!�Dؙ<cD!QQ�ֵWf��MV�jL!�$C�"��)BTe�(4PqyC5M-!�D�o^����
4f4 P8aAҎsvў��;�ʈ�EA"4[Z������C�I�J�����5��ٙ�'�)2���+�I�p|�H˖E��}�s�G�fKB�	�x��xI�Q$Va��#�҈��b�E{J|2����'��`���_�L�&DO�<���]�A�y��+�d��Y���L�<9Q(� y�zQ��2��	q�^�<q�ŦQ.�]K`�>/�]q@"OW�<��#rD]C#�%)5jx���V�<���]������'%ͺ1�Ii�<!� Y����˗�؟P�����@���<%>y��ۓ-J�P�f�L�۲�9�-#D��a!�v~|
C��n2�إ�9ړ�0<�QG�0=}X� #�t$�䀥�U~�'�?a��[�N\�$�gU�LKo<D�����{	nq�F풿 H�D��$��@��ڸ'��aҴk�.XfI3G��>!l�q	�'.Α8Wb
�u��WK�|J�'*f(�P`��#?���!L�'\�,����)�d)�f�������N�	RbS��y
� �)��P"#`���%��)6#����x��)�S�Bm,�І�<�0�t�܃S7�B�	/Q�伺�+�;Oq�a"n_3]� B�IEsvp:��^��>9J�B�X�C�ɟR�ޭɅ�ʥc70� �g^�,<B�ɗX%�|9`�@YJuY���*CJB�I4q`:�
�҇7.�Ȕ�5l�TC�	<r���FF�� A�88�<���y��)�&�A̽�f�	�V�L�vF3D�`B�Gf���UE���5D��b�
�&��-�3��<��*5D�|k�cǙv��9b�8E>�!�M2}b�)�> ��4�����Sx�r��t�N�;����Oְ�6�˻R||��V���Fl�%���$7lO�� Ao�5�r4�JڈoUB�q6�O���I�/	~�yJ�	_*�!�&�,!��mt\���j�?��蛳Gۀe!�Ą;4�"9�4ț.���$�*	 !�ą�-�⩣b�ˍo�h��iB'�!�O���a)Di��&(��o�!�䂿a썢�`F�]am��W�&�!��p�Fh�(O3$��ʆ��>,@!�d��yo~S�LM��ԁ��	&�U�ȓ�`���̉M��1���hq�ȓz��PЪ4��(��m�%vɇ�\��l�lپo��hb	H(�(�� �h:���[,�[�� $�Y��kI���`mܐQ�9K��ۤlR���Pֺ8�̅!D|b!�gE�L@��Ɠ_*t�.V�6���j�͟9$6�J
�'~I���=�H�g�!'�
�'}4��F$Wl"@C��!��l�	�'�:q��I�p�r��Q �4=�l�1�}Ӓ7�1���<E��N��p��|+�aKC�� j�Q�<��_�ȱ�P�P1$��f-�S�<�C%X�"�ry&X�O�����Lċ!�$�2���#���<iJ��	�wu(����'k�����ָ.q|�+rڜ;�`��'��E(�*vֺY񁆏64���C�}"�*�
��ѱ��� i�Fԋ�<dPB�I�6����EфK.2�A*!�"b�F{��d��7z�뇁C$R�I�SH�~��'��L�q+�(ò	��N�6.�p��M����i>�&�@�c�X����{�bӫ&Ѐ��E7D��	O�wc�Q��ăh�t�0�I}��3��=K^��U��g���a"��0| ��00T^��耿s��P���AܓE���D^�O8�SulݧM�n�R�	2#�B�>IO���'%�$$LM�n�;6Ks	x%���xR��:�c�m��UJb��f��$�yri�,W��Ь~xv�1�Q!�y"
�f�t�1eB� t+� ��i���y�����>���`�p�� ����y�AϚ}�:��a��:�F�B�Eڑ�y�B��ly�i�"^�h�H�ْ��y2Ƌ�t��e`$�Sh��Tqeh�y�^V����#
�̕f	�y��E Zve���w�8�b����p<���D.~�@ ؄	Љ�����Ư����Ps.|�`�ťq�L��S	R�q6�d��&f]['�Z*	+F�BH�+B�,qD|b��rw��S�"��
��I��C�I
zX�|Y�O9K&��7��0�C�I7ph@��P�Z�5�e��2��C�)� NYPc�Rf��t��A�f8�S"O��0b(:G�\	d�Y�
|��kq"OXsĥ�;w�a�f$�[y"= �"O �`ņ!����%�� 4���"OH��G^(NA�� U�.y�$�'ֲ��I����'K9b�ZH�F�&���A-8Q�#�Ϥx�h�b#�*)BJ����k?Q���Iv*�w�H�^ܼ�ғ��l�<�f+�3&԰�$�,k8�S��_�'DQ?��6e�'w	\�2���4� z��)D���gHJ@~Tv��4��$£f'D���1ɞ(��i2*P�+c��r�O&����>�C���O(��+�3�$���"D����*�:bƂ�x�AV/��� "D�d�'�Q�uȢ}-���P��}���p?	b� [� Z#�MK�|a���Pa�<�e+B����q��O%T��䲆��[�<ҡ�$?'���G���$;j�R��~�<A�i�* bT1tǝf���j�Je�'��'�>��4kH�uHP%a���\t��`+,D�[LKe���C6�Sh�j|�Fd����z~B�xJ?牮wХ��)
%W
I�#.�%V�>���Or�>��}2�\� ��R�ܣD��{�aX�hO6��dL/�����A-I|4����6
�!�䐈nXy��V3c�����B�?����>�n
�8�F�ڥ��%i��hr�+D�H��([�Y�Jջ�`�nҠ���*�P��$pN�>�ࡘ׀��v�X%�E6�	U��ϓ7��7��X�|�3�VK�Z}��l�"��QR��H6��Q"0���'�ў��.��)�x���=_�Np��e/D�8q�,Ah�{� d�>����?D����ަE�"�Cdk(�!��!D��Zu�8im<�H�lRE��	K5!2D����`�<\&2MȒ,P�gr��b�.u����I,Hp�����31��ؒ�Q->C���M*B@�U�I��ɒ��C�I��r]�g�\��*y�Tf^�#FC�	%z;x����� � fn8~<���>�E�E4k�rQ�֎�48�@��G�
I����p6O���$�Y�Q\*����3�b�I'"O`Z�#R���+�%�8��]r"O&��4�T��P;e�\6i��0"O�L!�݋T�%
�!�"M�=�f"O�ܘc��H|:�!��	�I �"OX`��!�qMr��&� DuZaX�"O�$�����ydc^#	�qx�"OF���)[zN����#�ƠR�"O��q��H19�t�A�G�w�Vy'"Or�J��(�@���JӾx�Tв�"Ol�a㭆0n�L��d��])Hy�d"OBpx`o@��\��Ӆ�:t ZI�p"O�qeJߛ=�(�C�#B;Y��ӓ"O8�H��ԡ2N�1�-�����"O0}6%�C�lq%��	�!��"O����ᐭbW&H�k�r�乲"O,� �X�BDU3��E�ӠP��"O����75�\	�@�
�p�d"O4�Y4���+�V�B�mZnHXX��"OФ;�����88��+P+���"O��5��<�tMba,��`��"OlZR甉^Rp��*o�pAb�"O�����7ה����Y
u�2��"O�������\�~��v�?c�Z���"O� p1@��P�P�.YB�X�p!R6"O�鸡c��QTqI ���v� ,Å"O�h�ANM�(�*F�O�F�^�"O�E����h��  C��|a\!�"O0�����]����B��c��;�"O��JF�W�q����@�����	S"O\X �Hx�)�!S|m�"O�}ӷ�)'"v8��;,�AB6"O���Ӛ_�F�`�L	()��\��"O�Td\�}����� QК%%"O���-א>��r�KY�.�pa��"O�t#��;4��B�
0�N��"O�D2֣F�~��]�'(��0"OH%�u�����e�J�y�H=�6"O�:�E�6'<���,99p؋�"OحQRQ�b4�� ��-)�a0Ff�"�P�#�
/n��DԞv��)2� �|Jy	a#Ծ@n!�	(�z��4�z�Ic��Q!����0-Ќ6�ڌ���B�
M!�H _�|E�ס�AĆE��a>>5!���
�ܒ�*�P�*��fA�Q!��.�V���
��pʡ,�!��X�����C'��$��Ab�K<+3!�W!,��\��*������D6�!�� b��,bQ&�?N��h�$�2z!�@� h���8s�x<s�M�*Oh!�P�*���"��=Ǽ�r���m�!�dZ�
���K*�d�b�lV�!򄃞3���b��N�zFơ��E�8�!򤝔r� "�B�Q0�ň�C�!���O(�`'d�(R?�q�A�FZ!�dŞb�2�Z %0R;*e*��]�X!��
Ҋ��F�7.2�I%�[!�!hiBҁM,_����GR�/4!�䕤{Ur!"k��{��y�ǅ �!�D�e6�KP�8s���F�>�!�D�8-,�"�Jie����%)�!�ʿi�J`P���5ZJ�З���p�!�d�;k=���W66zL���]M�!�F!Z.U!q�O�8k��3��S�l�!���/_dMcu��(!H2��'(�6E<!���)Mi
U)W�Q0��@��B�!�Q�d�d\�g���p9x�c@܆�!�DC�3��ٓ3�3!�P�"���w�!�d@�TR�(fB��� c4�� c!��&!;�*aK�I���s��O��!��&�&q �Хv|ғ��q�!�Gv���{��_'nR���K�'�!�	u�,�e�,�X|P�i�$3!򤈟��M2�O�I�8��Ǖ�:!�Q9����e��>�ޔs�Y�!�DB$FqBQX��L)�nɘ�ʏ!{�!�DQ�xA�E�d\�K�T��U�̒:�!��:2��eqѣGQ���!B�)H�!�$�3P"F|��RC�^�����!��&MBP�����G� �3��V�!��էU������2�@H���%�!��\�ؓ�M�^@�m����S�!�$O&b���B����n!�)�^U�F��'ҠM�!�Q."i!�gL�0���2m�	ʮ+H!���0�!��쌽s�|("��Q;!����$���p%�=7��;V$�35!�Ĕ�+�.����H.�\�&�E�*!�� �<��Ń�`j��:���4/XP��"O� ��"�� �F�U&h:c"Or�Z��U�#�� ��
���@"O���g]%`�pɐ���DLS�"O�|
uIN�Kྵ��뛺(��H2�"Op���>{6����0�&��"O���0X�
����8Qr���"O��D��3f�뤁ͬ1n�yp`"O�|:l�?K̈ ���o#.-�"Ov�Ҁ�)uo�4`��I!��j�"O"�b�*'N+ ��l_�>L� !"O�бWㅧ@��`J�*K�Q�"O�h0�锵L�v�hAJXn~� �O`�^��I�d$�5� 'J�>���ӂ=�'ð}/X9�w�ƹEKJ���w��0��3`��P"�	��^)��uJ���mS�Z���Q�&E�P��bJ�*��N�W��P`�W���p��{�}�����pRE���]�؆�<���'ل���8 ��4��ܔ�Z<�&(��!�a"�)pFA�򫝵a�~�a��W��l+��Ҕ+��]���!�Aש�6=r�{MʧN�<#>�b�i�2e��ǀ�q��O������)E�� �	�0'�8��'_�<
6H�?S܀+����X��`����`M9 �����5�蟂yRƢ	�U^����	o��єA+�	n�����'��	cpkФ9���w.M4E�����X��?�kN�|��X�!������>c�4BS��7��e����D����"6����dU�Bw	yD�׹i2��[#�Ɯ]��xS�&��v��Ц��97vh���'�H���6�ȭ�3�N/ft��h#�O�xl��/_�6���M�b������5�B"=�$b�.M����uf	3R�H�eB}>���	@�7k4#�"cJ�0�E��U"
�Q�FS� �b�X �Lxu 4n0G��U6n�ѱٽ=�9BnF:,/Pac�A֚���`C�p�h���B�����G�g�,��(�~��	MҪ�r/H�"">4�ҋ[f���TM��"�DR�"+��51V,�~�7*���#�4A���l�&����:A֙�`B�4)r�ضI��*L��kd@�?�mZ�o�4 �B��@Б��"H�{x���㇂Y�l	��5D��%K�'��k0j �u`JV�'��M����8a%���ÃBC�`��J���p�䋗�95:�p��1_���A�+�dɊ6GǄ�J�B&kP< -��	׭hv`|؁J,˚�˔�Z!DO2��!lB��(O$�k֪)����t(�#AG<��Lbݩ:2GJ>M�hk�n�$̶��B�P64DիtA�6�H|Ba,�(-�y��U�O�|C���0�Vc����Th^��jBztX�	Ӻ�i0�LO�°�ߜyĴR��$�J��dު���w��8Ã�+p���%7�=����50��a�h]�\IS��2���U���'D��
Y�c�<�f�ν3��x���L��lZ�¬؉7F��)��a�0�PƅO�7��`�D�9L��T�ȗ}ը��[!J �BL���T	q�ЌX��x�d[�����Z3sj�Ye.E0@�������uղs�A�W�Tk@d[=�Pk-[0t�t���V�O6��E�v�݆h��p���jOv16�.}^�GzҊ_��]�q��7#3� ��g��<��H�k��|������!z覹�V�׵{R �G�K�}�2��n;o�tA�W�A|�����O��K�<(��Ct��QKLV���՚e闦Y��ΐ7h�ժ��ڽ^� ����E�V`Y-\!���'Y:lx7�2V�2����!t�F��b��� �1[H	\^,R+D��~��Y�A����䔼.�j��@ۑvA���Gi~�7ʞ�V�LP�I9'���B�&G�u��,^L[��x��i��R�_�xS�T����DA�
;�O�LY���/*@����3_�$YAG<4�DQ�p�V�}D)��|�s�U�U�I�4K\L�я6TS��	P\��)g���l�г��"�j#>1��?�D�3`A{T�R�������><�C��@�R�h��*_u˓�p`R�F)�x�?٦�߀f��X�A�E�|�T���g}b���s.��s�J�ΟhC���2Yp��0�R>����B0J��Y#J9�":q`e�6�'�xh��H�8N�B�B5(��Cl���'c�a�G*+@�(r��O��z��%|�d7"?��	���#��3=4~��Γ�P��&!2� ��i�X�"h�M�^��'��\s�b�CLɧ�Ԃ@Izl�'���j���3jԃ�����'� �0
A56��5�"�Z�A��Q�O>�oC��Y�Ó@�b�9����G�,��eeN�X`D}��@�f��o"J�J@*��a�0M�Ro��/�TB�I�F��Y0N�j	�`ybh� �B��vc���J�!q���8;�B�ɵe���U)S
 ���Љ�?L3DB�I�PZXX��H^+Z�@F�r�<B�)� ���G�0XT��A�8]s�up�P�<Ђj\S���ɣ������4x�(]*�nO�X������?�<t���3���(�@�0��)7gÎ0!�`��'�j�@��8��".ҩ����X�[@� �a7r"�?�z��X�g*p�j2+T�D� 4!Ũ,D�DIb�(Q�P�W��U�4EC�`ה&0p��-h<���<E��'v��t*�w(J(�GF�W���y�'2�yJ�E�<;�ja�`�\�E*j��'X���3)�z��q��'6�=�7�ˈY�҅p�b�5	�Yy�F�)�O(��/�i	do.DN��q��]�D��W�T�r1g�8)��"�,i41Gx��M'c���
%"sP>!�A�;,��P�E��[��P�"OJ�=�(H"*.�=e'ԓt�����ӂ!8`���W�"~�3t� g��5%�
���D��u��$�&U���#Q�4x��Mj���L�z%*aE��l��n�<�g��*�k���)����G&�\bf$�/�.��ʟ_w�y��R ���(Q�B�H����{��9O4x�ׄސ#wh�0�,R�c`�IJ��{b/�Q�OgQ�6�أ�,� ����J��k�)��.K�0>1�L���p �r@��BQg؞0n���T<�t�'�IY(�w�Z�ȑ�C�sjx<��'�� �S���J�>1[��ĵu�Vt �}R�ݣ��R� �q�O�4���/k�l�a l5�����'
��3E�X4�*��7+�e�����X=U؞Y[��>���>	V�B�e3��)��3V]�l8���c�<i�DŌ	��;e�E�z쾅	�,�ᦡ�A�~����v�'ۨ-ysŇ\�����y+4i��1T����Nu���@)*���Ң���ř�N�Mq!��PD�{��#���
­Y�c{�O�`[֡YRP��I.ff��m��52`lF?Cz!��T������؄w�2I�K�mz*XpU�8n.��'��"}�'��X�1��w���4̖�&�8���'r���kF�2)��l�	��	�n ا���0>1�e��L9�x�[Q M�G̋u���")�>c_���!tf�+�jH�e&�!!B��@�!�$�L�Τqv��cr*�*e�ӭ;��ɳ��s�i�����Έ�;�(�MN9C���b�.7�O���+;^%|�;���]���5.�*.y3�a?�y��Ҋ0�,m�t�V,!�5C3)�/�O$��%
Q$f�A��4�S
R���ÆN	x��ĩ�E�6m��B�	1���UG�;yq��c�.��~t�1A�_@��w�y��9O�3f��	O>�Lb��S�l�l"O��c�C�|�xH�!##Iz��w:O8�����8j
��7<O�9B
,&�L�R�aO	6N$p��'y@�!�a��Sx� ����#CȰh�GKs�2��a��%H:��2a�.�8aN�Vռ��q!T���"�!.c��m�bv�' -ړ�Z&0���c"�DE���ȓN�AI�h<)�y���_$���D�A���������s��4KE\�*\������!�t*8D�0ʣ.M�g�!8Pi@%�I�B�x� kƁ� ��`�`�Tx���� L�B���s�L��V	@���#7�OX- �F�^�z8 s��`�^@ץ��k� 8�Ї�"�yC~����=e���)���HO�'͂� �ң|ڲbO��4��۟	���r@�s�<��(В�lU�	�T�5�GT`�<	������8t0���f�\�<1��a��pɋ5N6K��T�<��nG&��Ma�3DQ�z��WS�<�t [0�� i`�ê(�|i¤��`�<��ؾQ��d�G*��!��Âa�<6dE�i~
���e�pt�(Rrf�b�<����x�^([�ǜ(~ʜQe"^�<�.X�N�9�A�� u�c��_�<��⑮Dp´�� {��ݬ�S!�� ��&#I�G�Tx0�C�`$��X�"OB�q��\���0	�H�h�(�"O�q#G%{ߨDX���%<ľl�D"O
٩�N�c��@���U��C�"O����h[�]vb���@F58��8z�"O�����NG�Ժ�hڅ@�*4�6"O����H%C\ g�G�Jqq�"O�Qr%�t{r�Vi�rV��ӄ"O�ɚ���ku@M�VH�3sE�qU"O�����.WB ��U�FUf�p�"O�Y���B�!m,�!r�W  ^zh�"O4)i�I�@�Ly�bA,5�{�"O��F�TY���+�%O���!"O ���Qax�k�KQ����"O:��1�%:�]����|��s#"Ohٺ�J�"@[�2�"O�1���ֵY.��#I��a��"O���G��w=@EH���ν�f"O�T0@��E���(3J���>I�`"O|,҂lZ�x0��AȆ)2ݔ��"O\p`(؀ %��1P%�� � "O>���iD�_`�0B���FG��"O�U�����l����j	�1���yb(�
	�H¶�P�+F�mc�-ݧ�y�W?���P.Ph$�+��y�&�V�}�d״_Z��ٲ�Մ�y���xڒe��܃S�2�a"��y�G_�7'����8\�^�����y�J	dv�a��
�z�"Ux��G�ybF(�z���U�IK2���y���(v�Pd��nѺ��^��y��DL5���e�jT��E�y2�!m��*2I�x�h��ѫկ�y� L	\`���~�N�;��@��y"$��D��ys҂K:p���I +�:�y�@4 lZ�w�Խut}��H
�y2�Qc�:a�*B�p���M�y��"\�yA	�(���A�$���y��V�!:���vHIңS�y��JO�D�;6�-V���Ĥ�yB�.7�z웳�� �`�5���y©V�W��1�NO����D N�yR+�!8�a{�'��t�Y��X��y"F6D��z���2���eAҨ�y�W�`�<0HR�^9|.���
̿�yB�7f�Td��:li%_�y�)];�4�6j���|g	� �y��As��S� �
+Mԕ�Vl1�y2j�	i�����O�$�� 	���y���9/���E�+��qx�y2��G �	`��;,�<��*�y�Eϫ�2�X���..��b`���y2��`�n�9�K�*7O��r _��y2`P�$a{$�]s_U�w�G��y���`8�x:�웳s��=sG ��y�iY�e�0]c��C�:V���aT��y�J�%�2 �a�?��1�4��y���_��d"��޸+�D�tʁ�y��ߕ�&�
T%$-�.�tŗ��yBA�J��|�á�VH� �Å��y��H�Y�z�x �T z��3��
�yR����"y�7���>EƜ(RC��y2`C�i�n�c�S6&��A	��y��� o��H.o�W(U��y
� ��Qh�4a�!	G��u� i�D"O\U���]K���C��&rf�1�"O��2��L+
L蘒�a��k��x"O�!sj2:8�	[ª+}�h�"O���֍��.w���\i�у$"ODٻ3K�>y��j�E*� |��"OXPHD/ў:��@��S��I�"O@E�G˃& �"dA �y�r��7"O���oӪ@�(4��
m���"Oδ�V!á	�`0{q��!OY�H0�"O�l�d��1�`�0aW=18���"O��iZm�Xl[�Ϟ>D�BUS�"OjX��C�7l�7D[�ṷY��4D�p�*�>S�dܛ��+����5D�89ǏJr��$O�.-��Qئ3D� KЂZ%��Z�_,Y�T��u�7D��ZF� �D���Kԥ[7�l!�0�7D�t���X l�z"�WM�>���5D�4#�N�<��-17*U�.�AKF &D����iL4p F�1D�du��&D�xy���pG���6A�l�V���#$D��[`fB9c9܁�u��:v ����&D��0�&��y�^��,���,��T'D����޳*�	�C�e��iv�8D��B��ƺ��a6cܼ!�7D�����!]f�1��)Iw����8D��z�@иzlx3�)A:_����=D�DIb��g��C���u�htP�*9D�pȵ�В~tN�#m��C����!4�ɀB�����'"Bq"-�g��6.�����bA�'�@��d$X*V�R���c�*Lp� ���T��reOF�3p�T�q�(�Xbd�	3�n�)RO$��R���'"�
�ޑ�7��"H�����y�bȼ�b�bu�B=�qHrh��Px"$^�-ǈ��gm�d�|y�[�Zz��",ة|��txƉ�EF������-Ɔ��w�)]N%2#b�Y�`�F��x'�������ڐƋ4����M��_;j� �ć$�t����\���c���Nv� bJf���]C�� 5[���&z����
�^�D�'N��y�-�h�ʁ�O��n�ҡp!'a�꼃Diͩ%26 ���-H$h����J�ƴ
�c�J��{���!��)P�dV��EO �D��O̸b�.��-T���31	���")p��Q���Tj_�{<�Ybf��
��p�O��;�Y'B
P��ubK�,�p)�G<��IRT ũ^(�,��@��t��p��GZ������):�bl�F
_9uJPI;U� e��#?�5#��Q�ҙ3"������0}�4E��K�#�X�����ڰ���R�_�4ui��).����~���+�I<RB��	�;(0RH�OܶK�B�	0Y��U��=x�MZ�	��n���Ǌ:��C�!�05�:��3'�;@��q�3�Q='&$�j����=q��M�!����Ӭ]�9�A��U~�ʓM�|���ƈ�V�I#���d�Ƽ�t+W?B�d�h ���Ll���)'X�9�J�'�:��' ��"�t���
�a]�J�:���{���r�-�A�T����j� D3�HZf���d�'� 1���O%�`k�k˵*6��P!��$��Y˖�ɐn�j]ٖ�G(�E�lk�xS�KS2nx��&��;E�����͊T�85ۆg��hr8�Ck�,�~��Y6=����$�)T��B�D]9�f�3�hv���ͯE�9�c��8��D��5�D�����'y���pE�2n�����FE�=��v��e��G�`N���� =>��'`Z8xê�'M����Q��]�2�bL���_Iy�hɉ"��4�@�Y�iH�X�G���0?�c�K@AZ4	WJ�"f�1��kA48��JEG��r� ʓ�VȨ2���rΣ?���+M4�<���G�}�@��G~�'�^HB�iƜd3���'=�a;�I�G�NUy7��zl��pweDl��)$M�U��\;�2�8�ѥJ�-\��A3Aʳ�����̯W�j��'��9S���Y��N~*���I����Ĝ/�\ Ð)�c�<��] o�2�Gɶuh���S}R�Ј?L��3�|�OK���c#�@yҭ  Ԍ�o˺nI��a�!��y�
\٦mr���[��uȲ��;��[��a��ET��0<�P�����D����e�[P<�pH�2�9�d��}�`�[5(�r�8��1�� �£��'�<xQr'��[fB��"O�)��ߥc��1�f�sn�5*e"O2̳��Z�\P6�J��:k��5��"O��Wʗ
.(H�B�7<�"a�"O�������@�k���x�H�.O���
'���d^�`�EK�D��!h*j��|�!;����WkXWbB��P;#����
�8T�ȓTX,��/�SB
�k�*�!��Fx�`]��D2�	"��N@P���(j���+q'�*1� b"O����*+�<YԧU�h�H���f� <�l���̑Fy^�S��y�M��y1�43P41�5�3���yob����蘈4���S`�	�y�_l���(3�O�<�y�I+lB����?!���b&�7�0>I7�5��]cD�6�|Q&.�9�X԰� K�v ��C	�'���R��>�16gҷ	�%c��d�?g�(%Yv%˳A�"�?�b(�]� ��u�5?�x܈�2D��$K݅>��dCWgR,$�&�N��B��u�S��4ps.͖�����i溰:w����"��G��wj!���>n�� �A�H�(�GO�nA��F�6貔�
�~�f���T���ŧ(:���*׭�:8�|��\6\��|�@`��#q���V�Y%?�����,��02gJ�ow��"~Γ̾���a�<?ϒE+���B�0Dz�!�g�FP� 哺p�p�#BƏ)H��`��S���$G >'n踢�;�OV���*�)�p�[�^x�!���'jm����;g��ɯ>�y���'r�n�0 �M*�8C�	�n(Cp��#(��p��뉒{d8c��Z��K<���ө^��,�"ܭ?\~�B&k^�C�I�	>�c@�j���� �d.��� #O;���OX0G��Oj��C��#iuE�N�2�Q�"O|L{�+�<i|��jtcS�=���)G�imvy��mν_�dd�j�x�[�#�q$<x�7 �o�J���Ć��U�(�?�QIĬ�0����VR��N�<�F��c��x��#�y����!�s�?�2DXQ��]&��}�FDOV^HȫV�Ə*��e`q�Lh�<��"�(�"����?sࠥ"$](=+|�
@����	��H��IF�w�_L<�`	��Y�EVC䉐,0=�S)$�rl�c�T�2\$�$S�:��UB�'�O ��&� r�� ;E"W/"1V���'�~���N?�A�	;R]X���/T�L�W�J�<9Pjޭ�t��'�'Y��[TUx}"���<�:��%�'"-�H ���VJJc�qR�)O�!B�靃JI�%̚y�@��։�s_PE�:D�<�0cbm)�'�4U��)#��G�����v���fr��l|�P�`�lx�;���/X�b���B�8M�@I�@��SF1�2�L�	��qQdA[9���s���򇊄P#�2�A��\hz$�?D��p㘣E�F�A5MC*������f�0r4.R�,d�"_nx�xp�k�"}ْ�B���% MέQ"�O*P�D$��e��te��b�a|���A�r�B�I;�f���˻l?h��4|��#<�֯W�z2�z�����O��p����Ey�` �pp4��'���h��[Dr�T�G��k3�Zm��r����4}��)��<y�X!K�Q��B�9ot�y"e�Z�<	�_3p9Z���Y�cl
���U�<	�Ejޞ���.��<�Ť�50^|�4j�+u�f ��l�H8���A�_2['l!yЈS0SY�Pj�(Vr�ڨK��,!��*6jdjf�|x@u�҉'
��8A��401G�4�ʶ}$D�BdL�r�qʞ��y�)i�	a��B�1��!�y�BM�`�zC����� ���yR���L��qL��U��7�O8�y�m�5z4	n�\�{�nd�lF�yB	Z�M�@�f+�3 �~H��G%�y2Ș n��5˲H�KiҤ3֭Ā�y
� v1�!%1*�>Qv���a���(1"O �! ,�6	
<�Dg�|E�-�a"O��`D��V	��b%d�,59r�+q"Ox�"Fϒ�6��VdK� Z�+&"OڵR$��y�^�q�DO/��'"O���b��j��U�b�D�H0��"O�i���ĝrBzXr�Y,��q&"O��J��M��NYH$��4��"O*D�����Q	��3�H��1"Ov�#Ì12��x�W�F����"O��Aǈ4@�Z���,�@`�"O��
H�1a�H<j#G�,
Ɋ�D"O���D� >&�hH�/9H�ͳ�"O����D�B��0K�+7�!s�"O41I@�ߙ!$�
�+ �hH��"Oz�f�O�R%�+��l���"Oz���-Ә]�&�W
5w���"O㖤׆g	n�+��T�P�=��"OC�@T�9q��TC\��"ONU�a� C��uk���=6\I�"O�@Q�S�`,:�(��68E����"O,��֯΁����`\�d;���"ON)��#��U���e��E��e�c"O2}�酜͂�z��Էx�:L���i�@�1!̉.p�V���	`�`r�H �4q��	!��m䝡`�=v�4��W�X?'!���0�� %h�M�t����ȭ,:!�$��h��ٹ��)!5ģ��\�!�d�^�����Z1jQ�b�!�D�)c7(8�u�4|Gdc��E�uW!�$��Kj��%�#M+L2F 4SS!�D��j4��`ݻFdtd�ȧ->d(��XޭK���O�l���fݹ�T�'�|,�PEt3胢E)Z�l��gⰈ�yX��`�CJ�����O�$4��BB	\���L��C?
8h��B-,4��E��š(��iIa���שG�.MT��1a��e�cʞ�j�t�Zm҅CQ"	3��];�䉋ç'�pXA�ʕ�Li ��ߚ � }[R��V�TI�� ����)���v>��WB�.lt�u�Â?��D���Y{!��nڹLtP�b��є*�X,�'�h�RI
A��9:�1�62;��f9O��s�;��p�8��퓚/�"EH,V�N�R0�Z�[���q� ١�����S�O�y��%�F�81bٛm�J$�e�'X �	��y<�-�uN_>���MUa�00�ȓ1E���Q�G�F�
lZ@�q�ɅȓsU�d�u�Ȓ,Vx|;��/�"��� �Д��
J�v#KU�.z����W  y�(�T֮9�$�x�t��0D֠8�+E5[8r�2��ɂ,#0���nV��Zw�ѓq�n��ܼal\E�ȓ=���D�>'P��%�Rh�R�ȓ��z��^�o���jCI94Hd$����H��BC�r���@ֵW&��ȓ=(�@��F=U|pr��E16��ȓ|τ��咖_�ܐ��n�y0�=�ȓ5�nJc$˸2��-�5I�12��l��x�����^<R����lֵi�(�ȓ+"X�X�.F��
4'k�}r��ȓOj���K�#F)��/��]��o���� �QY��j���DJ����m�(���%D�j�T��2� ��@�h���dO
%Fn^��XG�E�adB.|*�1�A�}BT��F74�صD�,#�hq�5�C:��,��8��fa�8��06m�=w�B䉐c�9s%$è���Y֯
.j�C�	� �� �U�>˲,�'�ȤC�)� (��b��+q�� %���S "O�x�p�d�|i#5��"2��@�"O4�)V�S(+���*�.��"Op��� ��PN²o���f"OJ�Y0��]�T(q,ñ"�$!r�"O>�` +Ř|CP;4�ƣc�T�Ȃ"On��Gh�`�諢`ȗ�H;�"O���K�*�~%�↊0�B�8`"O�|SA"'.�Ah��В�ΈP"O(�:B�^��� ���8�z��"Ot���<Y��@���*5���"O2,Y��4P�[e��B�UY�"Od�&g¬s�Vl�Q`ϒf0�]j�"O�b�F*{���zW���,�T��"O�Re��b���^�V�UC"O���A��$��,�7Z�c�ЀI�"O�����בB�t YQl��֮�W"O��@�a�s��-��J�?)��A&"O��դ�<�Ѕ���Γ �p��"O���Z�z��TY�f��O�TpH"O����\4X��8���K�x|�]�"O#��>?�� ʔUf٣�"OB��'˔�0P��/7S&,�#"O`\Yt��F$A !ĢP[���E"O����nf����1eO�і"O�Q�ѫ�n%z�!�RZ�Ժ!"O���glU�LWԁ�F ��o:��"O<����<���I��ZN �;�"O�-�2�XTf1�"	�Q@���"OB�RhÍ7Q谀3%��p�Ʃ F"Ojd��&�<Eh���`8s+��it"O���r�͝)P4� �@}�p"O�qpVǋ�Z� ��WB�>@	�M�"O&p��x�QckR�#��<�"O<-���ZA1�tZ
�;+����"Oά�A!��)��y�Ƀ>�~)�"O P��?oOv�aIC2l�J�"OrI�P�ƑYH*EHW-�T�"1"Or�P�� j�L�A�B�_��B�'[�ݠ�kո.@r$�"��N���
�'\V�X0�3�Bu�E��NT�{	�'0f��既r�~j%��w�^�z	�'eH07�K���[� 8h!�M��'yd�2)<�����=[JNU��'D01@iA7�p�7��b��8�'�ʄ3�&�����Ĝo'2��'��@[�ǛN�x�A�I�k����'�]a���N��p�Ŗg���Q�'f�(e$R1�����d��JئY
�'�reI�,��QڀY��J=E��A
�'ˬQ�sk��{�4�1W��@�'�<�%�'��@H�*NlR h��'"� b�X�Ԛ��T�2kܵ�
�'��)j#m�-84 �(N���-��'q&U�G��5>@H vk�B!rYQ�'�tU�$F�,XR�b�h�N��$:�'��m��� S����턣T��	�'߾�j A��y��SJ��s9Z��'��j󣒐4��\��!�/x�N@��'/���T$  r�ݨr��<b�	�'�2=����#��x��ϼ?z���'~Z�Z!#�4Z&��1�F9B(�"�'���֦�ˤŁ�倍]��  �'��<�`$��t���)S��H���� :��aA��k8�@5�]�>�r�C�"Ox��BL`<xtbvg�S�j@:d"Ohٱ3��yG�
cvp%"O�i�Q2|#�앇v��M��"O<���mR+i
��`ܺ3vQ�"O�Y��MQC���(JYCT<J"OV8 �h "		U�;(W�Ex"O�6�V>gJ���v�Oؑz�"O.��3m��Dؚ����$2�0e"O���F��ͤ�	��í��Qل"O��ұ"V5S�@d�gI�O�
q[w"O��C�j֓t�`e��t�P�A�"O�D�� �o#^A���N�,��!��"O:a�
5[;x�I��V�.z�w"O@��%a[aq�0أaɕBUt�Z�"OƩ�b�
4�Ru5��s> ���"Ov�A�W�"ɼ���&ԥp��ѣ"OrM��M8�p�hS̙�y��HJv"O���k�H��H�0��w"Oh�IaG�᜼"���h�U*O��S�O�2^��y&�H�c(��' ���Mr�&u��Ӷ\���'e6a���+�R���J]T�l}I�'��	�-ݨF��!�J�b�T0K�'uRXx���Z�.��,�^�TC�'giR3�#1d@y�.��!�H���'�v-��MY��D�D�Þ�jd��'$D�"���&5-��j�!$b����'�2��'�ӜTt�"��V�"@���
�'��!qr̉�5���X��9d�d��'&4�a���uOtT;C�I& �x�'�b�!�d����b�9/J���'m��h�N�/Yg���ď{J���'��(AI��m.-�,��"OΑ�bo؋$e���˘o����t"O�=q�JB!���C�/�"Y�n4�"OF!aʛ
]j���K�����"O��Bm!dD���M
�8���"Oz	�eh�t"h�p��<�6ey�"OJy��Ϙ!j�.0c ^�mr�&"Òb $Q��0�@ ���X�p"O��AЁ�w�����B"��9�"O�����8�� ��Nԯ@�\9"Ox9j7�چK���#[7�D2q"O��(�Y{b�+BG�U$a "OjQ�Bd�"�(Yw ��3���T"O�4�`�,xs� "���
)�H��"OX-s��)9�p��τ?��-�'"O�Ԓ&LWPfN� ?�"O�Q���(r�x+�,U�K+�Z"O��I��J3u*nI��ׯiT9��"O����H�e
�IA��Z#���"Ozi� Du�ܢ�闱?�T�`"Of�@ ��"�n�Cq�<o�q;�"O�j���P��!8���=V�%�u"O,b�O|/������H�q#c"O����	���KvL�%^J�Q�e"Oi�gC�#R�#���7-�C�"O��Q&E]9lU� 1cȶ�Z5"O��0��-(�b��&�ۊ�1�"O*�	0�(C��M[V�X�{���W"Ol�"&$NW:���F�/vs|̓�"OL	c�]���`�>m,au"O��j�M�%q�J�s��:S��j "O� \l(��=���׋/H��cg"O��R�"���IF�C�0��Q�q"O.(���G*.9��@��Y�n�S�"O�|P��I�a䪑{T	 w���PG"O������(E�ڬ.B�c$"OJ� �o�t�a�lQ8 9��"O���CĀb�VY@��N����"Ov���[Dg ��&	%D�f���"O8-R�B٨hI��0��9�`1!"O0Y!"���v��b6�R'n�R��"O�-[vC�4#�Є��%	{��"�"O��#Κ]%&\�3�ƀ���k"O���a�q����J� .�����"O*l@�ą��Aϒi���1#"O�,��'F�-<hm��#׫9�켲�"O~A(�ҝ$c�{1X�p����"Ov��� J7����=-�P��d"O�(9UG^�DR��#��M
���"O��f �11�����6M��,�yR���ߊ����xH���J�1�y�%��;�Qۂ*�[zm��T>�yR�FU3�ڱ�˕x��2W�΋�y���BkD�(^���V�۶B�p8��rKx�.%��y#v3��a�<�$d�����g�O|ABqk�\�<���>0��Ҁ�2Y�P�d�m�<yp"ą'P����T1`�N$��#@g�<Q䎊�2	J��f(0y<�Q
�c�<	���de�hӵ�V-{�ƍ!��ZI�<1��@�Z�����,N���n�H�<�3�7�d� �_̼`!�D�D�<	��mxU���,#6D���K�<����cB"���ӳ�ҵ���^r�<I�ᐴB��e����+_b�5�j�m�<�T�L�%V�ȣ���l����l�<Q��A2_htq� E�D�X�����h�<y5&N�������].Z�����LI�<��f�B�:��[�9S�9��`@�<Q�f��.%��C$����r��}�<YQN��'��DC���q��x���D�<A��"�f�� �?A��꒩C�<If��s��9{v�Y0��H{�<)��]�/���$HǗ
fq�mEv�<)I��_>Yp�`P�/
���h�o�<a" ]:��|�2�F/>}1��[i�<)�ˇ {���k ��	dpa$��d�<����_X웱'�o�<�h��^�<y���a��H L@t���Z�<٠)Cr����!�ds���U�<)F�8P�����?�Ev �P�<��.�M�0h%%��T}Px�v��F�<	$C�8�\�y�+N<*�&���E�k�<��2N<�`N�L�c��S�P�tyw�r����?�}j��?y�46�2a ���搉t��+;�4Z�_M���O
y3��L>)�f�3 xE����O��V��!u��#��=}Z�l���U�U��Ybw�;�ө�y�/�"�lTP�� Ѥ�bd`�=�d�D�O�|m���\��>���cj^����������+ׂ!��W�����1.i�!'e�!T��e[�θmq*�'���^�m�ן0�ڴ��I��|6�ؾ����Ê�Zt� �+){����0)t�<l�Ο����%������C�P:1����!ݦa/d��֮�
?W�e:��<Xj�@Ō��z����$�Z�nڼ&�h)!�v8�\�l	�����Œ ��B��^rb����d'�����T'��P�Q�h��Pb�#8<�"ƌ�
ېx"FעY��5b����#��b��$=�DS����Iwy��) ���)� p��Oφ�j�j��bf�j�������o�i>i���da�՗��2�� �L���(v�v��Z�G4lO����A@�<�6��	ĶL
T%j7��J�N�T2tj"j�8t0�p��e6�Y�ҥ�	ڟ��3��f��`�"|����2�*faJ�	wyB�'��w�O&�
ҏK�̉se�D�v�%�
�'�FlR�Re�c�S�O�bmR� ږ�M�۴�?���,��&&?U��6��O:˓���Td|��4�[�w 4i�lݹ��O`����W��Ob��+�	_I�P����)���[ܱO������,O5���'3�'�+�,Ob�y�b�%���)&��.{�2�'��O|��LZ�h;�&�+B�$���i�1ڼ����'�ў�NR�M��<��ɰK��
��؟`N�z�Cp�����>���/P��0���(m����I��@��2�MaӜ��<�O�b�'���i�<�A�BI�8� ��}�kbj/��O�b��L>i�nR`v��
��W t���Rɂ�n�fy0e�ĴV���i�'U#}�'U��
��[5*�r�L��1�,-�S��O���W`y�����R�r�3掀�U~q�� 0N��`��c�"�'����"`��ICx�9$��6WH���{|�8�oZU���
�4�J�``�1C�����;v�<��0�X��i���'��|�O��vgG"(�������u$�mq��Rwwt(��J2�O�1J!+H	U�"Vˈ �pH�`�ij�� "CǌP���X��'X�80a��/Q�́�@:&"(��4&X��ٟ8�J<���?H<9��@�n.� �f�XF���B�X��-�O杓p<dqC�G�EQN���dޱ�M�O>��i��d�|��c�6 :  �