MPQ    s�    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h��G����|I��+N���
V��I�S���a�г} �7	M�9'�,x��0l���,���:���e�w��k�$bK��c5�i��xt�e�MFksb
�c�]�,8�����){+'DIt�RiC ��д�^�W�tx�I��[� 3W���w����߻� /�	��i��UJ��N)oJ\)��L5F�S�c�"��-@  �N��OL�k�LI}mrA�v�c���6�������!*���H�w��&Y�t�	�h�\�W��F���-V�ύÅ"/>^0'r�+���ch��.4���«��CC��h!*�ź;0��������t:Onm�1�ƪ���@5��/�D}�Ä��vڧ����P��6�������;����7�а~���c"�S��(Y�b��{F���ݢ~��C�o�Q'@�+	��"��eO�A3���e|�ݭ�#pi�z}l�O��VB���y-uHFV�>�,Cn�ћ�ɺ���͝4�r`�z�@���7G�v������tw�-����ߧS�==tV��U_Wz�ê�
�^��������i{�Ma��`r)e\�z���`l[�R�(A�(o�RXw)�)k=�{t��S>�0�L/n��5W���F���mC"/�\�� E��@�mdI������*,%�0+8�If4��&���߁-]iy�\ϛ��4n沜*�2*Y��U�����r�U{�$��7���,������{8eYP�@FZ(�ۖP RE*3{cDk�=���K��QRp{9�_Y��Q�Q�s�;;F��wR\g1Y�7����ע�i������x�\�g���ů$=MO߮I�2r��nչJ�-;'Rws���۲��=��"�S�m�1�ԙ)j�Ki�az9o�ڋM	��7��_�{!A���Ԇ��P~5g?�2��[I'��%�
�I�Fb�+�qZ�JT�K17?�ɟ���m��#+��}	ċ��]�#��V�O��kY�ᨏ�^0]7ӕ=��i�^�~(QF=e�uy�#�L!Տ�����&�z�͡���t�#����U�T��@����7�Oᰴ��q�B�f��-��]/�\ W�}�݈�8P�>`� ,���r��Mj�@�X��g+�º�������-ç���D��]���pQ��l�AP��}=���v�6���Φ�wb�.l��/�:B����Ʌ6�\&��8�ǰB�%cDΝl*�?�#p��I�8Du}�����ڸ5��H���D������������������~��:Nf�i�8F ��Z���FV4+����p���k�c�pu�i�QF&j[Ħ�g>Uam�s%Ň�xúHތ 1��r٪�|�i���a9����V�9~��<A�$��Ie�*h�y7QII��iwDT��l�M�����WBշ~���-��lKps��;��Jr�����h�cNA��j9��[���.����g�|gӷ��oT�DQ�ET��`�f�O�L��}��%�T�ǖ��WgVW%A	�J#å/[̷^�]��0p�g1h;(gS��I�J�3mH��^D�xa��W����o5G��)	dP��18��f'�Y&��D{�1�E�]����.�C�hۦ��3��ĕ��ب�fäna'
����D��H;x P��]��A!��;RDgNEX�H�~~�%��l��]�]�K�G�w�P��ry_��E��0�Ӏ��@ �m��ʀP\�|}	=��A��
,����ړ��wr?Q�'*^?���ˊ���]l=���ʜ��5�8���(O�+����޽Pߍ@q���D�<	E|h�X��T��S�����7EZ��Eݻ����<(�J�Ry��$���K��[�D]Ԙ�"���A���g���'�&�z������e�4��^w��Ӽ�0�l9,�!^��`yl(}q��\�h/hfb%C"���Q�b�%?��2^�2��|9�E0`��AK�I%=]+(�P�RXK���=8 [�%���:K��;,<�����s�TQ�m^Ix|fk;��>��{����)\�����GEa��g��O;ppi�_E���Tl5�?1�'��*
jfl�g��F3\�k�M|�.����I�:�K�l)!X��C���FUҥB�'����P`WY��9>5����QH�ƅ7ӣ#���!�]��Ǻİ�>a���O���V2Cm�����"���T�?"�#�rn;~��?���2^�����$�:��w/�/�-��q�,�x �ߊi��m$��VP��1�څxH^�N��@	�y	�[�V}x���o�Ȍ~��k�ُy6�/@��V��I<ڂ���VO�[5.�鏠�|t��� Mb���E}�9���_ܴL�OY��b����{����P��U)*�h;xdŢ��8��67�'nX���ߞ�°Z�8��zV�'e��߮W�D�9T�*N�k�
��|D޽]�F�O7��Ê!��or�u/�����@�NK�-�`�@��<k�b�L�QNq�'rգ�b�v��~2��Na�����0B>�4�,�[���ʗZ �F;�m���bb�ņ���VM��kb���T/B���k���y�a�W�Y/��{�z�NKލ
��@9�-?׺������q��|
8�}0o)%ͷ�SEV'�ؽ+:݁xv��%��`C\
{b8��k�����|[΅�93�1?�SS߾B&��o��<[䧯q.gL�*I�����FX|*G΂]�0����¿琙Ƕ�NƲ��Vj�J6Sx�9�<y�Ⱥ�7�0$3����E	W4+��/�������YA�0�?�wq!h �S630�#����}��y�����s����&�����m+�I��堮z����Z9��4��vp7+�֔�Y�Lk�����_�=�V��D���D�Z�a5U:�f�)�ro�=²���'�'��2��]<-�!e�mx���te/���Ѭ��c��/�'���j�W���P�7���1��)`{dKn���ZA�7�Q-�0�գ�GDʡ����d����j�0o=��%=�7UP�<�L����әV}ӑ΁}�Zg���[iB��qU3��I_��ւ�_W<�J�W���d
|}��7sm�r�$j��ߥ]��F{>��Yn�(�(�K�$捓g�/q�icߋ�oE^&j���I�L�{_Y�����h.crА����&w���UEL����JО����5�#S�@Ћ]���o� �q&����kѬJI��)AF��c�3p6��K�_��!%�пb�nw_��Y��|�hu?�W�6̵���-	���
"�!3^K��~�C+�Hc�d��ɤ���F��AG4CC8�!E�r��
;L�Z�|ʸ���d̗Q��O)gq1�Ě�@yc/ߣ��^�5Ր)�/W��FU6�*��u��B�;��|��_��c���������/�݈�VP���c-�����oH?'��Y	��B�N�&�#emݨi�~J�5�z-ƽu�p��qG�u�88�9^��H��>beѶU��5f@��ƾ��vz��L����GG�V���e�.Мt���]�~���?=�<ȵ�1
W�ʪg���y!�}Y��4�'QM���`mн\6o��04�{�C�����}�c&�R��$��N-D׶0�K�L�eW�>;������h��/49��h�m��ʋ�#��
�%��8�Qj4��Z��H�My��<�f�Sn!��*lY�hs�\+j����p��$jǬ���<�ڼ�q��eT�T�dlZ� Ζk@�E�Vc���x��Eh��y����{�8�YQQm��s�y�F�!�|P1T#E�s9s���i��&�1��x�E�g$ ��J�q=H��	(�2-28n�5��;�s��N�v���8��r+�S���1��.)�=KDZ�So�u�P	��S���Q_�;�A�X��|�PY2?J[�+(GD�f���
��F}G���?!%��Klgj�� 1��&�A4�+@��	�e�,#�8������ᣅ���@7���t����(,�jx��u�.�G�A�����ؿ�޶��w�Ox�#�����u�����;�8���c����A.�hǊ�@��W]�W����S�S�>���� ws�`�M"=�S�g���:L������TՄÂ+���]9Q�pL��l�ͧ۫������|(|���z�Nf�b@S0��/�穏ɠ0�\�M���$�����%��Νg��?Ӓ���S)}�\D���Y�L�5�z*H��NDގ �ms�����~��_�~<�:���i�Q�^8�ÝR�� 4�I��Ԟ��1�.��s�u�M���tj�ަ �U���s ^���w��� ,_E�g�7j�i�\�a�N���zV2���B�A���ߤ��L�yR�L�H���|4w���VM�4d�JudB�'�~�<�-,�0KKփY��CǍ�������c	�A���9\23[�).0fM�RO�wB ��<�o5Q����y`�V�O�7=��m%��c�� ](�VrM��#�@�[�	����+y�����;���
���3H��6`3����R�L�J+qGA��)$bh���I8��v'3f4�1�J�8����`�R.7ؙ�������3��̕�㨷8.��r���_� ��Ò���M�C՚܊|�6��g���{e�ˀ��Go�^O��A ]R ��B�0wW���-��u��K��[�x{X�m��K�|؛*�c�%�P��?��ۄ�Y[�r�闡"(z?�H��3��W�l�B~��=�b�5{N���w�O��ǟt�ػ���?ܫ����@��E��X��T��<à{��R�ՙK_ûx���w��J�>%y��~�𑱚�ID�8R��v��|_�����ҩ'ݏzi�)��DSe3䠃9G�7d��d0�a�,�����y�?kq��Cy8f��"g!�QW���䆧Xݝ�'4� �� %އ�ч��]&������RB{����=��[��2�����0>�75��s���Q�ERI�W�k�>�M�O*�)}��t˳��ga����/vpK__�Q��%-�5�+jׂG)*�@'f�|;�37��k�	������@�c�MK���)	F!�`�C�&�V�@�""ҟ��W��9Y���g�7H~�,7v��n�a�دa�g(3>|[����_���C�j��jkĸ��&��9�#�u&V�~��<����>��9b�5ވw�P./~�2�����S �����m�w��Q��H���@��y�u�bt�T�n��~}Oʐj:�٪���٪��Ѫ���dƄE΂:��QI6O!��\�骦L|��E~�A,E�7��b_7��
��}���:��;�U�0�h6R�d ����Hͱ ���<˱-P���*ZC��u�Y'�#�i'��_�>T?���F�]���y�V�ACd7.Wf��EƊ$�u��o��?�ˉ�S-}�>@
��<o���݉l����6����v(22TYka����f̶��ʙ��,�HǨ�~���Z|��X�m���-SJb��i���MZ��k=O^���b>N.���h�O Qaٵ�Y�ʋ{��~N�J-
m��9Քj��F�u�\q�1i�vd��x�oK��RU|EQYA�3/�:��v��%�C�{���������$�S[���9N
�1���S��&�0��qk�����gmI����^�&XW'�G	���'��z��B����N�7�Ѭ���S��)�׃�ȵ�ċ!53�[�ˀ	��+���Y\���
Q�TjW��`�?���!����d�0�!��b�}Lh����Y��s��&mՙ��m��+�ݬ��C ��ߜ�:����O����4
�~���d��!���g_R3CK��__�FT5 T���Uծd�$�4ox�J�mk~�B�B�i���8���e��Tx�̻tq�,�f���3o�	��
�
�M�:j O���;=7!fn��u�D��d�^j�Z��r�=-f�~��Y�G�?p�o<M���A�N���$��=z[P���L𕟻�\w�q��I��5����l"Ba*gqP1��Ǟ��1m<NF�2� �P����g}�Ǘ�c
ry�+��؟]!�{���Z�`k7�(�-$wÓ"�q��i��>�hƑ^a���K�I�ɸ�֫[�X��&7��$q���6dݟ�dU@�1���J�8�V/5	!�S��l�� E�c�^ ɴ�qyk���I���A��c��m6����Jl! �ڿ�ºwtMY#�u�u�hPB�W$�ŵH�-�x�C�"�%�^f�����+��wc�ͩ�d5]����Ԝj�C��!`R	��;���J��S�����旬�JO��1(I��wK@�|�/#ƍ�1��ԧ������6�f���G���;,�H�m1Ұh�;��x��W5�X�1���:����C���to�Ж'�>�	5�������+/��e��ݣ��D����(*a��wkۡ!d��"u~K�4���m ��2��=ɰQ��3ɾ��zmQ��dG��p��E��I��tm��8����=s%R�-�W0�p�"�V��$��ڥ�������M�:`h�R\���˃����t��B�������R��\�o�����q-��f��L%}s��Dڷ+�<���cݨ/�5>�\�پ	m	؋��b�E��%�9n8�y
4H�P�P�c�yx�V�A2�n\��*�Y�[M��}��[���$��ߜ�A��1ceO����Z�)$����E ��cқ�^��=�����{��Y8.�Q�N�s�׏F"�_��Q1Own��ǇM �i�����u(xiN.g_$���[=C2��d&Q2��Jn��@&�;ݙ�s)/����3ˢ��T�SQ�B1�+)`��KaB��c�o�	�Y?��C�_GwA�/��|6/P4)?�X���?ɷۚc
:��F�	#�gEi �K��ɭJXz��j�����+���	�� ��s#�fi��Bk����ល��7IwV*��T�U( ��u��1�Bê�Z�|���-a}͗��*.j#-Mꅋ����x6�s����x��p�g�����Σ�@�:DI�R�VWC
�S�V�n⥄497 ����M����N��g�s7������:Q�Ϝ]�]����1]�*�pG�6lRz��f�ӹ�%ױ�:�ӧE7���bۗ���/z�!�dR�ɻJ�\����1��&s%����bP�?pv�_�n.�}R��R�P��5%�zH�B�D9��(L���|Q��q��:O�~w?�:�Q!iҊ0��˿~x���4����J�lK���d�u~Q�-cj�֝��OUW`/s����K�~uE '.�(���i��a/#���4Vmة5	�A�8B�����Q�ym1�h�����w��բ�M��d�yqBK�u~��#-�F�K&�3�����cA���B� �c�,`A�p�9��[x��.kf5��V�r=�N��o��'Q�ߜ��`�f�OCӭ�P�%����L�[�X�V����O#y�[B�(�G���&
��r�;����=|�W>3#�q��®�}�M1��MG�4()?�����8��6'n���̋R�_ޟ��#�VSv.R�7�^��K�3�����F��*��$���1����>
7����~���wv�1�g�\6�2���
V�p�ӎ�]�}�=Zw�?��>�?ѵ�+��6P-��m1s��F��|3NX�iG�@v����}�C�����rH���Fr?k�D�w��0�Fl3����N�A�5�Q��`�Oq¢�����F(�6.���e�{TE��OX��TJ��[l�my�ƘջS]��#J!J|y���$���汵�"DS�W�؊F����Gq$����'8z$I}�Аe�����ԻIѩ;�]0�v�,ij͛U�_y�v�q��J��f�O
"nKQ7��P����BV�{'���9��5���t�]!^�� RΗ��=.T�[��)�����`�2����sW��Q�=.InS0k�l�>���)����+m�aטG���p&u�_�"���%�5}7����*�7�f�J���[3JZk����dQ��sܾ��Kag1)$��!N="C̒�<�*�ۿ��}�V�WϷ�9t]����HY��7Ih#�	�����:��>���EF����C�g��������p/#s�qR��5�����y�o��X�0�@w��/9i�<^�"�� ��J��mZ���L����,������,�����/o�Ѯ}�4�e��4c���҈���,�%"��ƿnV��i�L�mO|��������|jn���^J�|B{E�=m��MO_���������}�̻�����R	U_W�h1L-d{��Ӯ�q�"1�M�ˌ���7�Z�;��p��'z��$o�z��T���!���"���<�7��(���ƥ�iu%ԍ�m����L-d@�<ʿ���������d��"`vc|92�+`a��J���*��C��7d�,��t�����l�|��m����cbq�О���MՎ>k�����r�ڦ!Zy�
��a�3HY%�{�<$N�ր
Ғ9���pA��0��q��tr݀ϔto�7�����EL�����:S�mv�h %��C���{�\�ݡ���� 0�\+[D�{9iI�15�GS���&'� �(��q�'�-g�? I����e�X2DGD��f��-`����=R�N����Le����S�dm�r��Ȱ����^�3�DW��	M�3+��,��*��Q���O�ȇ��h?\?�!�ֽ�I�M0�?�
<H}�h��{�@��z��.�z&)C���Z�H:+�čK�֠����U���,1�jr��l)����
TY���z���_��*�_��z��������	PUp���Xso�X�(.�]�������29e,>�x�1t��I�!Fg���ٹ��J��L���j�fR��F�7|Ж�9��_�dAo���ziϭ�}-¥�/?G�Ԟ�*}N֚E�������_�c=�XP�^LLKVϻ{(�����Į�3��oB��ZqK�S �Yd1�L��<���꘧�4��q�}�3)z-r4ȱ����]�6{��5���&fy(�/{$�Hؓ�k�q)�i�Q
�C=�^��jE�I����1^�x[�A&DY����Tq���:�{U;\)�_��JF�u�,05�>�S��9��h���.� ���`3GkG�I�\�A<PWc~�62|��%�!����fw�wY>S�����h+e!W_3��*-��>Ϟ��"`I�^���t��+��7cWc���G�߮���FC�u!{ع�A/;���މ��ۼ��b=�`sO��1C��Đ�@Ơ�/U¨���J�$ܧ�i�����6��k'���;g*�#���@��PI3lX�/���ӽ$O�u��O��
��o��'q!	P�8fQiPuSfeM�ݞ��4_BҫNcCGĽk82�|��z�u~��/J�=�	�#%��ES�+]��^�;�#��z�
N��j�G�g�J���d��t�k��q�X�w=.��zI�W�$��ݾp毽�s|\��u��fM2��`c~#\�m��>4���g���ùT���dR)���!6���,J<��;?L�����ki�f�{�E��^Z&/�Qk����$��m��q���,À��%S��8��F4���5��~�y�d��"n��M*�1�Y�n���گLs��zV$`����M�| ���eJ��Q�ZYrޖ��E��c�\.��I4�{37��bK?{j�YSyOQc�xs�UF]2#k1J��) ��_Ui��z�'o�xDwRg�h�ŀ'�=>q�߿D�2��!n&�U�j�;�m�sd~1լ���.��(��Sl�10��)��K��+�Kګ�	�.��H�_(A'���PS�?���a!i:�Ƿ6:6
���F����j]�r�K�']���{���ʼ��+�Ж	��[O�#u��� ��<����o�(7yE���U�(�2uJA-�=������N��HL����n#h�h�&W���D���^h������8��� y��(n��g*�Mk\W��s��[U���� ����#�bM;>�I`<g<B���Y�䞉�J���8�|��9N]o$�pB�Hl�FW�!%%��tS�rm�ӂ����Qbv���	��/����54�ք4\�(�؟^��a;�%4S��]=?�*Y��SΉS�}��+�s*/Ӌ�N5�ϢH���D�	��DI����
����~�!:�;i��	&�9�!�+��4����ڏ��4p�4u uyuIb��j�� �6�U�	�s��;�)@��� "��䣋�}i��>a�U���qV��}��/A���Z���[v�y��{�Έ}��w���=CM��� �~Bg'~�j-"�]K�����y ���8�yo�cg7A�9R��[S:.��Q�~ymX����o��Q�\��~n`x�%OKn��N��%ɦ�ǧ+����V��`z�e#T֦[}�������!�(�xB7;Y��!�3�y�����I;}�H�	� �G��#)Z�����8{�'��l�g_�����V��E^.m
��`���'�33wY�S	��<��;���6!�鹡8���޹#l����,��g_Z���ϩ���������v]�)��8�w�ʣ�a:)��AY��-�(�m��P�AUD|� ��$;o�[K��y$�k���A�r㞭��F?Ʋ��2e��K��l��c���|^�5���|i�O�D�=����X��<\�|~m㶧WEMJ�XݜdT�[��ٿ���D�A��.���]J�uy6_5���|c���~DD�a����̯�I���]"'���z�����Oe)�4��R����֧�0��x,�>�� y���q���l	f"�څQ7&��v�Β��]�5�����nj�pR��L�])5�a�SR�����=�$�[jep�Zl��f�-��a�s��Q�U�I�nwk���>A����e�)��*��(�8a���%#p��_�b�[>.5xc0�8~�*;N[f�8�1Y(3�*�k8���Բ��}��])K	:)?�!�9�C��w���v�J������W���9�!��]\HH4K7�z���vJܤӯ���w�>��Z��ؒx�wC�����ϸ�q��PȄ#.��������y���oM�+�w@5�/�6 4�����m o'#mm����G�&���pڶ"a��|�X;��
R&�*}I:�`���;��G����*�Ѡ�s�t�i���r�p���G1�O�qf����|�w�����緖~EN۽��x_�������j���������U��h,f�d�N��i2��=+ʩ��I�g+�H��Zy�f�k�)'v����&"����T5�����3�]|����7�a7��R[S���u�	X�H����kz-��A@ �I<%�s���ˉ��ҁ��]�b��v��2�-a�������a��R,�,��b�OԱ�g���m����Tb,���a6MP��k��e��_t��ܶ�|�*��mfaҽY�m�{e�yN���
��9��u��Ƿ���q$������o��͈r�EG���q�:�>v��%��C���{��<�u�] ��8[�\O9���1��Sp�&b�g��:T�����]g}2QI�-��T��X�aG�v���� ɿ��b�ϐN���=�a��S)H��'ȫ#��A�w3AMT�g	��+������U��J6�AQ�?�'!�ᛴ�!�0x}�E5}}����v��.5����&D9�ՏjR�#h)+GƐ��:#���_���J�֊�So�������Ec���z��۽_������ר�<Ә�]��$�UR���-o.<e�����xJ�_�@���m1�e�
�x�lBt'#��ܐP�X������a��"sjV�Ι�q�7�Z��b%�z�@d��*�e�u��-��ݥ�%�GU�-��ݳֵ�&�7}����ۚ!�=� OP�L�6�6K��F7�?uZ���"�I�PB��eqFw
����~�g��<D&��*�Ɛ�5U�}zU��r�����*l]��{��2��.���`(�QL$-�͓��gqD��iw�A���^�`*��mI��猤`�Ώ��\5��V�sG+�>y�տ*U6���F�J'׆G*�5�{�S�6��E홾} ��
��Uk��I�AA��ccY�X6mA�0 Z!/��s�rw��YY#�k��h��W���~�4-�� ���"��^�S�σ+jy�cT �Ś�J�ڒv�R@CtD'!�~���;����ʉ���Зb�[OZ1^K���@��/��_�/_�ƞ?�@#��<�&6�>���&�]�;�����4������4���J2�N���氃����ÄoYϦ',�	kE����TD���FCe��5ݙ�(����f�=^�����W���ehu���*𝄘S�o4��n�ɦ�3�9I�^y�zS�B��ۀGX�%�]���tc����Q�ߓ��=�V��u��W�ߝ���.�ʻ��=?�Z���U��M�"w`^�0\GT8���'��P��ĲÔ����Rı����_��熮���L�ȡ�跡�r��Y�/E����_�?}bm�-��e�û%��8�)4�����P��E�ynR���K�n���*=qY��5�m�s��)��]$�Ԡ\OM��C��Bf�eE���< Z����`�E�`cxO��)�~�I��t	�3/{%��Yn��Q��qsb�$F�h����1EτO���ki�Aa���^x�&g�����=9����2^�nA�Q6�v;�a�s��`�GM��)����S� T1K�])V�PK�~�fb(�F�+	�#���Ly_�:�A#>��r�P��?�BL��M^5gb���(
�4F���]���g=K�$��g5�}`��R��+q�	0����f#P���;Y"�ףd�'���,7���`�t�J1�(�}z)>�u� �8�p�8�	C�c�"͍�`���#��{��/g��0"�)o_#]2���]�7�ҡ���O�p�C�H"�W���O���L�*�� ����^V�M��B�D��g��,�k����"*�ŋS��N�0_]
>�p=�l3��ܜz��W���]i����b����/0؁��7����W\�(�z�8ǜ#3%�B!�X��?&m|���Τ��}�ћN"����5[*�H�~�D�v���]���������t�~��:��Ni�\o� ��(O�F�4eA�e(e��=��ϥ`ut���� jG�Q�UM�s�肫dT��� ,���!�h7Ai��a%,f��\�V��%k��A��?ߵ
×�^y�ɯ�~�X	6w0=��؎�M����[�B�6�~2{-�{�Kܚ�
PM��p���e���c:�2A �9Ͳ�[.�.�ơ�#��h���ko@�Q���C�`S��O������%Ĭ���xClVÅ��F�#/Ѯ[�Pý}���^��2';��5�}��3���#y��Ô�CI�[�Gr"�)u����8VW�'�J��S
�����W���V
.�SL�Tͻ��#�3n�ݕ�g��n���f|�J��QUA�4Y��+����%�����'��g��a�'��ȹ���a���I�@]#^��3|�wh�*�^�UU3�������)',�Fmg���<�|�t��x��v@������Fs�
�hr~�|���?!�\��-1�f��l)���sU�׷�5LO|�w�@O'�̢�:3�)���,k��W|��`�E�*UXؐ�T ϸ�ѷ���]8��k~�	�Ŏ(yLJW��y��A��7�ڱ��DI&G��#�-mj}�A���'z�Ѷ��e�� �ʲ���eqɷ0| �,3=�˟�y�Dfq�9i��
fN�!"8gXQWJ�����5�x�bqR����x��Bv�C�]��B�RD����.0=$[Ee��g.�u(��F�;s�țQ��Id��k��y>| �� 3�)�ǅLC�6�a�G���p� �_1%���v�5s��דI�*��kf�F��*!3�+�ks�͚x��۔��tS7K��)Z�i!DV�C��"�#Q��lh��WE1�9�����rHb�7���?���Q��r8o�O+>�h��;��S�YCY�ǥ;�9���E��?�#�='����+��e&\�����
�l�&G�w��/�$MOfk�9� JKUq�m�G8�B�{�Y�g�q�1�,\������T*GK�}�_�[e3��3���b���C����ON��5!#�k~�B�0O2)�!����x�|`�������
6E�����_H.�; ��*��s�ջ���<1hU��h'��d1�h�$�f�Xg˩�r�B�A��+RZ���f�K'ѢJߚV����}T����M����J�ѕ2SJ7?e������u_Γ#�#�:�-N?�@�1�<���N-)���؁4#�=bvٲD2%1�a�^��w�2��șm[,���*/ߗF���qwm��>�b�t+��4�M�ۜk� £@t<�Dײ��0|��T�a*�[Y�{@~N7OD
>Y�9ƉU�&n�����q2�ch|���,�o���#1EB��DCV:ɴ�vqa%��tC���{N�����L�55�[��&9�'�1+ulSK�t&����^�,ī���g8E�I����Ϡ�X���G��<���Z���S&�m�N2G��B6�<��SdK�c�Ȧ��Ĝ9�3�u���	C^�+^���
'���+�E�����?҆!���?��0Sۥ�NF}ʙ�qg�j4�7�&_O��
Dv��p�+����槠��y�֨F���TF�bBKy:-ր��������_c#�t�Y�����B�Ƽ��M^ZU��/��do��r����!ƭ�\o�ɣ��v�eb��x���t�����]�-�����ۛ�ծ�r]j����F72���ѕT�d7�<�@��#k�-7{ѥ�;;G�_��^}��U ����ڜ�Շr=K.=P� �L7���{���h��[���~���`�B2��qA#�	7O��qp��W�<�PظË٧��X{}u� ��r��	��>]��{w����/<#�(��y$�+��S��q_�+i�����^��{x�I�����Pc����wdzO���N���L�prU1���J��\�bD�5z��SZ�c�I��4n! �=$��k�#�IG�A2�<c4SF6�����:�!�!����wK��YtD�抛h�
W�oj�B-�2��T="���^�.Qj\+E�gc�ɒ�5�e�Ֆ�ԭ��C/3�!�D�z4;woFgg�$sK�������O��1y��Ć�2@|H|/�`��%��8����_���46۾�aF8��;��c�>fY��6[�L9��k��e����r��wP��x4����� ��o��^'�.y	���.����F�e��ݔ�\��h�!z\y��a$�2�03q�uOC1�%�.����*eu�"���!�\�q���fz�/��l	G������܌t�x��ɷ��ι�=D���p��WA�$�S,���٭�iN�5���MMh�i`Y�y\�Z�˴�V��Y������o���OC_R_�>����2Dע���L��P�|X��Q@9ԍT��/��ł�GX�Z\Xmy�H�@����l@%���8���4Y�F���py�_����n,�*���Y��C��4L��'���+$Viy�7����9��0�e@�8�Z�c�� cE�$�cSb6�d=��~W�]<�{��kY�onQY�vs=��F��Y?�1@3���F��~|&i	�o��;x�(�gQ�Ŷ)=4O��u��2n\_��SG;nu�s�|d���m�$I��ސ[S���1f�)ї/K�=������	�8�� �_xz�A>u���%�P��?6�ĝ���0G����;
k��F���J�|KXh ���x`���X+,\Q	K�Q�#+F��v|�r��Ꮭ�%��7z��{����,(��_dBu�<�3&Ώk��Įt~���&#�`"�\(��<�� �S�7{9��;���b��T����C�WT�$���񿭌��n� sf��=NMq���?��g���&����2�@�p����k�c]�w]p8u�lc?ۗ4Թ,s�h2��8+ͦ:�Gb�%2���[/�b�Z��Y#\��c�U���+%jR�S��?��ߒ�Ȯο�~}��C�):E��&5��{H�L�DJf�Y��)� D��7?~(:�:U�Yi��r�Y[��� �a.�4}s�@�ʟg�j��uo2w�jc��l�Uȼ�slz����OH� [�9�_�#Ai.��a�`Ãf �V6��A����Dk��y��Ku���3x�wk���s M��N�F�B|&�~!s-F�K����E�������8a�/nc�<RA;�#9H��[	}!.'&�-�c��_f4o���Q#���t��`.V�O�$���h�%�ң�]֗��gV�-Tp�#
�&[��>�Q��}��.C�;ϱdP����Q3��"���l��>7��X�G-�)��Y�|�a81ȗ'�u��f���A����z.�����Y��d?t3��6��怨��r�5�����l�0�0�g���/HӚHq3�"��g��go�ݔ�S<f���6]��n�.dwÕ��Wmp]�7���Flgy/mR��7�w|D%b�֋ɑU��oa��!;��E�7r�#�`�?|y���ف��l����N�"���`5���r��O�����%�D�ҍ���2�-�,:E�+�XӤVT[b"Ì�S��3T�7��W/�c]�J�,�y���� ��V{��_D�
1�i�I�h\_�ԅ���'IuMzU'Ѷ!5�e�x�����_30wu,zG���?�y��tq�J���f��K"��Q��
�a"�D���|8���8���R��P[w]����R�X���=�%`[ ��Ђ�����#���ls�	�Q0�2I��k�m�>�&��� �)A���a(��P)p�vJ_lV~����5ng��4�*��f�t'F3�L�k�:7�5<����t��iK���)u�!��.C]�z�j�Ҭ��j��gW`W ��9�	��SK	H��)7��I�ډ���ͤkG�>�WF�]�.�KC���ֽ;�����׏#��o����[@�S�*d�����!��w���/j2�j+���� %����'m+"��=�������,4f��#�N����w��ɧ}��V^D�EL���ݕ�A�і�}�*��p�g��T�=��O�l��WA���|��z�gi��-��E�0_���_����9U����!L�[Z�w��U0�	h"�d�a�ߛ��s�4�����r��՜Z��.�a��',g��U�����T+��в�J��ƈ�L+�-C�7�T1���0��,Fu������u�q-�%@��<ۮ�	�ʉ؟������2�v~H2�cOa�� ��!Ƿ׵噈,�����|�����M_m�R{�T_b���(�MF2^k�&��{U�������2�m�;[aEn!Y���{O5Nr;�
��29�pqׁ4)�a�qM�G�h�`��o7�M;�E=a��4�:�ьv(%%���C\�K{��r ��7�Q�[u�9���1���S&�i&إq�����3�87g�wI"��JnaX�Z�G��6�7��Ͽ��)n+0NM�,��N��\S�n1�C��ȡ�����:3��z7A\	��+9�p�EUZ�"!��@N���8?�Z�!�Wp��^P0.YS���}�*��l۝�����_�&z��Յ=��ٙ+�.E��d���Ϝf�����ue�݆NT�ֻᏒS<�����_�lS/^������2���;�����UAu�wo���Y�U���U7*ˤ���ێe��x��9t�Ab�R���H�	�߃�vky�9�{j�m��'�7�ϐ���Ѱ!d�`��~�^�6-�]���q�GUk�[�����-�(�w���=�{#P�hL\W_��K/��l��5b*��T�����B�L�q<�Sd�[Ǌ(���D<:������<��k|G}pcq:}re-ܮ0�X]�]{Rٜ�F]rױ7(��$��X�rWqz_�im����a$^M��r1I��D�Bf�Dd���a�.m�)+
"�4�iQU,��pOJw��}~�5�V�S5����a��=} � ��q:1kx�=IlyA�I�c+�6���fu�!+��)8�w�LY�#Y�a�Rh���WN4���G-��yϯ�$"�t�^�)��l@+ ��cʲ�з��к��8C�A_!�*���0;RH��[dʿ���ϩ�kmO�'U1��s���@W�
/`I�e����������&6/���܅���;���ٷv���"��]qd���3O�D�o�Q��&�� v���BoN7'�i[	�IB���`�~hg]e�ݏ�LEn\��?��^���9O�!�n��u��K� ���NC�嵳�=�ɜ?r���3��ńz����Gy��{��/�tY/�=�	��=�k�k]W��K���� ��� ���6��dNM��`T��\����o�I����<S�J�4����R���k�t�]`?���L�W�������0�O��/�f�HO5�u[�m�҆����1ڀ%$�8�Y�4��&������yd�v����nH��*sP?Y�g�#e�GE@����$���?>�-*��x�e;�Wb�Z�f���E��c.�⛟�o�L���f+sd�{��`Y�
Q�ȇs��F{!��G1;-�:�W�9;�i$N���Exձ�gK���QJ�=/�F��_�2�b?nw�",�c;I�ls,<�}Z;��{�9:�S=��1�}0)L�zK�Eܶ��|�k	�mǧY�>_3�SAY�H�h`7P��?q�Q�2+Gl�G�n
&�FR��S�Bl�K�8P�����s�ļ�V+��	f�8�`�#&P���)�	_�3%�PU75�9���@H(ss���Hu���.�'����:����̓i��E�#R]��@���h~�ߥB�j|�Ri��S�:��CΏ�/����>��W��?s�چ� kz N���D�M�T�:F gM�������5������������]]@�xp3hl�k_�R�1�G"����W�ʦu��bG���;�/�fb�P���'�\aJ�0���T'%���NF?�Q��K���ڂ}�恛rH�<�5�?,H�:�D����D}j�{����~cx�:�\i���%26�j�6�|��4����$��X���giuj��sz^j����,TUCƾsG:!��܂�#X �1�^��
iI0a�l�A}VY���c<A���k�󗌤�y��O�%!�=w����ҪM�m?�˦B76U~< �-�0<K��K���J�����c�וAVy�9��c[�a].W���Y��^i淺@=o��Q>����$W`	�2O��t�[�%�ZǸ��[�V�����#�&[.].���s���̉s�;��ZkJBs��3���]F��5�9�w���G��)�8:��VV8Y'Z��8����:0�gD��Bڮ.�E��J��?{�3�<c�$�D��2�����l�����*(�B��j
u��z��gp�g"ד g��Tj����]Y'��)lw����I���ɵ���Ӣ���QLm�1P�2n+|�W��UT�ɬ���9���"a���Zr���	��?�j��c�ٜ��l�&�)[��-�d5����mD�O�}עnB��_��"(w����g3�EL�X���T�,�GՓ��)����׻�@I��aFJ��	y��%F�iϭ �!�YD?g�D@��k(�����[�'�~�z\��<Xe�1=��m�5zI�l�0r
,�{��A�Ay�q�N����;f�$�"n��Q��f！ϧ�����g�N�g�%�!�����]J��r7�R�.j�!)�=Vq[��%���7+����!OsCjQK^�IZ��k]X�>�l��V.�)��;�xY��aCeh��Jp��_���,H�5i�,�I@;*lRxf�y�-�3~�k������"��*��KM��)�#!:��C8��(���G:�	�ş¸ W�*R9�-���H�o�75q��uC��o�(1�&_�>g��1Pz	NCϜH�q�ո�9g�a�E#_c��z��!0|�{�e�̪@�a�-zwQ|I/%`����*�  ���wm���8���u���� ����U.㛺��g}�QwQ���w�x!M�1�z���
*ƫS@�A�A�8}dO��}�&r�1�0|VT�B\�hS�Elu��I]_�*����Z�-��i��6Os�U�1�ht�d��Ӛ�챎?�	���������ZJ�F�\'�K�T��PT�	6Ѝa������(S�7�ct������uj���W6˰�;-��*@��]<6�������<�	���!�vOi�2[��a�� �-�����f��D�,�ᶨ�D�������>m��R��$b]���&;_M��+k�l*��V�E�v�
'�������a`lYR7{�?�N�G�
t`�9�w�������qhs^u��;D�or�k�YpE83���E�:?
vC�B%y*�C7%�{�%�����Y�덋[0T�9Յ�1!��S�n&��X��sV����g�ʼI5����[�X��`G0�d��%��9l�	m)	�NhQ��8�M��Sڱŵޘ�Ȝ�}�R�,3r'�R��	9EE+�g���/��6�;g�R��?HN�!
�f�5-0	�����}S���goJ� �(&��!� WB��+��-���Y��]b��2���0�ֶ��X�/���PJ�����_����������|ڴ��25U�6e�lFo?������/ƭ�1q�!a~e�0�x�Lt8 �1��c���$��Q`M�ts�j'��۲�7蹹�P+��d-����9{ϙ��-m`A��ǧGfj��<��˅��-�RPm�K�Q=��P�"L����g�g��/䑰���|J����mBh%q7�"���E�?����<���y�ڧwe�K}k��;r �r�K��]�h{-%
��$�r`'(�w�$>���^�q���i�q��X!^�w!��GI�
�	i���ā�"�E�ʐ�]v0ݦ��U'� ��,�J2�Ԇ��e5p�S.N��IN�j-� ����|�k3�I:��A(2Rc�"6�+�Г!�򿄥�w��Y�SV����h�0�WKLr�O�E-�0�
N�"L�^�D�`�0+��c��k�����5�c��C�pq!�0)p��;-A8�o�Z���z��sY�O��1����|��@2pi/A|� ��̒�Qf�m�6Js��W��;�;S��t)��`f��)�B���)񿧣xK��að��R�����oj�/']�a	���$|h�#o?�8e�:�݊����җ%f��!�WzF��p����u��>��䄩p�&V�X����s���f�z$��z�Giiv�6�}�Т�t�?���D\�=z�m�f�YW����B�v|�_B��9���M���`OZ�\X���*� �̡�w��%�D���R�m�)6p����]��K�L��U�2G�R6�C��J��/V!�w��z�mo�P��.��lg�%� �8�!Q4vl��@���ry��웈�n�<*�qY����~�������!$Lz(���.�h���&�e6BS�45ZEհ���E���c	����B��IXϏ6ά�{VO�Y��QO��s�FI4D���16��ϕ̇��i?��zx�Z�g��4��U=*�B�+�2��&n������;$��sP���a�=X�WS�~1�	6)ǖ1Kf��v��?	����ɡ_�YAtC:��WP{:F?���͓�&g۷���
���F����@�GYK�(��Q��n��c�+�g	�3GQ�#�%���+��k�����y7��������(N{���u����)}�!���:�c�������q�#Tc,��y2�ʴV�:q$T���mw�ξ��cDP���-�A6�9�W
���4���䄛�I )�q�l�M��a�5(�g��-��8��Po|�6b�äTe��BJ]�Jp.�jl���ē�b�^w���צ���b��C����/Aނ� �B��\�^��R��M�o%���I_�?7�f����'b}v/���ɛ�w_O5,��H�H)D I��g^�_������-~�֥:��Wi��6�*��%���4s�����E������ueE�Νmjx`�����U���s"�x�Q��� ��]��$�idc�a�)b�!V�<��A����\�GIy��k��鵨w�{�թ��M�r��lo�B�e~WG�-;IKmH����}��R����,���ck��Aq�99>S�[�f�.�G���\+Y|�;�oq��QY� �j��`��O7[���m$%�~���t,�V��f��#��g[i��N,N�������;EI���'F3jф��µl�4�ԏl/�G�vz)��B�r�v8�	I'�OO������[���4��K�.�����j��N3d��C`���=��z�'��G�?x��ޥ�
�~�_�=9gˋ��^v;滔������]��]�$�OwyĻʏ\	�,�-O��}���I�m81��-a�|��������`�e2���*����rO����0?2���HIٷ��l��?�6�h��5p�h�iO8&�)���z�l�����5.�L/E���X�,�T���x��?�-�ƻ�I�مQJ(dyy����r�h��<ÛD�3����ޚ�N���E�'��3z˰}�W�*e�m�[o��p�SB�C0m��,0�e���y)j*q���e�lf�i�"	�`Q�v_�ا�}�����-�B�ć\�9���]�����!Ru$3�<֎=��N[�$��F�����{W��s���Qf�I��k8c�>-���[})��ǖ�S�a^���vpm�M_�����5dSפkR*'�tf)1	_3Y�)k$��k#^�̙�܅��K�)�|I!�k�C��cY�����=�:�Wv��9�q��I�zH�&�7pӕ������w�H>�R�b��c`C
:��'��ⴼe#&m������H���&��K����w�~B/���ܤ��3 �F�+3ma7"�3}��jόڢ���k�DI��v��%�}���L�Z��ܧ�3���L�"ь���5������G�3�(OCS�RG�Lk�|�������'�E��ý�w_Y�Ӳl$�ޜ����\��n-Uf�Th�dB���U����?���u�Ӧ��4�Z��։Wy�'�Os�˥��T!t�h��I��f��#��7P�׊>��,�vu�:�����9-��@���<�Cl��ى:����<��1Qv�tL2�(�a�P����M�K���D,y-�����������m�T&O�jbH��An�M<?k_�6��wK�!4�f��b1���Ba{�%Y�3{�P�N�s�
�9��]�7!��ס9q���١�� Yo�^��,�E3%	�Uw�:�jkv^��%���C��{�g�ݨ���F�c[�;�9�d1�\>Sܛ�&N ��/MG����%_gi=~IP���@i�Xy�kGkLǥm�:ǌſd����N����߽́S��yc�ȗ�ĭq~3-�1ma�	��W+����y�Xl��6 Ň���?b�!%Ne���0�^1Z}�K��b#�{;��ճ�&�Q��{���K�+3ʍR�����0��Cw����|��o9
��1�ؒ�	���CR_t_$����H��(Q�W����̐Uw4���o�M���	���f�KLD�Z�WY�e3}<x�,�t�����^�~ ȹ���,uQ��#Uj¼��]�7C�"�N�����d��<������<�-����=�G��)�Ѡ2�!�}�#��-�}ۆzo=w�P�c�L�?�"$�.�+�*�W`��5t�B�q2�yT� ���aV<0���Tn㧲A6�#�}f����r�ͮfOf]E{�G��t/o(�*$�od��k�q��Nic�Y��o^�i�L��I�ws��l��.)�ȱ���ߎ)�s@�A��U"4%�&dEJ��Ɔ�R�5�S���Q��=] ����'�k�̮IUA�:�c�:�6Y���JW!�%��2dw|�$Yţ;�W%�hr� W�j$��f;-���e�"܅^�8ۉ-+�phc@��9G��bԾ�fC`�'!W��;ZZ��z��E��ut��gOF��1�������@4�/|����9���f��H��(g�6eo���d�ɪD;�]����%&�]�������:rcSeK���VO'��B�o�LH'?�	�͍�����zHeT��݅Fa���R+Qʸm���	�����R�u [	��	��9�[�\�sN}ɒva��	�J�z��ƩuߋG�y������5�tO�q�Z���ݢ=9��a��WRz�����6���ڃ��ƪ}�A]mM9��`J�\�-q���{�85���5$� �$� ��R0�9�{\ˆu�ӹ`���L���G���ޕR�E��/��N�������jm����Ѡç>%ZUz8�	�4j]ңw�.�yZH�c�qn��*��\Y�����W���r�-�H$�22�Ȯo���J�P&e1�*r�Z �_�(�NE�c�Z��1������=)�{��Y��YQ�E�sΪF��*�S11������/iZڋ��.�x�#Yg��bŇ@=%�z߆�E2JV�n�B"��;�p?s��gճ�������S��'1���)B�TKA:gR�#ڲ�	�7���_���A�ڳ�^5PV�?痧�h@$!���65
��F:6��I8"{�K	9L��M�i�¼�|+]h	�t��a�#�E$�'��C�ဿ�6[�7��<�6��()��uQ���$�Ώ|y�������y���L�#����-���� K��\��Vሥ��I���>e>�����ٹ4>�We�O�������d j��J�fMB���0*�g��W���ks����P�����+]v�p)|�lt$�Ȼ��}ັ�IQ��0���ROb}�0��K0/�u��Ƃl�]�v\�{���ǈ�%;A��D��?���������}�b��A?Ӳ�a5��H�v�D[lK�� ��z��q��\@�~�T):&Ki����Bl���.����4�P�џ[�΢��;��u`	b)�j3���GU99s���P� ;� 	��J̚�T^�iԎa����+�Vϳ�P�A�t��!���uyz���t�Ąw&z�D�HM�����3�B���~r��-�e�KH¸��d倯������@܈c&m�A��@9�Ȓ[��e.���$dT�ͷpUo,]4Qt�9��D`�e�Or&>�U��%�[�nF5/�V/�ᴯ#��/[��i��� ��?4�; ����i~�3E������P&��/�M��ʖG^}�)��s��y�8��)'�;J�na������x��c.����@����Rt3Z9�Z"Ԩ�v-�Fl���%�eo� w������)��Lg&�m�]V�w��8=�{��5�/]�p���!w���J����6����X]\b"m�P�(t�|U��˯5��Tu��JZ�R����r�*���Q?���ِ��W�l[E����ף�5�es�cvO�����ޕ)ƍep�ó�݅ET�XĠ�Tl�ýr �v�����ur���J�/!y�0,��;�#���W�%D5x�������6�؝��O�'Z�vz�%*�r�ee�0
�6�ٻ�Rݏ0h��,�D����yDa�qx�7�@��f:�B"�ٓQ���r� �uO��©](��W���C��!b�] ��(��R0:@�W�>=�[������S�m�?����s��%Q��`IPذk�E>hY����N)������%�ay����pH��_��b��5_���	*�fD�����34o�k_���G��0���l�K��)���!0�C�b� ��}7f�/�x��W1�W9���ġUH{� 7����F�EC�ީ%��>9��'�&��CE����Ҹ�	��]#�"�����\��\��v7���w�{/�*�:��� �A��m�q �.i���]�\6��ſ\F�Q��3J}P6�G	`�VUX��H�g���yg�E��!��w�e�.�O���$��gQ>|L��������EUCJ���_���'���:�ݝ_�x��6�(nU�~h�/d�����ė���Nˮե�o�5Z�E߉R��'=t�߆U���CT����C�e���	�"ȕ�7��Z��@��G�u�`��A	�&�k-�_@��<�
�:�G�)�����2��avşL2���a~6���ķH�����,��������26����m���e0b�#�\�MM���k:Xӣ,�x{�	��C^�l/Ta��cY5{��wN#�<
���9��-גGt���7q���T�����o�b$͏k:E.7��Ȃ:��vy�%o9JC�{:ʷ�C�*�nW�f<[�C�9d 1?GS�ͨ&�����a��q�I�/g$�cIk�Wܻ�XT��G��]����ڿ����$N����.X��	�SP��N�Ȓv�o03�X#�!	/�V+�ݥ���6����1	�ۉ?���!@�k�+*�0���l�3}�<�]���֎p�rW&��<����j�%+n����렆{;�w�2���s�N!�I��l�;�$���}�_�]`|8�����@�2xl�9��U{��o�!�i�����Ɔ��5��˙e��Lx�,�t�ߛ�����b#�v�������j]���(�7����	��I�d#r��d��-����ӄG�������<������F���`=�$�P��`Lmxp�ݎd�.���5��2�݆peeB�6	q-u$Aǻ���O<�VZ�/O���=<��}a��K��r��뮁(Y]~Ac{�U��3�(���$�p��?��q�K*i���e��^�{5��I�E�SBo�u摁�`H;�)��pQӐd��V�U������J�4݆��z5f��S�'��5zX�l� �	���a\k���Ip�
Ac�c�r6����7��!��4�:�Pw7A�Y�	�Ҙ hM�
W��J��l)-�V����5"¿�^#ەVH6+���c{.�š��������C.�!�Qf��;�,2��ʐ!
�p\3�)�(O�u1� ��r&;@��/�_�6�����������U6��
�MA�9�;�ǌ��l���
b����������w�\�.��׍}��k&����o ��'���	򿯜�|�����e�)�݀��V���Q�啁�M[�۞pN�Vu�M���_�c�h�ю>�B;�/��(�zZ\��p�G�,��G����t���5��ߺ~=���\�UW�h��?���Q��U�B��;)�|	�M��e`E��\��ˠ>��S���m�~���Ԗ;`ERˊ����&8F׎�G�#�L�����v�Ț:y��@�E/�|�y&���me:���2:���%�ɐ8�4�dX�2J� xy��ݛ><n��.*D��Y����4>0�x^r�H�7$B��� ��s��I��e,^�s�#Z��r�C��E}��c�퇛P����9�AA��`{�VYY��QE�s���F�F��1,C��KT��j7ziu�:�	�ixf�g��D�"�b= ����92 Bn�#y���;�as����N޴��%�J��Sn�1ҁy)��Ky�����MzP	��D�jh_d��A������<P1��?"�p���X��
Wj�FUش���4�\KDi��=��d�[��+��	��=��#����bA,�ސ��{���7f|�謱Z�(�VP]u�k�j��Y#Ⱍc�v���\��'�W#�内�Jݘ��[��g��n������
����@rF�w��/�lW��p��+�\�� � �UG�M���+LAg^}�2I���f�,��Zbz�W]��p$i�lϰhۃ�c���g�T<�Ӥr!�&�$b����Z/�,$�%��x��\y�����Ì�%�з�?E�?��|���+�e}l ���2��e�5b�NH���D�y��E�A����왎�7��~� :�x6i���6{ǿ�;��Z�4i������	L��x�u[�T�Dlj��ɦؾ�U��ysؤ7���f�v� W��Zً��i�e�a�r1��o�V
s�r�aA{��|i͗��y*��a�@��sPwW�C�ߦKM���"�Bh%�~���-�K#\��1:��,���h���vc�g9A��94^,[u�1.�@�*UO�۷ˏ�o��$Q��:�`fm`�UO�!����%����ɫ��-?VJ\��#v�h[�ߵ������1̚�X;�`V�#���j3 =C���Nt�*5�"��G�~)��̼h;<8�˺'H��	�����d�x�|�s��.�mݻ����i3�"�� ���Hy��}��:���9��� �M����Wl�W�g���S�GqD��x���m�p+^]*E��D�w/s��5�E�#
��3�aS��mn�Ȁ#��|���농����Q�[��㍚s�1��r��1���N?�B����M��׆l��6��	��S)5S{ݭ^?�O��(���ް�'��3���Qo�ߓE�m�X�4�T��	�x�,�*�T�#�(�P���O.�J^y�	W9��޽��r%�D����Օ�TY|�/���y�'�Z�zA����%	e������DxQO0c�,��֛r��y_x q��I�H�fuT�"?_Q��$��_I�0������m��K�������d]��>����R�o��r��=��m[�D���/o���=~=stL�Q���I˳�k��>�� �')� �LN��qa�NV�*�p#��_X[���q=5Z&�Z"a*�vZf_m�"�3�k�k�͡����j�;�K~s�)᎜!��hC����0��@��B�Ӝ"W쐰91Z<�?��HV�(7�,�F0G��g�9��Wf>TT��N���C�Ԡ�B5�~!��rt'#��.)������f�Ev�6�v�wb��/V������� ��|�m����)�
� ����!Q�S�:���,C�n}���B�a�������ق�т�"���\C���)�O��+�R��W|�P�ӌ"�0YE����__����`�U�f�ڳ��ڟ�c��U�� h��d�>�����s�zI�ˉ$����PZ�_�M�;'��9�A%��7y�T����9���\Q���C�7R������b5Hu��3�j�:�a�-Ue�@�<GX��i��DT��z6����v �2,n�ay<H�>wٷøB��|,o$X�q�S�m����Ům���Vvb��w4�M2��k���g:��~��yu�'�	a�&�Y�VI{���N^,}
E�9�L:���M��q����Z|����o#ھ�*�#E)i��:>:p��v�5"%��MCȹ�{uL��ކ��k��[ak�9&�q1�A�S��&�w�e�Q�ki��� g߂mI����6�]X/�G�\(����������Zb�N�У������S�;{��X\ȍw��c�B3�!y�'	��A+�0��1Nh��7i�,2u�c#�?y�![�z��X�0������}$��X���1��KQe&��qc��E}5+��� ���:��ҭ��p��':����T��i֧^r��V��x7E_*�uqj�7@2�POw0�ta$U�;:��
�oP��E�n�5C�A����ϰ�eiv�x}LytI���>����&��9����%��j��ҙ�	7�8��ı����d�b����Q�Jr->(>���=Gwjh�G�J�W.��ţ�����f=R�mP�EL�!��:)�I9ڑ!�[��L��v�B9o�q(_8����vCƩ	^<&(�
P�(Z��J�}\���&rQtή�!�]�]�{��2�2:�C,(���$O�����q�/niY�n�@��^9����ZI���箎r�0����/P�8+��r�Μ�w;�U��2�Jc���5�S���p�+�;� �L����kd�0I�@�A��mc{ʜ6�"�ҟf!������w�Y����M,hh(�dW�� �-�/<��;"}Ë^>V��&K+��9c����<:Vؼ���t;Cּ�!8"�Ü;��mla�+��k�.���O��1 R����@�f/����k�#�b ����6��������;R��E>����/SP�����0g�	���#��������Wo{��'��M	�y���fң�'e����{\f����Ȗ� �]�����y Z�uV`'�t脺���8�ѩ��Ɉ-�[����ކz��Y�k!zGz�G�g���!�/tEI���|��?�=K��W��W�(��m�lP_��f.�|���\Mo8q`@Om\iZ�[���ng��%ö7U�v7�RfI��~��	��I��>��L��������}[�T�;E(/g���4�Ҿ�m������t��K%�^?8|9 4 ������;��yP�X���n4�
*ߎZY�s����I�3���c.�$���~��w����e'n�L�Zv��^E�5�c��������j���@�EQ{�
_Y�Q�BEs�FgF�%`B�1'��Ϧ'�%vii�����#xA�g7��Ž8�=���<��2��un�$&��;��Rs)���������S)�1�m�)8��K��I��Y����	ˁ��f�_�rA�h?�T�P�)?]N�����ѷ�|
��Fp�E�?����%K��"���_B��t��+���	Ү���b#r�8���*�ySu�v���'7!�^M��,��(��l���u��/�Kf�2Z��k�����oCz�]L#W�c�֘�X��K�����a��?�R��+�{�`��u�*W=�+:�F+�� �aj����Mx���&�g���������w��XX�5�����]�w�pv[l*]��>ҹ����N{��^�amb�<ӑ��/R��<�ɓ��\��؜y��4�%q�1�:�?H���7��F�}��s�p�v�(�5��_H�22D�o� �I��}�g���Z~O��:\�i��>�Ӣ�V�7��5�4�� ���7�D�qi�uV�c��[j�̩���U/,s�]���m�V�� �%\ 	؋�1�i�aG����VER}�Av����B֗x��yE�q��x�z��w���z��MzA��}�B#�v~�|D-�K�f�l/c��B�z�p���c��AG9�r[P5..C�����J���&��o��YQ�H��fb`ue�O�X��e�%�p��$1��^/VeV�+B#QR[�u�e���P��tI;v]�V�_�3��zI���%���}a�G���)�M���8x��'Ft\���t��D�ӝ@�.a).*�L�6�����/3�Y_��?Ĩ�:!���?X���-��F��y�VS��O�&�	�g�@t�6�#���@�K��x�]�99�̚w��m��T�D���������m	�`��S|a��A���������h�lX/r ����'?C ��O���x0l������5�?�Y(pOI��Zџ����"��yh�SX�E��X��T"#��3���EB9��䛻+$�����J�&y�#��ϙ����D+a8���;����܅�ë'�z�n/��qe�����K�!#+3	0^�,A���->fyz��qn����`f��K"�R�Q���(?���}4��=S�Ϙ�`�����W��]�5}�ޠ�R��&����=X�[g$30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��*I�HO�@kQ����^|�e\J4��\2A���;٤����U��'qH��N�,}�(0��qp�2aΖ���I��6 �*�J��#�_���q�W��83CS{`�!��K�$sL!��c��X���/g�BX��w�u�tKN?����K=\J�\%�	�fؠ�X�2�}���I�ɲ�dۓ�YP%���K�_�$)!�)"���������/�1'�g��c���-r,���1���Q�ϐ@�&ٍJК+����L���מ��}��if35zǂ8�������R��*����Yvf�	mKǡx���6�o��aJt��� 8��),�/�Q����x�Z+���E�$�R܉��0;iw�H�l��&5R�S�_���^��g� i�d��t���,�����tm2���ܣg��Jl:Ρ�㻡��OA�f��t?o%1���`�K��.ԩ/��Aj���Ո²i�j���ޮ�κ�����i��A'(ǈ�Ɏ���G�����m�O$,K#$��~6Mm](�6M�� ��i�xu߂�J�ci�5��B!���A��F��b��v�8P3�]���G��1�":03�R��|�-�����sW4��!g'r`��,�%�j%��6>}�bn!ˏM��6�����r�O���G�{��6��Q�9�d�{6����H7��g�rV����1Cx`����M��2��]��枯ΐ�S��Q(�"�Xh��I��٩���A]L��"�^1/�`#.gH7�{��qI����O$���ʑ��@D��5egx�7m�K<�ÉZ���Z����*f�D��j�iS���g�Ûڞu:���<VJP����bsR�Ǯ�Z���i��B�tHH�p+��ſ��g��s9qp�Đ=މo�������������^7��}IL�MKRm&�3�P��Y�-��/㗢H�[1n�	�
  AcR=������d���l��(C�C���ւ�:���0�b3yc�u:��:�u<�Q.(D>TT�B���A�g��Lyj&��PpK��@�9�ST��T�J^S먷�"�K7�<`m���uS��kL������ه���G6b��]_Wʈv\�?����<1s�����dS��	��~�#�����5'�I1��
v�Rc�ؓ��ń����=q�6hģ�IСtI�A����� �}1�X�U:p]c�=5�h��\&s��&=��Z	"�r� SCJ:��	������׺b�4�/�W@��vr�t�S��*��#��g�@�;�<�����n-���Pk
ę~Z����2qG��^��}=#e�&�/�m���7�x�-N�kE:�XWSs�h�t��)&*ːr��8b�W\x|�"��!UKs-4�c,��>߽�}��Mi1��u��@�
�S&W$qк����sORM�����+SYa.'��Ш�f�ڭ�?lD��O����֙4`ӪUI�'���,5�xy6P�k�������v4�6{�;r����Ѷ@�A�-�U��-��F� ��4azR5\<�	��X�g��+�sB���h��Zj��݋���c�:`❉-����5fi�.Sl�����I �z]�Q�rmB	B�#๵�Y!z��D������4��?��nB�m��T凭��XԜ�5�Ÿ�HT�k���9�R �G&i�i�*��z�i�A�س.��G�,l�W�N"i�����j�;���t
C�*/D_��`)�ۂ��:)�'�$�PA��M,�C%-+��.��E/uT^�d��^�� P/8eu��%^AI����	��$��ϗj�����9��9��j�jx��ƪTU��\.�� �[�:�R%����6m�UI�]���vш�!���bQ��t���e��u~�#^��p�v��g"�e�b�c�">@H�=n&�Ւ�^�d�C3V�p�B��Kv.��e�Y�H�V7�0/�p�9�����	���q��	ݨ�"J ^E���f���#��\J�WLWU|�Vf��_ln��ژ�P+	wU�&$`c��ʣ�l^C8�I_��d(O��L���9�:�����l����S�6-{�|�V�S�'�F9�22~W�p��S�j_@�r"�.y�W}ʫS��$V)�%��  ������r���.e57$����1�.߱� �d�E�]���8�F"#zC�][��Y`F���
�L*�J ���O�Hy�z�.��-ck�E�+]���=^��ڂ��RU�̮\��bX�	��iRb
���o�ym .fxT�E�8.��%�W��blJ�U�sR3a�r�{ ف|Z�.{���@��_p/O��C)�|{	�* <�r�̔�w#�U����*ވ]�έ���T�yl�?�6����U�*���'��&��//������_��}GvO6��dƓ_�<�~�]�/�Q4����"���Kd	�����J<����T��)�Ɇ�:���o��	�o�N��c�q��ZJ�@c�شӖ�u{�'�����*� ����6��4h�,�5��8�_�̽��=��y�L'��m[�R��h�J���+ƾ��Ђ?@ʏ�n؎c\�ǴVJ�=B�.W�\`c��ѣu�LD ��*�U�a�����	�(��q�s�2OD[�NE�I&L�6K����U~�_���q��μMC}��K�I�L�V�8^�T�M��/U��X6w����K|�"��l�~B�\�f�%�ckf�@�X��}:C����I	�$�m)��� %�B�9���Ҕg����ќ�������� W
ĕ�c���|O+-������|��Q~n����ٻ���\f� �*�,�ܲ�}���f�cF��<�"R���p� �U*|�|�<�洵x�f�K54�x:���ܳ��a�!³��18�(d�a�Āq����H��{���ˮR/qN�k������~���|R�U	_�0�^<�gO�R�7ɂ_�8H,;}��:t@p�l��g%�l(%����'�.כAI��T��t�J��4��z��L��ָ/Y�A�q����p\v�ؾ�&���!F�h�5��|���3���z�(u  ��k(�ba���m��,��b���6;�
(�ӌM#�����f��d��c� !�ܒl�~K�Ǳ��P��Ϥ��P!���d����Rw�P�'3ɶ��*���h�Dϡ\��Mo!0`{�F�j�������nO�M��q6Hw�1�v�}�y�5��{O�$���,�m��Rz�6�;�F2He?:gt ��<5�1�9����o"e���ϔay6]��۞��]�jm=��w�"���,����g�B]z�"��/IHD.�%C7�~�_:G�o�YOp���<����6D�Q�e��47���<揉�R�B"��@�,`DL&���L��0>���u�#� �y�%�,V8$���b��f�H<�H"(��W�v�L�����^��s�f��*K���p��S=�З�y�����p�r������Ċ�Z&還gR;.3h��Ň�芃-��Pi��b��7�� �R��X�Rd�Jx�x�����ͱb[�0󤛍Q�kgI0P)�y�yG:�?�#�KQ�u�>�OK0+o�cg2+�y����x.K^��ʍ�S�̈T����f-���P�7�A�`� j�S�C��0e��e�d�-��n��`�W�HqN���Q����I����--|�YZ�ǵk�-CX)�6�,�֭f��4�0��k��}�x5�����Y?�I��[����4����k׀��!��C�ޅ�$n*���Z+l��&�$����a2�B�+�Q����nVh�S'��m����=�2rin���T\�@�Ck3����L��H��d�,���4��Z.h�_B�"�����l��,ZH-�g��bfg8o�m�{�"2j�yr4�y�2,|�D���:6o'	)t�B��Z AyI��7
9|"��!u�quFv�|��U?(7�8Is�t���-��6[#E��$�6��i����K��,����0��Q���#V惨�u.��4c�u�E>�B�0�
�U��D��!v�U�u�k	)�O���RH��y%�FnJ�[]nX�eB�����p�K�y;%+%����ӿ������ �)6gAha"�ɔ>r��I^v���:v<QUK��>�"���݃��+����<}3���E'��\>�cO#�>4P�7�oh?����9��ҋǁX�aݙ5J�;�eꊴ�EN�g_B�]��*q�!��=���#����Ae��*�J:7��I6���?�>��'o��8˷WZ�������KL�l�m�`*?
�DUFבY7�����g���,��L��#���m�ߏ5���S�Z�4��[D��,����A6��@4�~�	d3�����0N�D���#�N�Y@��e]rS�e�1�E���{]
E&����Cߠ҃�"�s繅�hٙ�L��-��1��K͐#���k�C��N5��.<!9h�x��a��*q��ߞ�J����g���*e�� N3}��c���jVؓJ�?_H�\m*��u�N?��3,�`��@n���\I�J,�e� H���ql�߅puhW��L�Q͉E-:��l��;i�}��uS�:��7GȚ�F7�&O[��Ч���)hg�eG�㳏��\�]u}�r)O�C�T���-��p[)����D�\��j�����)i�����X��)tǿn���嘙z�B��iY��������y���~�*�S�/��-�y���BU7�I������Ed��Q5&��H���t�j^3�K�K������ͯ_R���
�l6@8�`Oj��fϖ�=|�c�±c�@��;u��ѓ4�k�	��rH&#G�*�R_�?�bSei�V���58�z���E��p����Tc5��Gh+k�nlO�IV���0��O�nWx�i���kXf��h�@��|���E�G�61x e}�2f"
�R5i��U��ܳ�gE��
�KHg��,���Ơ�c��AMd7R����v�d��,0�RM�;�T$���qB$e�����E���,:�т<�8�.d��+��X�����>qr����zJ��MӸ��Ե2��� �k�n��lݷ�� �1@�P�B�y��X�p%��?�(B������x�'ீJ��r돷ѿa:���"�{�r���޳�~҇߬���:-��ו�L'w��v0���eS�dtȇx���I��J7*aU��"��5��29�߻&����p3wO�xua��O�SUH3$&���;b�<�C�,����� �%�SHI̊�T��;t��uRu����L!��W|V+�H��/m�T �d�9f���h�t�_lio�ڎ��������@"�pA�p��&��TR��cS��:�^Hi!���]L�5�AY�*�� ���Na��8�[���+�zmrCV�؇�K��i% �/��J��w(�{����V@O�;N��hqD҇���Э{Q�����](����n��}���Mg˰�c��(�BNn@�|�
L��h�}��TB��O�3N-W��?h�
T�o�.KB0w���d��
�MAmW�@\�U����߾1@�p�(�d`�	p0���d���Ҧ�GSW"J1��vh���􁂙c6���� ���K�>x��n��H�Ȅ��z�~GO�B�0]�B	bu���Gl&���3�=�|��O�	�r�_Sp���53�E������8�S�"@�(r���׀�~��z#N�B�M�n���J�@���[^�0P�P�*��ݣZs|����q��^�z=30&S������MhޚJjkR�y�#(s��t�F`&����g8܁�Wɑ��/�!t�s_k��P4���䓄�R�M6�&����M�R� ��qR[q�t;�b:����M�η���DD'뢨���:1I?��g��$� G,4mQ�U���'���,"jwy��*��A��9�-Uu4�qK����_���2r�ΰ��'m��=F=���AY�R�U�g8��E��bXso]��vÿS"������P�۰�`�S-���bK,��݋�T���:���z���_��B��
#A�q�~a�zX�����y���+�&fwۇlBV�(�!�@T��bw����r&��ka�XE���6 	�nihk*X5ӜvWeAM�.Q3��q���ӃWۧi_�O��;�S�.��CAH�DL�����ۯ�%S'N�-PN
�����CrG�Ƚ�#��\T��S1�^7Z�P<�u�|G�S<�A6��9(D�Q����.�"���ڈ��x�����x�f}��U*���O[߷��%_D��\G����DI:����Q��U�����^�+�!{���4uk�*^�R�����4�S�ҽ�pS>"�~��y'��^1w+C`��p�,����+��tY�4��?�0�����&�#x��PƉ�[��Y��U�Jmc��|��M{r��Aʅ)�=J]��Wb�QVH�_�p��������w��l$-���7_lk���B_F�d��S��9�9�����8l��uf6��)��i.���!"'ܺn9z�q~ę���Ԋ��Dl��Q������ ��-����d -����{:Ei����Ze��~$,���.L�� � �ER�!��+3�zЋ�[�b6�&2.���Y{M���r�*@�Hf��zHf��Z���>m+�Ԋ�J����z6ǟB1̛�Qq�VX����56bwB�|�yu�f�>E��d.�؏���/�o�&�^s_���#�{m��|�*�.��2@��L_ݮ[�İ�)8&�{Vd� )L[ͤ�����_Uq�-�~���jڭ��5]yY�y�����"��U���"��'��&Lq�/�7�t?8�#�kG����g���̢�<�"(]��4/i��4�LG�4��*�M	����a�Q<���>�E�v�ƭ�h�ǥ����	U�N�ͩ�~��Z��U����3V��#H{�D����ǗS�˽��,�����/h�H"5 �1�ؽf�� �.�Y�2���Y!��� dJ'e�+�f��q�+�������֎%�]���[7JoQN�[�\-���>(��YV��p~����Ü��4�gZ�(�{�qkT2��ߤ[I��6��(E���U_%��q� �;{�C	��<��KL�L���びJ/�aMXC����%�K�N ����J\�_�%̂�f39�X�օ}�
9�2� I�(���m��3��%�GVꦜ��W��D(r�W���@�*��X�b�8c!����-�<�KF��lLQ-��ۢو$f��3s���ׅԞ)g+}� fn_������d}�_"��4*)�:��El��S�f?�Kb~3xqi�\f�*X�ae���*~F8��gרĭ�9���Bεť������R|��l��>���㘽�|,�R_�a#^�hgP���?��Vr�+,�T�s�Zt(.��Pgeʏlt��v�[��Agx���t��mL%+�����i@�/���Aer��U}ľ��(s_������x]����d�i�f�(�%�ɩ2��� ��;m2�,��V��
6�	i(ȵ�M��d�5l�S�ǂ�זc3z��
��eǾ����l���2�P�{��&%�$b��36E��7C��������J�!��`L�D���jkB���f�0Bn���M�V�6�N��^�L�J��O{\j*�Q����t�?�6IP�s��H2�}g�娐Iț1^.�=q�����m�����]�� �
��w�?�l�/"_�H�y2˔��]G��"6(}/VU�.��h7�Y�LH����'O�E���h�D��e��@7�V�<�͉��EȬ\v�҅�#DY��鄵��}�*����*�����	{V����.b��f땷�50�e\��c�o���ˠ����ә�MX��t�p�o4=����g�����7l���yZ���=�o�mR�7�3���T3$�����]Ȗv?N��T� �ARx����d�d��c����^�ޟQ�ݤ����݌0}q�y^�B:��0�QQI{>ϻ�
p�sGg_P>ye�3���Kkf@�:�S�5�T�LI@W��C�aK[7&�:`(a0�S��I��4��d/�a-W�qnb�`&	��%�$�Q�x麫����-ҽ�����Ԟ���M�v/�{��cU�^���`�kUD�5�\Q+i���Ỹ1�����/��
��x:��}����Cn�ʤχ~F��A&��r����2Wd�x��r!�n��*ST |�:1�,~�?�iv`����@�!�����'й�\������%�u��$Z{���L�."���v���sZ�V�g�S5f��Uo׻���"����ԥ4ӏ&ӟ^n|�X�g�#otT�t@��g: n�Ii�v
u{]|/a8!"�<��i;����7 gI@�s�LH�:x+��S#���$�%��SH��/K��Pw+>�0�)�я�B#�(ƨ
��u��4�����
>��o0��U>���d0t!cp�dHk6A]��0¿E�>����ר�}X�+9�����eŜH8;���8q����-��냷)�'nh�������rO�[�V���6�Fvcr�U8��>~ �(�ڱU�W�1E�Iy��vV�y��o�r>z��#�ʩP�I�o�VH��W)9t�\���Q��&��h&(e����n�t�o�
�b*�(�����U�x��?�e�O*:�>7���6��4?�h���1�ż�W����)ƣ�7L�\�m0R�?WHDBWB��eS��54�ڙ�3L���ɹ�t'��v�S��_������<^AQ��ȟ�jLm*�=N��<�mF�%q2�2�F��� &��ܘ����x���E&Y����7A�up ĝ�%G����B���gqZ�t;'*�'���$ԟ3��i���ɺ(�YZqӿ�Z-l�Ԟ�G��f��<����#�Z�y�08ž�A�mBT�'���MY�� F�M�%%�,wo�	e�б1��H`S��/�(ז[~�G\,�L��	���? H�?z=h��	��[Gy�5�r�M�lij05��v���h������=YF�V�L�ǟM5�-�~g��}za	@�[�A0��'(�*Ԉ�Ps	��s�7=�!?��N?,!a}��������~+;m���F���C�v�%$��@��5�.�����T:uTf�W	�2��v�..[6`�]�>�t��D�q�����^H$56	 �ԑ՘�������в����|bjZ��|�*�%��@���҈bI��o�}�ne�wN�����*=� =�<�+ۻ��r���vOws�i|�m���P�pC�Q�׌*0�T�`)��uIo���,�K�?��Q�D�x>�#�3Ǣ1�#+�Qj,���箄����,6߃q8�%x�eB�+:Y��*r}4�}<*���GqF0��8RW!]��Dʃ��)c}�P�sX�_�πʃ��XӼ����O�E`.{ �X;������;Cރ+��%r?��\�����1�ěp�3��	Ҧz#p����,�8~�]��aF"p���|�Pu@�j|G�&0�
^	�Z[��#$F��+�MXH��w�! #�Az�t��F8Q9�Ϗ/�2^�m�JY�����auŘ~�2xS�N8��7�H�'m}�C2.��?P�>���G�zT��/��~��_aJ��Q�p�T�Pu�YG��L����'�؀o!ׅp❝�Ts����3��[��>vW�Rd�K�!4f����q-r��Q���W���X��碓�<����������!���[��X����^M�k���b�GW�%���B-2�����?��bz|�C�h������Hﶧ��Z��0��0�æbZ��ǩ��t>��s���a�
���bȴx��$5@��O��J�R3���a��N�D-�L�S�w�0Ӊ+�dΟ��[��N���c3_d��MR�7��G,(�`{G�S]p����cn�`�=�t�V��t�T�==%~��p��ܕ�Xmp��a��'�ݾ��y�9=�]��s(���z����Y�ʥ9�/b˨�^�{��	$�uE�������NiQ��QI�������.I$R��ə)�.��k�T~���+����6��8ÄEB��u�&A��µ~U��c�Đp�"��'��9KhyWz�_q�P\��BlS���6��������/0��-�9jI2����2��=�����_j��Gw��	vϿ�֏ H
�2a���sD9��F=��E���bMb4%������b'CY�9~��M�i�31���Cc�)�A椻IG$��Yƨ枔�+���o�63���4��ȩ���?\�]c���l@!:��+��3��͸�}����D���x�aN\�@���eꀁҒ�w1S+����{j�����7�ߍ`�ޯFZ��Byh������"w��ށCK�)���1`�y�{�����9���x��h�lY��݃��+�����ueX�N�s<��D��;Mg�QI��9�a囉�g��OhN���39mM`�:��f^�x^Ip�5��O �T�h������u�g�N�ܨ>���:L+N�9i������+u q�:�ZG��~Fā�O����tNZ(��g+v��aϳ�t1\�66}\iO�T�闡XF[���9)j�L���\�y����2�g���ԶYAe�t)!;;nI���ҫ�z��K�s�&Mض�h���Ȉ���@X}�$�0��s�WP�U�������r���-�5��n�u��6j�.�Ke�ݝ+�\Г�LԮH ʷ�O�8��vj3vϣ0|yK��w�-�?���:������&�	L(H3Q���GR��N�OwOiK�6V��5E����娑v��K�c"�I��F�k�Gtl��T�*Jg0ƵO�BcxwǡI�k��p�5���OF|��}E�h	���>x`E����
��iV3U�^�ѳ�E�Ǔ
T�n=´0#�a��Ү�7����n�̃���,��M��$h��$os�q�R����8��6�(,'�i�L��e�F��U��2,��ej�;s�>�7���UKJ��+���~Ԃ�b���k�9�s�r�L�;�L���,7Ӧ?HX��H%k� �5ʳ�-7��yr��)�<��r(�ь�":bY�`��(�;rAk����~���"����:�G��LԺ����|H��񴍇A�o�uoaق�UD�{a8�"1���n��9D]K&',}r����YO��raq�����3C���y�;��<Y�"�d���T� ���H6�����;8]��Ba����NL.��3�VxR�H��m(��ڑ��93;���A�l����c[���u���m�,p�͢�H������sSFjY�K�\�_ ��7��)A�>'���ɿ�����%0���}�X��m�t*V5O�&5>�Q0��2��S*�+���u���7V��V;[;(h���QE%���QV*/�9�?(q�5�����w�}��Q�����7Մ�)B{b)�I��
�u뼉i}s8�B棅O
G N��~W?�4�_�
���o����"�8��d���]�WD��\����y֍�z�1��c�u��dM�'	������՞�c��]�/q1, v�0��m�&�I2e_VhT�0��K���]����{��̹:Nh����G]]��oG$�[�&-*���=Q!���qg	Ѐ�r�S}?R�@�Ū`�r��]��n�S����@{�r�3Q׍p��H8#�1��:�s�vO�m���(���P�3���οZ�����-q���^�i=�&�sχ�Hƙ�Ժ���k?��'�s+@{t|��&$i����8�f�W׀��!��ms��O�D�8׋���|M��/i��:���*����q�ʖ��IF���M~m?Kz%	���m'2�Y{�ڧ]�?�o��Ɋ��m�I4Z�VU��<'�,�Vy0�������z�z��4�E�uD�ƌ�!���֎;��[8�DoF�6P�..Ro�8۔�'��/���Xs|�m�f�򿠊�����S ��݁U`��-����o�ﵨM���_w��ʎ:�`zה7�,�B�v#NU�+."z�P`���0�'ַ�S���H�B����.ʰT_6������}���@��}�%�*�3A ��i��Q��|�ܹ
H�@�jj�ާ���שh�0횄��������%KV��j�X��s�����9��cx�ZW�d����<��� �
s����eP&N���F��3�������#ğ����$����N�Ս31�@`��#�>�p5�Ih@ś�Ę Ჩ�`5����u���F�6���:D��1������Ru��:
��G��rF�'<O�E��lR� �g#Xy�j�Դ0\�u}T��O��T�e��PA9���t�7���ad҈�y��h�� �%?���h��9	�ax[����x��`��l��5��Ev.
h�w��a�PYY�&��_,��:�5�3����M�T �1����l%.'�6��[0s<�>�=�[|MH3�a����|�`��F =L�:̮:�����vb�T���a-.)�ѻ���:h�ê����v���[����0=ħ�������q����[XH�����F�ڀ�����E��8Mb�^���
|*��KHM���!b|>Sod4�nX�w�f����{*+��S<a z�� 4�E���B�w�o|�I�|/�ДQL௄�`�)�ڻ�\�����^{�?D�Q�>Y��wy#z�n�$׶+��g,\}l���'�Y���Y@8�h��X��+�9?�5�}G��<�r���Fc��8�|�]�v+��n`)�>s�FS�ʶކ���(��-�ߢ�`���&r�����ֹ>Cɋ�t���E߯�$�e�1�A�p3S$��߄zV8)�>�{�_�~mi]�k@F*$�U���#�l��������
Q튓����BОF�O�+z�&X�w��Y��nAm�8�.L�/���5Ϥ��+m��z�%Q۠��pŋ�2` *�� ���@:ۻ��mP?2a��?�x�>�i�Gƫ��,���_�����4��>TTC�u�
�G	�rL5xƙ:�[�� F!�e���w�T����f��g8��1��e�����!�6vf o5�hu�r��M�������J��|̓
tT����6gBNte��Z�?0ӀB�1M�c*����YX �t��-�-��Y���R�b�׎C&rս`�{�&�J�Ǧ�2��/f0��4bmt��_ti��_���z/��+'��"8�+�4�E�@$�ԉ�DFJ�>�=�*a��tN`��-з���w7҉��D���[��v����cp9�d_�be���
�(�X�G�EpU* ��c�����\�i�t��=(�~��pc�+�����ba��5��k«�F=��Ll�"��K�G����ʸI�/��L�־�{n�$cW`E��s-�+qi1�\��k���-Q$�F�Ɍ�㶁����~,gpߞ���Tf6D)��Bvd��y�̕��~h��c{,�Cou�,���ՔyJ�7˲�`P�vU�^篥u������f� �2j�=OɏŬ2ĝ-���菹j ��wiP'v�1��C ���2t,ɗ��D>������y���v��b�h��Կ5ՎcY�����%���1�ҼK�܁<��G��Y�!*�Ǳf+�b�3�:4<�a��4��[-K�0�v���@�:�J�3Z�������D'igK�*N���@�c�e�2���Y1&��{�
���W�j�K� �ޢ;�9֣hY�&���1���a���]KM1��1��S���E��9��gxU���?;Ȃ ��z�(k�O�e�N��l�� �����i���n�ě�=�RV�N���3��o`��3�����Ic����n� ����{⾬_u����g���'�	:�� ��u��Y���Lu�$:E�GH��F�O�Ec�'^�;��g�>��8��&�\A�}O3�OX�Te���k���Eq�)=�)��$j\{4�� �dͩ��%u�%")�W�n|���eIRz�J6��e1����l���[�:K���бP�'ʩ�
l�U�_g�Ef)�^�[5��âȇCU�j�#K��w�p������HD�;9C�솀8f��jFe��k�|L��BR����
�5k�Qd���K�	_�H�#d����R���⃨i>]�Vg+�5�l~�)" �o�I��~�c��c��(Mk�g�l���������0��XO%��x
��<8�kض=����b�P| �Ek�]���x�z��&�
b# i	d��q����fE~m
Jl	��0mn9���	���m7���AY���U�,�8�M������$"��q��v�o���5�i�,�E�}޾�Ct�6�r�E���؁��4�>�1�t�JtZ��8���5f�	�Sk=oʘF}޷�#�py�������X7��%~���ĭ >3��Z��/1:/�xrk`U�?Bw:u�5�����rt��^�}~�D��_��3w:�C��W�L�-���C����4��H1�(�Rٕ�o�*�aէ�"d���cF97 &zM5%�T� �O�paD�����%3�֪��{;��<����M� d�YJ-	H�����;��v���G�	8L���V�EH/rmY���A9���;��l��3�ڛ�EB��h_���r=p�'���� �/�|��Sycz�����qD������A��g��ɒ�D�΁���2���a���dm��wV,IH���Y�鵾&Ѝ�C�8C��a��R��V�?`;Δ`h�T9���ٰP��QI��%�($4��߂�	�T}{;���m��x9�w�`B�>D���A
̲U�/i}F�B,fO���N�]�W�9�ؿ�S
�W�oX����7�k��d�1��jW���\�b�������'1����+Ad��	�p��L�A�Q3��Ê���1�D�v�A�S���$����	��C�'��x��.i�H�{�-����}���(]p���9�`�N&`A2~�=D�Z�' {	��TrP�S��Fު�e��d>R�a�����@.�(r&e� E�w#�N���N��i�������>��@2P+�]��Z�J�w��qt^�^^S�=���&�+��!���l�� k�t����s~z�t/'S&7��hL8\��WI���!�!��`s߻��Д��KU�*��M�^<�b�Ѐ�U��l��"�qyU���*�� �MQߕ~&J�U��n'�;�	�ں��?6��K���$4��Uv��'Z��,�J�yC��B
k�(­uF4�@�hOM��b��>�ߎN!����zuF�k��	Rb��u�ł��Rs�]�9�ÿ�B���ȉF���01G`O�%-�d����d�{n��Ԛj�l�-[z*���ߠSB�#��b��q�z�)�C�����[�;B�j䧡"jT2�t��~�|:����c<��%��F� ��Pi�{?*�U7���MA���.у�]�?�9DW[(!iߪq��c�;!R��\C��D̍5�m��/�b�5�'κ�P�:��z��C�)�=�T�R��T�_��%^���P��muI=���A�{䪹J�ь��r⢾��Z�\��i�7wx�_�a!��� �7$�[��|�|%���D�~p�I��s�iR^�����r������ߖ2V�u��^�4R�#$�Ѵ�Rs���"kV8�
J�B�J^�g�C�8pD=�8�S��'�YuΫ#��0����}K����V�V���	Rܸ[
��ղ�J�3�����k��QBa���J��MW��V��_9�b�GE�]eWwn<$�T�÷�l���;��_���d��o��C/𹋍93)�|��l5�C�v��z���,�`��'\;/9�B~D:~0������<�)2��d�"� y�q>b�� �)��3�?Źb�jO�ec�$����k�.�@� k�E�[��v�P�_�zP|�[Bc��Bز��ؿ٫��w��Ǫ��H��z��������_+Ju���D��;%������}Xz�� F�b�b"��8�y���fE��EXL.�������Es�X�sߓ%�3�M{��|�.����~@�_]ϩ�D�)�f�{ִ� ����$hA�$A�U�B��f���T�>��pFy٨|�C��â��U����"'A5@&̱�/�)���S��G#'N��1ٓLCu<��]D�v/�rt4-����&���{	>����<44a����5I�6��Gu�< 	�6SNyn���c�Z@�����E��I{��c����%4�K�u�W!ChW��5��Z�#0��
��dh��o�Ȧ���E�ozJ�U�+sg����;�,ȭ��,��KA���@s�eJ��H��\Y\�K���$�����>�"��xu���J0(K|�q�+u2<#��D�IS=�6^����b| _�e8qj�p��{C���¼��K�ݿL|����l���Z@/B��X����f�KI���u咝���\e��%Lf�ٿX9��}g˯�^oIv	Ѳz^ȓ���%?X��&���_���h�����a����{�Nt��4�c���	��-�#���OM&Q���[���5��3	�
[�Wƴ���}C� f���ǝ*��o�n Q��47*����	ݴ"4�f�/�K�~�x��Η܆���{a�����ο8��G��-7�!e��5f����#��R�젱�`4����c�s��<R�9R_�_^i��g����������,���y�t��0��Ug�"l�Tn����ەVA�w�A��tz&��RX��(�q���鰮/+�A�^����t����/�9�:�ui��2�������ү(V��)s�|O-���m�B�,fm'�f@�6(�[(Hf�MP����<yӧ�q��c�3�)��k�0�>��}���q��P�N�q�x�⃔�]�3��ܷ����v;�n���K+�!"�`�󾩓�sj�b��q7恰��n�M�6U������Y�"�n{���J�L�K����6�@��H��Hga֐��l1�n����qV~��J�}n]E��E���my�쉟"��V�)~��i����]ǒ�"�H�/օ
.�7��ɸ̨�|9�Oƭ�"�,��8D7�e�!7h'�<rq��ƴ�,]�)���D��2������+�Q�0���&^Y ��V%;��+�	b`�������U��#d����K��� �����n�pO�=� ��&��A:]؄�[K���x�X���R((	3�6��C3�p��ݯݖ�	�� {�R�h̷�Qd�T�`�&�6��\��o��ǯ�x�n0�q�y��b:�0Ƭ���Q�L�>OW�j�|�Qg�Жy�c���=!K�ʺ�gSO7T- �GQ�Ür�[�7���`�>�p(S��a؝�����d�N�-�J�n�]`��(�u�:��\Q&Yq�+�r����-R����]�T���Z���ڈ��2��Ź^���}�k�� ��5+��9��YLt��=���+@����k�j��&q�-\���Wn7;"��q�W�&z����Y2�$������nc�PS� `��A&�pMdȿ!�i��P�!�@\��@�!̧P֕܋v�QdPȥe��aw�Z���̝�"�}�f�K�?��Z5w�g<�0f/�oWi�'��"?��&U�4S ����|U	t   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸���r(K!�1�#l����_�)��ToڬrN�'|W�lc4�MS�i��(�gwGJ%
qAڲtva�V`o�,����D��	8ZZ��x7���l~$�aF��'*��[�'KJ#<A��v��c˔7-f�YA��ɓ.�:虖^�T���=$Lt����9?1�Ά�{�b7��\}RND����Q#�kubDIM�o����sM^�6
��	��yRn�.��g�ɓM��]�2���t.ܙBf�-S*�C䉁X�,LÐ�|en=Ph� X�dC䉗O�}� &��A���%ۥ4�xC�	
/��˴���#����.22B�ɹec��`vʌ13<�mh�̘�B�I}j�����Þs���d��%1�0C�	:>���Q��k.���E�}G�B�I8$yhM@�D
�!d��t��r2�B��<'��Տ��6>4�%�?N��B�.wͪ\���.a�X	r���l��B�	(�L�����{.TQ�[�&����d�>�q�(]fpX�	�)(�0�˟|Ex�W-��	D?�Ƽ���!M�n�Z%�Th�5�䐺�M$�I�{������>���[�\u�܈��)F��@!�[}��S�'�<!Gxr�R5h�Ҍ�.G_9
E��Kp�<yg� 2  ��$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Z    �q�5�oN�b�ǐ�o��h�"LO�L)����u8��'���J��T�g�.u��\�z��Ш4�.$�(�!    ���v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   �  �  
    	&   �m�%O8���b���8f��p��'l���4"S
�����?�)O����O��S�0��t	�>=��l(լ��h��m9
OX�����s�f�(w/����e��Px"���}���J)X0i!����&���9���?�J>1+O1�r.I�b�~!R��D������y�#�Z <cEfذ:!�]C&�)�'P6��O��`������2wꕈ|@��_�l2�����$�h�)�gy�ν(-��2��6���dA�y�GA��@)b�E�V�\rWgܴ�y���)b��w	�5!��P��]$�y��M�(ez��k�-��]��J3�Px2�PQ8,�벡Ԁ3�jUQG��>�tuF}r,M�h��uJ0c�8Q�pІ_}��x+����	CX��r&ET�'̐�$�	f��/?D���WBL�P�*�i�k��F�	r5�:D�lp4*T3��Jd�@�S� M�2�-D����D�.�+�Ğ�kt܌�!.&O�PDy�Y �Z��7jчi����'��/�~"%��O�I�Op���>��F�]+�8������@]�<��a̋b���EH�H\��M�W�<�@�e� ra��9Vi��nV�<)F�B�}2���peA�'���J�ƃQ�<aPm�i�(͢���J�Ɩ�7)��'�`"=�B�ǐ09�����9d���!�,�/Du̡�pj��$�O����<�'�?i�O���A��=S����r�E�!ٚp�)��2]�H���A/I�i�R`Q��8�D�w�'�}���S�3�r��0
C�;���bR$��?�s�iD7��O�ʓ�?��}�សrx-Ye�T�zU�$��y�
z��D�1o�x�)���<��':vmB��'��	�g��]w{�S�� a��
���r�)эn�:Ը�����?��E%�`QS�:�$�,-n�e!^�^=�$`ӆT�}ayn�$Ѱ�$��y��٨L���рGOG���",OX�+��'�B\��GO1z����fG$1�LQ׃����I���?���,��T�Q,ސ;������x(<�ዙ�f:~8�A��� Q��	b����$_*O]F�o��b�b�IS��+�hA2_09fKk�aS$`��"���'�P��e�'1O�<9"�s��|�g���_�AKuJ�L≙U��"<�~Rd������2��z}���!��G�I	�����O����b��A��!E���h篁�����A��kX�����Q�p�ݎ~�T탤�"O�5Dy҃��A�x�C'l�t���0fL�$RF���O�ʓ!���S�T�	�L�'�h���$&�z�v&Q(c�(��}b.�%��<����:t����A���qÔ��k�Y��5���.cj��С�IJ)�fG��q0�,�"�|Ǉ��?�}&��
#+��^���SRDRr@Vtqw�*T��'�Q��dq�&��!6D�B�>1�i>�'�`��L,�N�}�6��gm=id��s�i.��'��V��S������5`j����bCL��`�f.���l��=�O֠�&��0r590�1�B��.uh<�s�ڏ1#������t��	x��=�v���S�| �H��ݖs�N`��������!�M����$�OLc��@��B0^��'�M+q��'�"D��Eb�}q
��2����vV8��l��F�'��IPڶ j�4-�xpߴ_JI��e�����&[K�@��U�'N�I؟��	��|��L�:ܚ]��A~�lz���*وT+$�4�?d4Zr
�8����E��I��4@�bܵc)�T�łڠ��z7I���� ��@,iBb�Ê�$K+���'hJ6mv�X�!ďJ
s�4	�G(P�ę� ��_y��'��O���C��ƹ%��L�Q�(�L�k
O
��P,
�xi�g��7 jdHt�ûB�����<i�9�^�c�'���?᯻3�$�ho��N�"D��b!E9��'�"�\7�y�T>�*��p�怦W��В�&4t�h'���&�)�!e��{�̜�36�X���S�iT~OdԱ��'�2��D��$��4r��	�TA@.$�V1�U��5��'���'{��ƨҹ*���y aʹU�D��5Q���� �1/2 !Ǯ\3� ��c����g�u������?�O� ��ـ+Z��Ɋ�L�,'�3�"O,,�g/��#����L���U"O�����'V�J��JX6$	8�w"Op���P,xtk�� ��*"Oܔ*�\;sj���Ò'C�����>���)��'pE����$	�'���ǩOǬ�'��}x�'j�|J~��n�%V��Y҃��l����blB�ɵ4����ۘ#xY���:_nB�	*B�1k�!�D����γj�*B�*H0ၡ�'p}�Q&ϩp�>C��-B�T:pj�Uݶ��W�Xvp�O�E~2���?A��6=�@�v��5J
�S�QTxҒ|����ɤa���ܡ [�}�4��Ou�B�I�q���	��.m����-����B䉙h"b��.O�bY�<N�&B�I<G�~��B��u�E�B�R�\D"B�I#?�	ç.I)�6pK��Q9 ���T�I�l�}"$�T8_�i3u�_�W��%:�g�7B���'a}�,y�� ��k٦	��]Ytk��y�KB�N���>'���F ��y�l�$�T����C:h����� �y@4[+l��S�Ϟ �d�h���p<I��I��:<YD����]3ee0��	�}�0#<ͧ�?1���G�<
������<*�*IQ��S�!�d�*g-t��5/L�Y�:�A#�\�!�!�$�#|Xx�*A��+l�L2�@�9A!�ġ=���c�_�5nbp��o��o'!�$�;���e+�cN��nA��N9���?���̤u��W�W�$?�e�4 4}2@C'H�'�ɧ�.���s�ß�ȁB�1Q��u��;���{�K�*l����2Wø��ȓ]&���V�������/f0i����{�E�8?�̤J�	R|0u��{1VmQ�d�.x-���`U�qX���=�G�ɩB���ձmgN���T�X��ʗ+ZP!X���^�	̟"|�'��a2�׋s�\��2��<~F�@�'�B)��j�>Hf��1�ÿr�F)�'�4	��9ج�k
�w�\1��'���Ù1Hu�6��p�	�'�t��@_�iB�:\}\m �o�R�'��)��)U������^���8�A�_]����؟(��	"
]^�e���Q�Pi��P�VC�ɍ? \��Iȫ,�!�Z�=ӀB�ɼ<���g��	@*֡�5%T2-5B��]��Tk
�.��`�Q�Q���R�'ݢ-q���giz���˛>;z���'�zŰ��4�x���OZ�&��I��NtX[nR{^�}����`��8NH��ڥ��a������T�$�*�$h�#�*t���gĢ�Y6�S�!V(�6g	1� �ȓvM���C|:U��NA�dR��O܉Ez����O���Ĝ�w$<�Id��2��I��}��ퟴ%���|l�]%pi�Q��/y p��"O��#�N�a4��/̳��أc"OĘԈ_�S2���V@�W�Ri��"Ob���E'D�S�G@�d��"O|��ɻ/)�碉�V��d��$�T�'�x���a����:N�a$��	�6���'<�'���Y��F,��\���ѷ&̉Mv��7)D�c�ݩ3=ʬ�e"W;'����F1D�#$�3a�҉!���._p����/D�h9��24k2�a!���j��S��2�`
vmZ��D)��8��ǌԟ�Q�(�g�6�'oȈ�����7���U)�:P8Q��'i�֧� �� �!�\$؍ ��ؾ�4"O�u��Ϗ	?��B"�FN����g"Or�!���l J�*
��}@q"On �f� @6	���V��Y�'}��<�� T(&q~ȣ��\tX%��ɌU?q��J����'�X�H�6�G15�������wG��D�(D����<EB�TN�>�����#D�h��!��V�k�^7���	5�%D�L��]�nܩ�Ѡ��
��*�&&D��B���8*dy*�* �f�BP3�I8}��*�S��`�D���#W���c�I�	Y���OP�Hf��Or��5�����OU�=�歎�E>��(�!��yҢ�?���Iޖ;��@�wgK;�y��ݍs��+Q���n} 7*��y���%5
�r�H�u)z��Aɘ��y�JO6rx�x	��ڷ6~�1tFGĸ'$#?)��՟D3U,ɪ����D�6.< �C4�?iI>	�S����ʔe��8�S���^=�@���Łs�!�DӒkg�,z�X5	 ����F,0�!��_�J��S`��1g�&-ِѨ	�!�E+j%<l��A6A����-�Sԡ�Dʊ��)a�ڹ%���ω��p؂��D�.m)�>U�IM�1v4 k��Gu	��z5�N��?��ΰ>1vÍ������A�x6$�$�	d�<qՆ� V�9s�TZ�
%��e�<����,������Oᮄ���G�<y1,A,6���׉�;g���y�KC8�\ً�ĉ�{�=k�@P�qw�����)o���y}����m}��	e�BQ�`�Q�KS�|�D��y���rˌA�%�պ5����C-� �y2GT����!5�Ԁ$�̪�yRnSIp&��b�"v�\A��
.�y��ÂF
�;�M�6t�ryA7d���I�HO�c�1\�F�
6B��:�h1�Ւ>��[��?a���S�S�j��1B�ҏ8�=�/۱`��B䉕9�Ġ��`ӥa�t��Y�hr�B䉴^D����A2b!˔g�O>�B�ɶo� 1��� #Ԛ!2J��TTB�0":��H��L$���R�үP4➨ҍ��ޫr�bhN<̡��TZHfR�~����!�D�O>�EX��c�Z���h��Dt'���ȓ��LTj	$-�H"`�n40Ʉȓ+�h�9�%u�
�����OVl�ȓl��#�A\�)��ۓ$V�n{Bȇ��-"4Z�U�R��	�+RvHedN.�=�^xD��f#~�n�s'"�v�"h���W?[od���OB���\"t�Jmyb�T���'	J�(S!�D��A9�m�;���ŊI�1q!�dEj�搀�_��+p\�5Q!�d	5�H�`,�,'g�H!B�+K>�xҊ<ʓ�F	�' �*O�,�@�A�8�΍��~o@�Fx�ONB�'���6l�`�Q�sv�1�S'H��B�I&r�� ��F�<?�!�Q*ѧ/�`B��z�� ��L��e��O�� �>B�I�4� �ױ�n�˔�X�Om�C�	:) �$��@�`6 b�3V� �'>�#=��s��0*�9A�lSԘJ��K^�$�}Y�D�O�O�O���P�-��^c����!\�I��:�'��A1�؟P�D�5���Lf�\z	�'(�2Ц�"n�����C��@��'ඐA�o����T�t扣.}�dh�' lBC���r�ؤbO�nG�pr�{BH2�Mc"��	/l�8J5�m��U����|��������?E�,Oe(�kسg��`q n*"_P%"O� $��&ȉ�f]�mKc>J?xe�ȓx��QG		[6�E&M�.0� ��6�$� `��>O+jM�-�9�⭄�R<��IքE"	1��ÌEY�c%� b��G��	�U| �t��J����&Ƃ������O���d?W����c��5��)􌋘R!�D��  ȣUAR��=�I!�$� y/�𘑢�	���%���!�D�*�Q*U�ć(F8�氄]�Ǔ5ZQ������� I�DG
 �8�⭟���%��|���?��O�2��Q'<3Pn�&�cR"O6%q���$+L��sJ�����"ON(� �?ز ;Ui�%W�t��6"O��+p���+��SRۢA�eB"O���Č!C�h5��aG3G�4Qǚ>���)��
d���lv|�Y�� ��w�@�'�Hq�'���|J~ʕBбS8!iF�k�~U1r�ZJ�<����(�=ؒ�W�{��A�gÛC�<A�,
����X�j�D��c�d�<�bb@)PK���F�"&��g�h�<ÁU��fŸ�OO2&(L�6� yܓr둟�ѷ��Oh4+�+ez���q�\5r��Xp0�F��&�\�)�gy�@��l4�r؞Zd<m�b\�yrF�%1*�trO2R�2,qw�V�y⡟�qh�|)�#M�v��s�.�y���<�:�M�:LWjaj��Y��PxoT.�
�_�W��a
Ԝ��F}REϐ�h���д�Q�$�d9a-¹�����X͟��IRX�\q���=f��K�'��A�聠�1D�@Z���7�rue$X'%��9�"D��9)9jl5R������葃%D�����	'��a�s�H�HW�H�O9O�qEy�͏M��+G�� *~5��	 ��~R����O���O���>��l��k#��B0�Ҵf�\����g�<�a䏅/�mbQ��*Uz�rPF�_�<��R^Tض�)EA�B@�X�<���3>0�Uq�ԫ����@kAj�<�	�7cj��D���ˌ�B�l�d�d���Oپ`X%�=6�ɓLV����kJ���d���`��S�)��# ��q,�Z�.�I�,�6K!�D�?W
��#&KU+L�b�� ���A�!�Z*κأ�,���*Ua'Q�,�!�$�v���ƛS���aGF�6CW!���7�X!��]U'��x���p-qO��G~2˃4�?ys��{�(L�p�ʑJInus��������?E�,O�8 eL�(e0C7uZ�X�"O���c@֜?��2���;\d���"O�X[�ƔM��=�㛻fD��
"O�������+�-����1%�ݲ�
O��eG��f��w�N%(���y�Y���O�|B6퓃Vl�5"g�B���p�����D8`��?�	���*#�^8hӤ5�udX�!�f��;��yw�[�f)*�D�ܕiG*Ňȓq��!@m^�:B� �T�#�<��|���2��'���P%ƀ	�l��	;�(O�L@�C�8��MzԌ��{��R��O�9�3�i>I����'���� ӦK��#7�_�t���3	�'^nLB���8��1�f�,ji&h��'x�1#�?�hTH�!(_0^���'�"��(���v�ߞ^�Dԉ
�'��@v�D�<���(R3nꪬ(J��x���)�)AKT���e(�@]s���8
@�W�&|����?�M>%?����Y��l؆��28A�� &&'D�,�e��M^:9B!ς)?����j#D�� h�y"�R�Ā(��P���1"O����5o�<ѩ&�{8���"O>���N�E?(��g�o
����QH�';����7}D*b�ڄJ����D�e��x��'��'��Y�@�0��,Lp`kC��"RQ���!2D�����?}rʤ!$H9Q?n���;D��a�O�50�e���D
u4x��<D��0�#.�����H�,�6)��<����"ل@c�hi���� �i��ipQ���é4�'3(ܱb�ĳ�\�
�$ႄ1��'a��'(<�*bn�6A8�!�c��/=�E��'�,E�3E5Q�6����
�`c�'t�"g-��A,���o	�-W��	�'�Tm�FJ܊2<v�H�@�'���k
Ǔ�Q�к�n��&�!�F�BM��ɐHR�I�6�.b�'�lu���r���?��OZ](��Z�X��U��B3�Q��$"CT����F�3�ZY�|&��sO�_>\�X��K�;Ǆ����Ԙ
��p���X�2�b(�C)D��c?OFq���3'W�P��g@���\;af��h�'>����|�����'�"�2�"A#o���vB�l��1
�'v��f�K,
��p��Z /p0�I����4����>�Gd!��Є�_,FXbe �ҍz��b��qӮp2g�O��D�<1���?٘O6�- w(W-6���`��=@�x�W�ȟD�U�L�-4zR]��o8���䑶N+�����~ˌ� RKR"j4�՚��F� ���nA��x"��MP�0s��ճ`O��G��92wz�	Ο@E{r�dʵ1�pH�ЁJ ~[v�^���'�|q�%߰��ʘ�9��9ˍ{�#v���$�<ٴ�����!������ �P;(�#�I�C�@�<`?j���<���?��O���k�FNv��� ����B��1�zaZ��^�BNO@Cb��D����p��#���Dt3ԅ��#u��\�\�0����C ������9o���$�Op���wCT�C~p�r�O��,�=i��<)�o��z��q�t�"N�piƆ�t(<�N֭e�DI�Hϣ6���$�-d���R����$�n��)n�\y�	O��5�V?#��qA��}q��D�U�Pn2�'$�mI���P��E@�@�*DDl�|*��@��n�:T�6��`3-���X0�x¤��Q6<��fZr =�=§Pft�t�+a�Ij�>�.�'��� �O��D ڧ�M�b�Y"{�R�a��M�t����*!���%�(�S���p�����	��xҡ>�"��c���(fX��ٳ�Vl��s��@���O	��'�	w�l��v��-׎�(Ԩ�QZ4B�ɛg�`0d��>ydi�0g�%`$B�	�]��XЕb[qJ �	��VV�C�Q.j!�v(Ì;��$�!� IRhC�	��>h��Ծd���b�$��DxJ�'6�"=���C߀n&�T��j5�Bh�c��b�
������OR�O�O���[��]�0޴��Я/e�DM �'�ȵ�Ե߮89�
��b��Y�'��Ds�
�u!��#S�:`�<��'�`IA��zF
�KGJ��RC���'Zr��R��=9�Y���>J��{�.>�yT���ɃD����Ȍ�[�X)9J v~�=H�����?E�,O�Y�'��1fT	���T<�h�U"O�%�G��W������� 8B�"O��ä��5(�y����0�E"OH�@���D����K�]x
O��[�(�h�X�R"[�	f|� Wg1��O�{a�/Z,��@
>m�&X�	�!��J��?Q�N���+�3�$ pP�B�L�,ф�j&��ǿYJ��2�<����ȓ��(jbJ�<;�r�a��T��u��R쬝+�,�.j.n���BB;U-��I�(O.Y��k�/��˰���* �m��"O��z�@  �G4���'��ʓ:�Pg�9r�E{5,��D��?��.Kw���$�'��e��сs"<���LG��VL[��' !�V�t��U��Ί�&�D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  5  �  9  !)  "4  ?  J  "U  w`  Tk  �t  �z  ��  ��  �  E�  ��  �  #�  ��  �  ��  ��  f�  ��  ��  G�  ��  ��  �  �  ��  � � # g 4$ �+ 3  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9�ӄZ���1.*��5�����5	��9���ͺ\4X}�]�=B�=a0T��&�U��8�e�� B�=p�>1{����y於m5c��C�I0d�����̈́ -�\����C�	=ڴ���M$k|$�QT� !��C��2G��l���5[p���C�<�u �
�X��/���C�I>0��[3㔶%��}��j�5 d^C�IvQ�ղaɌ#��I��^@�B�	Z̒���Cv=@T��&_<�B�IK�����,�)f����ס(�B�	�3�ztx�G��J��u��/��C�I�	��,��̚0����F&l�C�&	��M� �FU�<yFb�1�����>Y�B�B��Hɐ� )7�T�u�c�<� CR�*�Ny�tb#"t6��d�d�<�&$�{��4 ��N�i4���(�W�<It��o��13aԬ��<K7h�L�<q��Q�-���34D=@����D�N�<�W���=�����E�v��@R�TH�<���$w�t��4^X���
K�<��mM	a��(F�}�nD��a�J����<A�(N5+FI�'J=���L�C�<q�]�+/���B+����At�X�<��'n/,ds$\�X�x��@�^�<!pj��V�r9�!�!h�:��ee�<)�h�=7��j��o�)�a��a�<9�C�<Ϫ}�W,�(6���R娆[�<1��"��ݱ�#�d���S�T�<Q�'�ޠؓP�%P�L��bK�<�qA���a��]�\;t��F�<��� ~v��`΋4�@���DB�<� ͸�dH�j\/{8����-B����>Q�E�FW�A�`���~�0 mN|�<�1T� �Q�.�VE�P�O�<فn=<���&�*�L1�GGK�<�A�Gx(���21q(����[�<� "�X�'�z�r�I�,Fb�	���`��+���O虺�畵 �P��a�^��0b�"On�����#*JpJ��� E;B�)�"O �s��V���p���+�"�["Od��ŎPG}+6
�qZ0a3��x�)�Ӓ4��6o�r���c���0oD#>i����_5bhzKҤ%Z�Ti���
c���	"N���q��2����/.5���hO�>yi�V:*^�`t�K1N��Dsf�(D�hZ���	_`hd��l�v���AKf�G~��.1�����C��]>��f�?e�R��o̓�P�3U�@�]o�r��x�%����.
�P40-ۃTH*���QȢ���q�\I�OJ�І ��
m�ʅ^"W��J$"O���+���09c`[#�iV��t>qB-@Kdb�:�]�@�b-/D�D�W��T��d�S��4�)��/D��� 	^� ���[%�];`��e�B-D� sd�Vr�d*Ĉ5::ta�!l��C�	5R�p�і�	^��XIW���˨B��6/d��ᣊ�6lB�BNآ�ԙ�ȓF�X�f\��2|!'J�"D����	l�'Gt�C�.@6��-�2I�/��h��'�L�AB>o�B<y�/̕*�`x8�'�2� f��/;(��Ke�
�79��'���!���T`����ڪ����'�h�ڔH�?ӈ�Y�fK�Hp�'�F:�×��@����E���'������R<�CH�.��y��'�X���f��e�X�G��w����'����ȋggԍ�$!Η�.�'��1H�$��"Z��H�U�	x!i�'�r%Z��-�4x�Cc��}��a�'�.�1A��jZQ3s��804�'N������.r��43BD5{*(��'<4��W+�-�L�a�۾[c.Iy�'A��io^|R�)��Y>ʬ��'����F�C�Yi�@�*L�܂�'�	&@�k�T85H]�z8��'����ː�bp.(aDMH-	���3�'mf�
�V�/�x)�p\
N�+�'���Q$��2:w���wH�/Gbt	c�'��B�7	�x�xb���g��a��'�u��i��Ok=�!I�0�zI2�'�#���
���pf��QPz(	�'�d��i5r���p-�^�`��'�:]Õ+�m���K���+��d�	�'.̈b��׺g�v="`aR�R���{�'�j�{��I�?��j׃P,LX(�+�'p��	�	Au��[�E�1z
�'� #��˯7Ü��2�8%��	�'���1�)x
�� rB̭Sy��z�'Լ�8`刣m4�����N#�$��'���p��ɉf�j�� F�6�6��'#�4�v�N�+<N�� � �4s�Pa�'�ri�2)*/w��q@�͐&����'��`����*]���7��v��0�'>� ����/� ���4Č!�'FE��oì�$UkSo�	8��q��'��2hJ.h
S��0@�yC
�'պl�u�T�����"h�.&���	�'M�Q��@AL�ܺ$聆i �
�'F�]��IϭLX)��&m���	�'�f\20��2k�$qb��\�hϞx���� �\CO�0&��@��0�Đju"O �n�/�*<#�j�(v���1r"O����A*h[h"�/��R*mq�"O�i�V̖4����V5Oi0�"Ollr4��S�č�d�� ?��a�'p�'2��'QR�'���'5��'~��K���=k@�3��F6Q���'?B�'r�']B�')��'n�'1�Q�N�Jc�8ô�̽k��m�4�'o��'���'��'U��'���'a��	E��7+�1�aL��h��AxU�'���'���'���%��� ��ß�{�O�r�`钥��#}�$:Q�Oԟ��Iɟ���埔��ß��	ܟ��	ڟ8�b|8� u(Tzw� s�ҟT�	ȟ�I�<�	ԟ@��۟(��Пl9�E͹|�RٓТBH�@�Cϟ��I���	ş�����ß���ݟ��G�#jGr�R*�%�ȴ�2�Aҟt�	���I埐�������ޟ\��ԟ�R�տY�
�k��� s���t��� ��Ɵ���ɟ �I��@��ٟ��I�8Ȗ�+9P�������He��"埌�Iퟔ�	ǟL��ٟ��	ڟL��矴�a�!:zb�p0G�� j��������ßT�I˟��	��	֟��	��rqBܜMsب�g�X}�L���ן���͟���şl�Iڟ��I؟d��՟������|+DY BDٛ}�&�ë�ß���ڟP�Iϟ �	����	4�M���?Y�ԋ]�´R��P�d{���� �rK�I�蕧���d�)� �Ͷ�H�C���To��1�n�h�'�D7�(�����D�O,�I C!���JTH& ���O����R67?��O5��)5��ݮg/n�dC�#l�5�qh���'mbX��D��^�e|�4��������pۼS������OB�?5�����v��57
�h2$/S�d@��"L���?q���ybV�b>=��+YԦ9��:�4�@5\^S$c�R�M��y�E�Od�"��4�z���r��SG�@���s�HTu��<aJ>�u���O��9�C�mF�P�'i�,"���p.*�������Or��s�$�'u��S4,ZRp
s��=�:9��O��H&TE�uz��	��?q���O��q֮ 3ܘx`E@�;"�TY���<y+O���s��K�+�:��CH�b��f���hs�O �	����4�%Y%�e�z��BK1T�z�	<O����O���
;X��7M2?�Ok@�I��}�����"����C�P���I>�,O�i�O��$�O�d�O��qB��oHͱ��ߒ}�b�b�N�<�5T������h�	c�S�� #�gȖ j�L�2�F8*��`)������d�OB�D+��ϔ<a�x{���TF�{2�2�X!�̈́�Bj�ʓ"ʬ��5d�O��I>�-O*��'�13�����6'Tjxb��'����?�'޲n�td��b ~6��q���/�?YA�iX�O�}�'|��'~r�L[Kʘ���;T������.]�)B��i���D���)�ן��������%��` �I(�`��C�QA�.�O�d���#rl�&n5N(��l�O����O�ԧ�i��)$��g)ԾKT�{�([2U�q;P�a�Ip�i>��������u�,T/3.�q�.�)z���$,P,#gt�B�'��'�d�'��O��������ڕ��2d��"��I9���O��d�O��'	�ZH�a�`@��� N-_}p��':���?�����S�D�(6f�d�2Ϙ��H@��ne��cs(�0�N�<�'K���`�30�H1y�!�+#!Ju�,�P@�Iڟ���쟴�)�ey�j��11�Z�B`�a��RzI���C;O��1r�6�S^}r�'�6 �ԁֲ!�(M��ժ�:6�'R���LM����l��iȠJ��~BAA��C2u FL�B�T]ǀ�<,O
��d�CR��)��ՄjJ(��L�A��'�R�'N�	�Ѧ��z%�A2C�
 e�d�Z��)j��	ğ$�b>-�"@���L�Rق�́� 5h`c"�6'�ΓHɜ(�@���$�T�'$�	!w��#1!^'l��9窀�
����dE}2�'��'6��A��<����dC3w=d% C��Xn}��'5Ҕ|���&Dx̙�%[�����c�%��dK�%�����dӠ@&?����O�����ن�;JDL`bb�bF���O����O���4�'�?���О:�\a4 ������I�?1�P��'% 7$�i�)�V"ճA��A��h;�|��sGy�<�	ğ���V��qoZV~R��,_����'X�
J��ѼO�t4�Ũ�+0�a�M>�-O��O��O����O���I�#'Fe���]�z���H�<��V���Iҟ�	j�s�0��,g|�Y0�Lф}���*FΜ-����O&��7����5B�>�s���#�Ik�HҪ{i�i2q�P�I���A�Ʃ�<'�$�'$�耵j��5R��hp�K�yPB�y2�'���'������_��r�O@��P6䲰�f��c������'0����=�?��Z�p��ן�I�Bx�q˄�A5>_ҕ@���)E^���Tצ��'y�|x���?�`Й�t��� ��ATn�|��hn����8B�2OT��Oh���O���O��?!��ς�|ysF�Z
'��d{���T�I��H�O�ś��|bB�
��ѕ'�^�ޱcs�ν��'	rZ�8*��ئ1�''��� ��)N�$�"�!�\��Is�)B�~���/R�'���ԟt�I؟D��>�@U��םj���rUA�2�����ϟ��'"���?��?�(���ʔ��*h�A��	6`IB���8q�O��0�)�釘 ��Q ��y����V�P��	GLV�f��-O�靱�?�AB>��Q�`(��C�'d؅�2,��:���O0���O��)�<�U�i�� P�2b�p=#�d�4T@Ü'���'��6M*�ɑ��D�O���-� y0�!� IJ)��g�Ox���!Yx6-7?�%C�$J��S{y2@��ᢼ�Р���#bkӟ�y"^�p����������I�,�O �0qt�\;��H{4��L�PE)�>	��?����<�1��yg�ʍ!g������#<��� 2�r�''ɧ�O��(�Ĳi��$Lz��q1�!h�у�X�_l�� s�J�'��'o�i>��	';�>D��C�+!���4��6�����џ�I埼�'w���?Y��?Q�-Z��BR-Ҡ������'����?���|m��+��C�Co���@\�'��1�'�����J�gR��#6�	�$�~��'J`���*�pu
!EM�Xd�M���'�b�'r�'Y�>1�	�ºi��A�O
���.Y�	���	���$�<qd�it�O�G�H���R���!�S�\����O��A�0��ڴ����/�.����Ef�2��ߎr�@��.@�-�bQ9H?�d�<���?���?!��?��L�`�0�Z�-��,k4�bW�� ��D�{}�^�,�I@�'^�D�`��؄�v�+挘�%�h�3R^���IA�Ş#p��r��66�B��e�ɲS�B(Ią˶"�� )OLM������?���-�d�<�%�*:�|�`A��F,���U��?1��?I���?ͧ��G}�'V P����!(���c��X�'�Z6�%�����O���O��F�H�D��1CԈэ`��ũ5�L=��6�/?	'�2��i0��ߙ��O*bD	�s�+&� �`�/d����ҟP��۟x�	����R c�gHH�U喳!�j��6 ��?I���?�CX�(�'O�6M.�D�G]�q��
� Z�͂ ,�|�O�$�O�I���6m'?�!�[RV��
�ꎵ^��
"儬�XE�u%�O�XCH>�-O���OJ���O<Y��*Ԝ	Xң>;��e���O����<�V�L������Iq����	ca�~ݸ#�����Dd}"�'1��|ʟY���:F �-)XHU1I��_��a��j�B�S��O��O����͸	��@СK�'D�d�83��O���O����O1���:�6���_�	����V�V��wOX��y�'� t����[�O�����i~`�p��Q�`��e�]q����O�	�Ox�,�X�2ƴ?��'Ap@�W�Iw�<3�lV,���a�'����	ٟ\��ԟ��e��g&<�^�qV�R5��퀄˂2Jf��?����?�K~�!��w�а���OjJ�N6B*�Ab�'��O1�N���l�p��%��X�A%�*���h�3Zn�	�e+�@��'��&���'���'[(dAG������cǨ*VdXY�'}��'�W�0��O6���O��E��}��١2� <r7��h�����OV���O�O�@��A�<!w�	�-�#q|�u����d[�<��$m�a̧Exx�	ߟD! ��=tQ��*��L'E)$q�cڟ��I� �Iߟ0E�t�'���r�P�@���
*�p�K��'Aj���_��?�;C7(�s�f�*3t ��^�����?1���?���M�O
19�冫��0�;�����
�Q(� ���_8ΓO"��|���?���?q��7���\G�t���S@49(O~��'&�	۟(�ZqBMj�y`�퍉	*v����h,�	۟L�	M�)擝`�D�2�%��&CT�"�֕zˈL�'sS��*�6!��O��YI>9.O�xs��,G�z��XA�|�� �O��$�O��O�I�<ѕW� ��? �θ#�*�5p�*p#�#��:@��ɇ�M��R��>���?���a@zq���jJ����J�bt�!�M��O(!�d�Y�(���N�7�"A 8a\�m�G�K0`	��O��$�O��D�O��<��<Q��y�V&�?d\	 E�¾L��������	��4���$Qݦ�$�4Ra��8[:$�Y���3��0��c�	����i>a+" �Ц5�'�T�ա�3����O�=\={�%��@
H-��䓄�$�O�d�Op��ώ\"L� ��0P>�(9�-]�_o����O��l��	ş8�Iӟ��O
�� �-S�c�\qÑg��y��OH�'���'�ɧ���02m&��6���m���|,*S��X+p��6�!?ͧg���It�(
6h���)YRI*��~�J����4����)��by2�d��Xs�K�+p���E5`�����2OR�$�O�yo�_����I���Z�g^�a��e�sD΃#GШ0�Ǆʟ��	_��lf~g�mV��SS�� ����A[>d�b�pQ'I�$Tz �2O���?����?���?A����/渒��ϿdD��U9��r�R���I�����~�s�D����CcЃ1I�1�����įT$�?���ŞS8ԉ�ݴ�yb��L����n���
1(���y���n���ɬ��'��i>��	�x���G�DG��!2�@��8��Ɵ��ꟈ�'*���?9���?��������Ƅ�B�&"X!��';R��?�����7�$�E�7MW��@.
���'���@�b	-XKd���#��pK��'](��C�&:���'F�1�,y��'��'P�'s�>a�ɷ ��b-p����ɠ~��H��&���O���¦}�?�;%��l��O�(*��	��:�~�͓�?����?���M[�O��0�p�	ζS��)���ʷ�via�"JSJHAqO>Q)O���Oj�d�O���O�A	ץZ ��	dc�|t)PN�<�vW������d�	{�s�|p�#�)Hm~�h%�5
9Zu���F����O.��*��	[U04�ËV
�a���1*�*�� �F#>L���c`"aڅ�'v��&�h�'6�A�pqJq `���
��q��'LR�'*�����U�l�O����PZR�
y�H-�f�Y����禍�?Q@Y��	Ay2D:+Q攱��>Md�)F��3xq敃�i�I;��%���O`�$?��@�� ��
AF�I�*X��j������ٟ��	ğ��Ix�'[���VI�<4M0��샯'h�@����?!��6��i>a��$�M{K>��i��U�ѡ�a�	F���4���?���|"����M��O�h��Ď:50e�#��?�Pi�%Z�b��'u�'4�	ݟ��	՟d��	.R`˦�<�k%�Z�G
��I����'hZ��?y���?�*��1Ѷ��(Y�}�  	�q�v��"�����O6���OD�O�S`@p��N�Fv��#Z7C��=���=�i`9?ͧNz��d�2��Y a���h� 
3d�Rpc��?���?��Ş���Aڦ)#tϞt�����DD��|��'�66M>����D�Oxm��F�D�V���a��m�!jd��<�e��M��O��+�:��vh�<ف+ٮ ���
Pl�5D8�@��<!(O��D�O���Ol�$�Onʧ-�@M8��<�ҤSI�~�\�R#Y�(�I���IV�s�P����&����	�Ax�"��5bA����?9L>�|24��*�M�'��Xs��CH�*�Ÿ1�,Y��'�8q:�� 韤S�|�U����ѵ�2c���!Jԑ2E�|��XПd��ןH�	{y���>����?i�A��:���!Owl,Rb�F�[�^���ı>9��?qJ>�3-YJ�N��&�";b�����g~2�M.EyJU�W,���OoHA���7y��^ �ܲBoJ�>��<�������'���'�R�s�yc0(�"A�C+A;V����
G�����O����OHl�n�Ӽ�Q��G�! �/�H�tkeg��<����$T�	c6�,?�T��StL�)��R�z��K�ji�̃�]"�\-2J>�,O����O����O����Oش��NΏD]b(��.�:&���D�<�_����ҟ��IO�s���-X�&�Db�.�Tlju�Ƨ���$�O��$+�󩟾�n5sp��<O�Z�HeM�^O�"P3��	�-�h
`�'.�$�`�'���Q��Ń+��zC��Vk�����'���'�����Z����O��$�3&��Ta�!ąQE�#G	�V�d�צ��?IRU����zyb�+ �a�l��� ��rD9a��i
�ɓ*2����O��!&?��&+��p	�0c��Ep"g	�t���Iן8�IΟX�	�L�	z��:��q�5!$%�FCSC�r��ͻ��?1��.�I]yKwӲ�OL1�苄h���z嫃�2���G4���O��4� �3jmӜ�R� �� �e&1C"��\j��8�eșe��$�����4�,���O����:��ROO�h�R�KR���gn*�d�O��N.�	̟���ȟ��OB�5aWFQ5!"�;�I�@|0��O�i�'�"�'mɧ�IS�s�$`�a�-*��B+R�H6UHv��k!�7M;?ͧ]���V�ɰYZ���%o�N���LȿjY������I���)�py"op���!ϕ �B�2 Ńa�z��?OT�D�O�l�M���H��M�9��a&�ߎ}g��a��l�d�Op��0
`��Ӻh���j��<1�@#kAv�k&��!bj���cV�<�.O����O��D�O��D�O˧b�=ywO� ^�J�I�⚲.��Z���IӟD�	p��Sߛ�wm�V
�Z�ty�!�Y�&H��P��Vß�	w�)��-c�Ul��<Qs��B����b�_�A*�����<!��#����Z�Qy��'2��;/|jUn�} c6�DGr�'�R�'����$�<Q�>��`�β.�v�(���"̾>����?	N>����b��	�d���M�A~�)�L-�� e/�{:�O:�����{s�NW�8nɂ5�Ϋ@�p��#�r���'�"�'0��S��x��Ʃ4�:�{��Z�x����Y�LʪOT�2�f�4��r�Q� �WLC��ͫ�4O����O$���F�7�4?����A���3� `p�"�mҲEGMӃ9޾�a�I �$�<ͧ�?Q���?a���?	���"#����:6����)����R}��'R��'��y��]�a)�5�3�>p|2 I�h["V���?����Şg�ڰ2��C�L��	2�1 J@P��Ć�M��O�(q@�
�~��|�V��c���t�\��֗O��D��m���	ӟ,�	ȟ�Cy��>��/�8�i	�ah�Z',�hN�<�;��&���f}��'Q��'e�@+��	�q!����� P;����M')�6���@B�7�Q>����0Q��C���>�[��Q� �
�I�����韔������j�'>�L�PT쁝��ir3 B�#]�����?��/3�i>1�I1�M�J>	ƣމ,��-$W`.��$.֚���?���|�P��M�O���vBUK:(��0��Q4�0"c#m�Nq��'��'��i>%�I���ɠy���Z�EE��pb�o�b-������'*���?���?�(����d�{x�{C�F�P���)�O��D<�)�V��!2��mK�C�<X����%J�k%�W�pz���q�DLy�O�����$x�'?�I��;T� �� ��#v�s��'u��'X����OB��Mӥ+�H��y��Fޞ"���w���<����?�E�i��O�<�':2뀹gQ�mҐ��$1��XA#߱+32�'�@չѱi��i��Ы�?qA�W���!M�
t�b�]_[��bMi��'��'S��'pR�'��S�n�j=g@ʊ"5�(9�/���D{}�R���	E�Sҟ$�������е�(8#������#^��?Y���4�?a�V0O��I�_:_e�3����Z.vE�v>O��CT�ٱ�?��B>�$�<����?���^0˞|��� Q�������?a��?�����~}��'��'E�M����U����N!j��a���o}��'�R�|R��
j��t"��ɂgL�;E�'��d��;�I8E/�	KH1��M�NH(�g��G�*,�D���ĸWZ����OH���Op�$=���I�t�J|p���ȼ�V�?��^�����l�ܴ���y�H$6t�XC�l(�IX2(�yb�'d�'w�, �i��Iu&�pHD�O����'s�x��� bX���@�i�	ay�O[��'���'��ǭvت�q�eRRj$R�f܁Lm剛����O����O��?ͩ�ҀR$m��I��C8���K"��d�O���?��	^�P���Q+)Cv�h'%('�����bӊ�'�@9 ��O?AN>�.O�e�2�ĨE����c��|B��a��O���OH���O�)�<�$T�8�	�pӔ1sDK.cB�q�ę%"������M��̱>���?��({��#�H��X(ȩ��]2 �h�����.�M3�O���'��������d�w�X�+`��[]�!2��X.,1�'���'���'�B�'h�@CQ��Y�!�	�	�B4R��Ot���O��'V�I"�M�K>Q�$�ɬ9ZW�J�ش17�"���?1��|*%Q<�M�OV()$e0f�ZԂ�$� �	�6�R�8}�C�ML��O���|R���?���P9tŀ��R<谰��:2������?�)Os}��'<��'g哐�XѲa^+�����l�+;�	؟�?�O�l�����1rQ ��2,��tA`��"	��mj�%W'�i>����'h�%� 8��d��2�ځqx��q�%@�����O4�d�O$��i�<�q�i�.��Ň���J��cK@�X'x��'G6-#�I/����OP|��_J�����0����W�<a�(��M{�O�E5���"��<QB�Ԓ<�M��B6P i����<�+O���O����O��O&�'+�H9f酩!��hc`�-��U)�Q��IڟX�IL�ڟ�:���%�O>sj�����$�"e�ׄ���?1���S�'>Ř��4�y�O�QC�l15��D���A=X�<�ϓ }�u��O��O>9-O���Oft����<O����9ʎcP(�O���O<�d�<�eY�l�IڟT�	�eP��`��H'��A�3��|�?!�V�x�	ڟ'�H��L#4�l���3_�@�[�`9?�$��/?X�bܴZ�O+|����?Q�͛]��)�E��B���:A@�?����?9���?I����Ob4 
m"����4�@��ԣ�O� �'���2�M��wT %��פ2���#ʑ!�@D�'�"�'<���?�����ra���4$ڭi�B邦�C�@{4G>��&�L�����',R�'�'0�X��(�_A�Y��Cʡ+����WQ����O��$�O�$)�9O�4���
�E������<%��n�Q}b�'|b�|��D����Ccҵ5�P����/v���i������9�7�Oj�O�O*z�)C)1�4u��,	�K8�I��?���?���|�*O8��'��CK�V�~1��]��yv�Z�?r�v��t��O:���Oz���I�rI �
�(~��� ���{���XxӴ�b�n����?�'?����\ԓ���<�(�K� ��B)��	��D����Iş���M�'9Ů䒲��'{|Xa�H�F�!�+O^���o}ʟ��mZ�I v~�*vȅ�D3����*��/��c����yy�+MO�ƛ� �'� �C�G�?(>���P%Ht����A��?у�:�$�<���?��?a��F�+�~��uF��c�J��Ё��?������EK}"�'���'�)i$^�Q"�0N���̊�'dj�Kj��Ο�	o�)���8-����C����aZ�@S�i{*��,>��L��T�P��|��:{;|u�b+��Cn�``���^�b�'���'���dW����4u����'�!nT�١g� %.�Γ��DYܦ�?��W���I�6@Aٱ��+7gzl�(N�B�	֟�����'Yv��Y�'P$9���|?
9$A�*?,=�����O���O���O^�Ĭ|���O����ռ.�l� ���0����O����O���3�9OX�mzޡ$�=��< c`ȼ(DX�r� ꟼ��A�)�Ӈ�f�o�<$��#
$1�4��>8�nR�<9��N���������4����pfH�t/��N�8���H�>���O��$�O �k���ğ\��ğ�c�
�!�qTL�P�ڴX�x��k@�	��Io�%BJ��!'$��h5���C�6�&�2��L�s)ǍG<��|Rc��O����M��=b1�!/���bu螋Lm0m����?����?���h�>��ʑR����F��,����AدD���dp}U��b�4���y�ᝬ]ol���C="�Feh`��8�y��'�B�'L�J�iK���QIH�`�O�v���I�6#�(9��lB�p���봁@[�|y�O���'�R�'}�֜id��'��|��ľ���,��D�O����O�?Qj�FK0C�Lh����H����D�O��D#��):�q#U�N��u����!UD��s�tӊ�+�if����%�0�'��Ёd�R'T�s&c�+|<��'\B�'�����W���O*�Ĉ5g|�C'gF��NU�*�����P���?�#\���IƟ�]�nvV�Qwi!O�^Ydo�>~p�Ѳ�����'��]��[�?u����d�w�xh#�'%(�[��7L_ ��'#��'0r�'��P�b>���+��jqb	�T��Ο���L0�Or�3�V�|�j�;s���i3I��a,a�-����'F�������ʛ6���Z�ܹe��� C��R!p��J�T�&�S�O��O���|���?���c��+D'�0j|�)�E�XlA���?�)Ov�'��I���Oj��	��?'�q�bͤ<*@J�O���'���'
ɧ�	�< �D'�"ư�C5`Q'L�j� ʚ^=��xb���5�R�FV�	K��$8����QJ>���Ĭ�����˟��	�P�)��hy��tӎ$�.I���Y!��%$��P>O����O0-mD�1@��ɟ����| z�"��MN���i����I>x�f�l�C~��^��������߹l��a�u��5X����IޱQ��ĸ<��?��?Q���?i/���b��,�����$��
�m@}R�'#��'��O"��q��́*�!�̆=uI���,��y�Z���Oh�O1��q�fӚ�=|����a �A�td����;�`�I�F@%��O�O���?���c��1�"	�l�fd��j�$X�����?)���?�)O�u�'���'��A�v@���m�0�2��K�O���'�����G��@{��S%<�DQh���Y'�ɧJN�E��XV��Y$?e���'��}�I�|(N��RHS:�M@ei
�5r��Iڟ�����I\�Oj�Ϗt%0@b��\�r�ڑ��	�b�>1��?9P�i�O�.ŌN疴��*'�ns�AN���d�O�ʓR�\Y�ڴ��Ć1<�L��'L�Z�:��L3H�ӥ(�Xh( �<��<)���?����?y��?�0!�[���Q����~��p;4�N2��d_v}2�'��'��O��B<0�:�F�>q�M�a/�p�8��?����S�'t��t!ɏ*_-���6���~�~�x�`϶��h�/O��*�"��?��7�d�<��.
Z�����A�;���tnX��?)��?9���?ͧ���Bz}r�'8���q���br��-�j}���'�&6M �	����OR�Xk�!ÇcE808�D����ѡJ �Mk�OPdx2NW�r�'�i���A�+�-��-C���"�.�$>O`���O��D�O����O��?�Q�N�4��S���y�*��ܟ��	����O�ʓ!�V�|,�#5a� Ǿ
�����ǋ6\��'����D�Ќ]o�V���J��(����ꂋ��Tz��k��b�O^�O
��|"���?��"
ٹ�K=?|pa� P	 ��U��?A+Ob��'���' 2P>��󠖳([���F�K�Z���9?�"]���I��('��b�6�)U�R
%C(��P��%�<�;�m	��2aA1��R~�O)rq�	�%�'����
�+7����j�o��;2�'���'�����O��Ɋ�M+��'7�x���)� x��hL�<Y*OD�o�V�,��I�(��0!X`�J�"�9�4RcΆzy��ɡ3S�����E,�d/HqybG�
Ov�:�Fҳ8�l|���4�y�T�(�I��D����,�	�0�O��y�c�+;Ζ�8��1������>i��?I����<�b��y��.j\�5{�� 1E3�=@��"���'�ɧ�O]��IQ�i��� �����:U̜H�#H���^��v=O^���l��?���%�$�<�'�?y����v���*�X�,�����^��?1���?������h}b�'|��'����`�e]� 邮��U���2��R}��'��O"|���Z0t��ܡ|�t�2����P��o�:}#5EV��n�bğиr�G .u��V�F$c#�T�t��ߟ`�	ܟ �����D�t�'���D�N�f!��OY�.w�\bu�'� ��?���0ɛ��4�l��Ծ#�h��@�E�"|T���9O����OH��Š6-4?)�&����)^*b���V%�#_��A�D�zL��J>q.O��O<���Ob���O��S��X������5h�!򓌾<	Q������(�	~�s���5���VE��&@��~��5B	1��$�O���6��)0d����V[{lٲ!�>$L`	y5�no��-}|����'���&���'�x퉂GQ8 �53�R01��'4��'������V�X�O��s>�ˆO�gW���Fh��Ao�����?�3^������	�B1V��qIF�C�����I6�8;���Ӧ	�'.&�1���?u�}�������3��x�\��
�H	�U͓�?a���?a���?���ON���p,�"B'���-�FX���'���'�����æ�&��K`հ6�vDq���s¬H��(���H�'��ta��iD���T6V��-N�N��- P�(:��*Y,��	�P�Oy2�'G��'mr!۽Sb&h�͙
����N d�'��I4��D�O����O��'cg�ͣ@�$GZ�(x�l�2Eh!�'t���?1���S��-	K_�+�ڙqx��)��TFݒȰ4�N5�6��擏:v�$/�ɮ�ĐH���3|���+����Gy��D�O����Oj��<ɳ�i����W�B�쑪Ǌ+xUb�'�r�']N7M$��)���O�I�R�$~i�ԏM"�(uE�<yu�T!�M��O"U�A��
 ��<�Fo��w^ڵ
*�PInH��l�*]��8 �$_�n��Щ�e�?�r�J�\v�J�(�Lq�QCo�$I����gjѫ��y��៘.���
�`�_䔽�
��T'a}�J_����t*�';�f�f�?|���ī�C�Z鄄GB^�Q�Ď�W��P��(�-'���de�+T��Ud�6J߮���C#��Y*�ᅲr)���l��5'�@�1J��1���a� ^��8�2A)����Q₼f�xBe,�u>��3�e�f;�Ѥ�] R�Nh�I��M���?��?	dV��'[�A����.IZP6`1�SG@7��ͺ�(����~��s�X�B}@�i��[�~.-�Ÿi�'HR�'��	�0�	ɟ��) �p#BZ��������_�Z�m�[�ɧ;U���K|j���?Y�5ܘmI`$*P*�k��]Sjn$�#�ilB�'���ߟ��I՟8&���hm��̫Sp�� Ƌ(=q��-@���K>y���?!������IoJ�`�ͫQ�bE2m�$ú7�I}bX��	a�I���	�]��Tx�#�k��(5-%X�ޜa��	E�	韬��ן'?��'?���Kd��%*|� �J'v6h`l�������h&�����<9��IL?��nr ���@'cY�#��C}�'L2�'L��y�OH"��3R�Z|��jK/V�X���KG�6m�O�O��D�O�e9aN�O��'�bD��-�"p��+�G-	R�`˹��I󟼗'�"]>��	쟠�I<H�.�SቮL_ryy�jô���0H<���?',�������{�6�P��ƞd2ZX����7�f_���Iß,����<�Iޟ���5��@'d���E�,���h��M���?)���!����O��|� �ʸta]�1Ɇ�c*e0ٴ�?i��i���'��'��듵�ĕ���p��f�	^"���C��8@�l�0����I^��Y�'�?9����~���$�1*hu:����j����'2�'����>�(O��ħ�@E�8}�B��D�f�v�J�&�ɝw��'�P��ȟ��I�>�\lE�[W�|���ܛq�d���4�?���+s��]yB�'tɧ5�%�%�Ĥ[�l��1�����섺����[� �O����OP�$$�(�N���B���.<^aQ"���M3�Y���'�R�|��'��� �X��1�*5��$x��� /��|��'�'��OǊ�,}�6�W%� 6h�8'��9�`6�<������?����V���'8��e�E�y`�r�δ-0Y�O^���O���G�S��ħ �����Ɨ4,8̋PHPk���B��i���|�^���ϟ짟����g�J� x{(��/�T[�i���'N�ʟ��K|���?��
@r�D&	�|,��	���@��'�ȕ'OR�'b��yZwP~|�6͈.8��a�B`�#��h��4��$�Om���i�O2�d�Q~2��"7bj	���1�P��P���MS,O����O��&>'?7��pl\LxC�	-:ɰ6���w��	Ο��	��I�䔧�	�G-�,(��W4RaQp ��^.��'@\l���Sצ5��)T%~"��2ǏW2k����imb�'�b�'��)�N�!AJ��&�:����^	q1d�QDn���O6��~Z���~��F��}�F�N�?2��%��8�M����?�/O��O^�O�@XāP��"Q��#v�4�:��|�ɥ9�b���iy��O� � �2@�*7�2D�#gL*QƜ��T�iU�	ڟ���w��?��'n�,���f�ԩp��!/m�a�4:�ܤ�<Y���d�<��O5Fb��0sy����ˀ-I�ߴ�?�����'��V���{ӊ��Ӎ��L��n�,mY|��`�x��'��ly�[>	�ɮ^������ P��O	<��e�ش��'XBZ����$0�dÍ}Wl�3����v�"�ҳ|���'�Q������'�?���C�	V�/��	�g��/f���c����Ŗ'-��'v��'���yZc6��HA�O�2GjԈ���r��Xx�O�ʓ�?����?���?)O�Δ{@h�!�,�%8�dR�Ȫu�v�'��I���"<%>}�W`�;	D���^�Jq�AdO}��DVȦy�	ܟ���џhI<�'�� RaO�@֙R0D\㶍�E�i�B�''��'��J��'�[mr�yQ��9+NT4YU�?|7M�O���O
��Zo�)��'^0q���\���b .J�PF�U�ݴ�?�H>�[?�I�h�I�t�&��6 P	C=���C����M{��?a�P���'U�Q���i�Y
��H3-� Y����0�ܴ(S�n����S�$�<���?!����$��S��F�L�`C+��{a����i�L�����O:˓�?����?A֦�H�ـBc_�	|6-
6Οcy�X��?���?����?�J~r��i�
�ӆ��J�^dI�'Jq�j�.n���d�O4�$�O��$�<���\9��ϧ��Rv$��R�Z5�p��w���P[�P�Iɟ�IFy��'��꧈?Yv�e)8g��2�dځ�Q!vX��4�?)(O��O��dW�v�0}�
w����_��>E���M���?a)O���E�D�'��' (TbT�X%�X��t�_�P��2�J�>	��?��;����9OX���g��-Bv)�T[�} Q�P�o��6M�<��:����'�b�'Ҩ�>��-�L)��KE��k���&N.m�ԟ��� fE����9O��>i9d�W�V��YH���7��t�0�g��$���M�	���	۟�ʯO�˓��T�CP<6��)�)�9N}:|��i��T��O<���O�r����l��o��H��̥e��7�O����Oz�d�~}�_�p�	P?�2��#��@��S?o��R�m����%���#�p���?����?��oY	2#��2��E P\ċV)Ÿ"��V�'��o�>i*O��d�<a��KP&DX��<2Q�Gx�r )�C}��y�S�l����T�}� ��AI��Č�?.be��æ���Onʓ�?�/Ol��O��D�v�>�:���7G���9�B�۶�#�d�O:���O蒟f��'Y6��*fe�1���Z��F�tf`�o�syB�''�����I��d�o�֘�Gf��
�� #�T��&a;�6��O0�d�O��D�<	�6���̟�� 0ഠ��( ,Yp���
,6-�OD��?���?��G�<)����F�ЍU�̽��-�T��	�Ύ���������'O�~���?y��K7����ꑘU�1Q�D2=d��vT�`���<�I(��	ǟ$�'���ǜ����� ��V� �`�	F 39��'YB�'�>7��O0�$�O��������ݨ
"�9j�EP�5ұ*��iE�'��^��'��i>A��� XVHÏ'iL�)��ݥE�(���i��ImӬ��Oh�$�O����O����O���	�;F�!k�IĐ~��m��LT���a���{y�^��3?�'�?�AC/DDYk�+'"�W�;E雖�'b�'�"G�>i(O��$��T�s(��Rd�<�p�;-X�� �>1+O�d�ם�����˟ʂ�Oi��q�h�%Gl�����L��M����?q�X��'~�W��i�y�7��3^�}Ƀ��H�R��u��>��R�<y��?����?9�����$2�)�����,�2r��2�i>듿��O��?!���?٣��
��hՆ��PĐ���,��l����'���'���'��i>�ȝO'��*�-c<�XJd��:e��	޴����O���?i��?�vX�<�U�(Z*YhP��&T��PjBfό#��	͟|��؟�	T�$tӘ���O�h9�������G(	�O�R�Fj�즱�I֟ ��Uy��'�F9ۖT����a꫆�7���)݂%.A�i��'"��'�ge�^�$�O�D�O���T`�F��WBy�bѦ%��Sy�'U|���T�����ܴ+��лw���<�D�ς(�hn^y"�'�6��O����O$�$�B}Zw*�,7��-6x��օ�(�%��4�?���Xn����?A*O`�>qh��o��� `��
�j�"qz�6�$ۦ��I��0��ޟ�S�� ���h0i�o�X-"6Y�5��TX�B��MD'�2�����y��'��`�	!C���ɥ����,�mvӰ���O���OF��'��I����R�Qq@��V�����Yk2q�'��	$?U���|����?��|T~�����&�
�{0a[�N{N��i1��'� 6��O��d�O��D���O�P�o<7�����Ki�*=�X� x��/?��?����?�.O���q�ҹX3*H�'�
����)e��A�>9*OV��<1��?Q�y���OY�,QDE���"{�Y�F�<�*O����O��D+�	��|� &ױw�|��V*�Q˶%̦Ŗ'�B\�����@�Ɉ�
�ɬcK���%��8�*yjD	�\�½c�4�?���?����4��8�O���7� �]"�&^<L�P�;����`O=!�iE�X� �I����8P����~���X"6Y�%�G�7!R0 "ᐼ�M����?+O���l���'��'�b�2.h�N��uK��2'�m��>���?1��)�� ���9Ov�S/u�TI�e�*N�pF��Om.7-�O����O�oϟ��	֟0�	�?���U�0s�W�hn�q+4Ia�0c�Op�D��2��$�O���|�N?�ɰ�
yLb�-��?ުT׋h��������������܉M<�������X#e^�r��Ѹ_Sq�i�����'M�'3�f�d����"=�HIc2�� �M���3�M;���?q���?�1���OL�Ij�^]ʐm_2!"�����E~c�X�v�:�	ğ�����zU�;iݢ�����I�� ����Ms���?����O��OkL�~� S7H�t�fQ�Ї\�k��	�Yl�	Fy��'J��'�W:xU���=���)��6�X�m���?i���䓱?a�e(����*a��e��L@r0�#3�D�<.O
�$�O4�$8���|���GPm<�
���}9K@g}��'E�Y����Ɵ�Ɂ8�z�Ɏ ���W��WX��1ϖ�o���ON�D�OJ�$�d��%�ħq���±$��4Y�I���:@z@�iY��|��'X�i�o�"�>Y�5D�-9���:m��}1���ۦa�	����'B�:���O����5qCdl2-\�h}�Yp�I*{�N�&���ӟ8��!�̟�'���'o��m	�ǣc|���n=L:�nyy��'�^6mJh���'�b�%?��0��薫B�'�hׁO�%�	��`K�ҟ�%�b?5*�a��#`L�y�b�/3�D��i�4��X������<��ޟ�0M<Q��S�tϚ�'�K%�^�8FL�r�i~��3�'��'���$׽c�����4t�4)��(h��!n���������	���'��Od!�Q�F/V�6x�G�ͽj$8h8�i=�'*��r��O��'�����.h�E�˗4�d���6T6��OH��]�Iş�	w�i��q�"�.����hM
M��@����>��(ѵ�?y,O^�d�O���1�td()r�I����=e�|Ec��.�M��x2�'���|"�'��/\���� ��7 J�H�#(������'��I��I��&?�I�O�J���u>]�����B�ȮOv���O��Ot���O��`-���x& \�u,i3��T :�9�>���?��p7�OEJ��s#(֐! Ġ�k�	��	���Ʀ�G{_�8�Iw��E��,huHZInlE��ΐp�ZH�q��R����4��S�(��7/���@����	YO(ə�Td�
���+�2���ro�^�n�+��z}�p�����H6o���`(�{P	��i�r����a�*����N�$l�M�����r�`��ǅ�Bx�a��Wrt ���%�Ȉ�ć7d1a1�AV��J㌋VPD!0��2.��DAuCٙ^�����&��xА|C�jIZ+��I�H� oCZ�)F��8:����AܗB��\P^��d��BB�p�1�@-\T�Ղ���T�a6ĝ�� �ʡg�]m@p�F��@B�6��O��$�O��)�ͨ��Y�M���Q��}m\u��Ğ
�\�uo6L ��G�g��xi��&B�f�6y
O� �j�z�-�z�I�W���W��|���b7��%ʵE֊��D��S(R��+i�O�)&ړ�� ƺ5,�bg� �a����z �I�I�9dԨ�i"��I�6�'7V"=�O��Ƀe�>e�v�_����C`E�S̨p� ��M���?!����Ol��|>�3�HA>V1��tMV�4V"��"��0I�X�	Z��q(��Ux�kU�Y�ML$��X"8�$x��וY3H���#�_3F�C�[x����C֋z�0�$�3F��%�O$���ON�=!��8pN�lA�n!�6����y� �;3
4i�Ui�'c�-X�W��'������":%�']R痯�Z9P G�$DD#�
9!rZ����ͧ~a�l����"�y�W�O
� &�
EAĩ�f��&"��Ӗ�'{��XTė)��l��h��t��F�)~�0!v/;�LCF�3O�=�t�'F^�"��ånJ*��g�fv�6�/�IB��0�p'�)L �J�@7&U݁4
Of�o�:�R�Y2��(�1p oʌX��_yR`Љ2bꓮ?yN~�����xҲ&B0�$۴$ȑu>��;��?���,y$^�)��/3�^�S��^>����]�u8$�W-�-9�lzCk9}�JW�5������!D�ڣ~�"�S�e�J!�`E��:���T�$JH$�'o�>m���B?PwJ�?��ĩ�9ئC䉪:Od�� &R6�$��b�8����Ċy�'��0{S	Fx�R�*�(q��	%H�>����?q��V�|����?q���d�#Re E��MG 5fH���"C:�#�"ޯ��D�4=��#�|RhR�L���ZUو�z0��B	 2��塖*Qv}�fT�#%��}&��I���m�5�g��	����џ$�'"ɫ��|���(^Hn�k��Õh�L�@��s=!��N�EB$HÕe�8�>���X0/�	��HO��wy
� �l���Y�����mM$���
��=�qo�����͟4�'�"�'V���SM��pH��y�ʱ���ʩf@���Љ,�����X)Ԭ;�d7Z��Uؐ�̪W�t��v��C�����1�az"��!j��vj�f�j���l��5�(}#���?���i�V�H�	ZyRV���G�L>.�rX��e�$�@U��>D�H�0����4�&�Sw�.�Pt̓�M�ıi��I�|�n��p�I������BWX@ʰ�@�e
�y�	my�'I�?����������O�u9�'\� ��A�w䆪!2hP`e�'��T�E� �bX�'JL�S��A�R��a�Q�B��IǓ�J��	ɟ��	ҟ�8a�N�`���3v�B�(3j�(�My��'I�O>�/N3�@Ia�.yX����;0!�ā��%�W ĉX("�3���6�6�x��򟘔'��4j��'��'��s��ɠ/�J�����2R���w��X���O�d�9ow�d>�|�'�vUj�B.W1j��R4(��O�(�k4�S�'d�|�إ���0 �b�<i����O�e@&�'���'�2�iI%D�Z� ��D.�����r�yB�'��y��!��M+Ӈ����T"�0<)`�	0Uٴ�A��ǰ5�D�2$�XS�[�O���O<y��1�����O��ı<Q5),m�JR�M@�`�d؛��܂�`�OPi�*��1��'ҜM;ahD�7��t`.�"r^,�#U*T���q�X��v��|Ҭɲ)ܺ@Srf~�0�`���q�B�'e2)fk��,O��W�C���6�\���I���)�@C�	|��c��'�ic����6��[���h�O���S���D�4=��
�H�Qk�m�$���M���?Y����D�O4�du>}��ƴW���[�F�6����G �5ФB�	%`��d�u����]3���hn�i��&�x�u,� ZW�����s�͉V&V	I����;�ObIҭI�U(�lf�ޞ<\y8�"O>6��z.�+�,Լ��	&��C�bx���Ұiw��'p�P��<�^�� l<#/�$���'�����I�|
4���('����1,��è�.d��E��:O>�y�D���2d	�s� lׇ.��x2�ː�?�J>�	>*�����ʛ67]�|딎v�<q�$
h���-�t�L�!�b�o<��ioL�`DJ�:1"E��L�����yBg̺G����?�K~���S�x�i�� l�}[��Z�v������?��#�*�v��I a�@����Ķ��|j���,��)*%���@%�1�O�D� #s�9K7��3=8"-#A�R���P�qǢA�'�f9�b���#��eQ6�>ID�O���7ڧ�?�`�
ȺL�2cOZe�T�sG�R�<y&/��\.���a͓Ŝ�:��V�����٭J��n�<@*�)ʛ=��n�ҟ ��֟g k>�Iʟ���Ty��:F�� S�l��	!VR(�1OX���':ڑ�l�I�Dd���t�z袏{�#Y&��<�	B�v�!%�V�)Z
E<�?q�O�5R�����?����?Q�)�%Q���f�X/|'� 6��x"mԒU̜�1�ON*�teH��H9���@c�����'/�Ɏi�>��T����^ j�Aԫ&��12��*�M����?�����O|�$r>U�ЕU�NAxgA
V5��Щ��
��X$�Yx����T�{?��Y�LD*w�)c�/�/}?���ևEx����'K8���zbϓ�	r��uѝL�^���O��D�O��?!����Qe�iP�#*�4 ��Ӣ�y��@o��0�CO]zm�F��'��6�O��vdu5T?��I�V-�=�6����Ѻ�צ5kĩ��GyR�'��<��CJ�l�"E����B?�cᗞ_ �b�oX>6�r���Oq8�@I���V�@�`O��~rى6�Bj��E)q#�mI��ڣ�p<1��ҟD�	ByrH�/A1�ƪ�<\������Ԙ'��{��CO�~�s�V�M
��1*��x|�ԝ03@�M�b��dB#t���9Oxʓl/���3�i���'�O���#o���Iv)�!Ulac`.D&W1��'���'�1O�3?��-N�s���si��I�ެ�]�	3���?�Km+w�T�qo �EN4ҁ�-}rc� �?Y�y���� .j��3��y;�����^&�y��/G��,����tH��"��C0�0<s�ɲze�-a��D�Y�T�7�B�)� h���F5n1)�҄s��xd"O�=�e[�1�F #�$�r�rK�"O���5&١J	Fܲ�@IhZ(�Y�"O��ag��t�d����.k��(�"O���).X0Ѻ��Y�:d	�"O��Y��
i��84�� �2��a*O ؠ�+A'���$��:GX*��'�Ь�u∍z����S�T�)�T-p�'�y����,oph����o��=��''n��f���Z�,3�e��J�	�'�8��J<��c�b�Y��'�zY���2��'p���'tB`�@�,:���S���i�
��
�'wb�R �,x8�W�Kf�
 ��'���Č�?[D�{w�P�d�:�	�'��M���(�P��w�Z�v�"�'5p�z�яu��U�'B�JF��z�'N"9��_� ؙ�Vìz���'�$�'e �E�\�(�J�wuB��'�n	�w	C^%��`ɾu�ͻ	�'*��'ʐ�7Z���ۂ�A�'R��Q���� ��2����'�&!�CG�6F���'�]�M� tz�'���5唫V�z��4>�qb�'�j<���j7񡢄K
ir��'5D=ɇ��u�b锂s��q�ʓ7��ʂ�H	wK�����|6��ȓ7 �퀑��& �gz�`{�'`$��!�~�(PkA�8kIx���'���� S�bj�{ �5�����'<H!���4�,�ワa�B���'JBXK�n�R.�ٙ��I�z��'�iQ ���,)b�L?��|r�'��͡���� P�L�	�&tZ�'Nf��*�+����Sm
6vf%�
�'�޹v�Ho҄Z&DV�zD�Di
�'GzZt�Z��D��"Mp[��+	�'����GB�pU<<b�	I�aT���'}ĸ��iK0����?l�]¡"Oh�2��"w2a��ֶn����g"O�1c�%: 0q&DΚ4�I�"O(����C�[kR �M��t�&x��"O�]�1M�$뢀`V�;F���g"OZ����0!��KrLE3�N]�U"ORE@�@	:J0�8��m�\ĸg"OΌs��r�$�P�������c�"O��Z�"���	adLZ�d\0�q"O�t���1.�B�2��D�7e0�8�'1δ��ⵟ�bQ�:�1�%d����Zs�#D�X��kN��"hkRi?82�80�!7�7by�"k/�"�J�1aaH�Z$R]�!h�C�Ly�ȓx�ԁ;�� � \Sƫ��=�¹��I�w�)�=E���)��&�׹8&p*���2ys�(�ȓ6P0i�'ҋ)e~�1(]+h0X�u�Nlis�1�O��agLYj���� dyn��e�'���zQ�i���U�P�T��JߛN^�� ��'D�(aF�+Vb9	��݄K>�0(c;D�|��(��3(��	-;-qd�U�:D�� �O�1�4��'Ț/-<���7D�T�q����Pjf˙�\Ys7D�d��9��0,Z2P��dh�l/D���.*[	� 5J����۠�-D�8!���W�����c���#�O,D� (gnHY/�U�@c�I��,�q�%D�� ��8���I�;�8��0�'��RRP��A���)��4�̯hp��h$D���`�N�bq�VK�q��!�`	8�$�,  )1�'K��eW���S��)VI���݆�&��%��`X$n �e�
�y�b�L����"~�n������KL{  :��Z�T��5�ȓapF5r늫,"�\W�I�M0�g0���&�;�O���.�)$޲8�QO�6VP�+��'"v����OA?ye	-{��bԨ�?�Pa���\�<�E���^(IAծ�<Wr�=� �X�'��u��NK�OAH�h�9qj���B��5
��8	�'��ju	Q�BvTx)��&�b��u�[���=E��'�I:G�W��]�VlJ3s�9�'$���M�S*D�y�,�=�(%�M(~]��9�JT�wH2y�׆B2Pay"��'>q�혃e�$W�laK%	_��0<��g�<l$�`bK
	x��V��=?�p�q�Y�=�$�0�N¿kv���k9�t����$���(E2_�hS�J;?�')@� 6Ӣ���N46�1��ן�>)��UF�A�%�m����8D��� ��?z2ܐ��ʕ��p1�BU�Op���#�	-\�j�@b>Yʔ�>)Ba�qX1�ł�	t��`�͔k��|1��1��h���N�yy�tʄ���-�T�4D�ՙ�O\��H�؆AŠ�p<��a�Qi� �w-J6?L�t@Q��U�'׼y��HD�p��|���{�P���'��㥥��t���
�cL$P�F�P(<�Ak�3?s��ga�*�:���I[��8�7�	>�f�P������Ec&?�|r�eP�}��r�Z��dh�eЩ�yb͗�$��5���-96�a�X>GV|�J��H�kX���(cG�8�O؊��kSl�$��s���HBm�2�Iᑦ�X�~ڌB�����j�)��}�� sQv�xC��'x(�0��7�z2m��w�.}��I6=�E�u�A4VN�d�B�>I��?�M�-GQX8c�m�3x$��S�]/*����:w�>t�pm&h�4$��|(<Q7cN��@E������4��@]V}"Zl����IDj���5/['�~���#��h^����3:7�t�I�y"��B$�\"'A��u���p!�� O�#@*�2���+y�y��ęZ�	i�$��!�1;�EX L?�uYSj��f�b.ЮG�6ՋЩ7^��K�֐��;�dC�H*q�IߚDn�5�O��p<�'K�M|F��d.ˁ(c�e���GO�'�6��B��l���ۓi��^������#?�̰q�(Y6RUZ1�a_,Z<��'G♋#�^	�^��D6|�Y�O���3�,��=���X3�$�)E+`�q���(7��?ڬa�];3����"O���ɚ�v���w�ȯ`I�\k�����h�b�09�7-��+�2�>�J�Hhᦞ�Nձ2�z>4u�!��rW�\ v��xK�D���P���2��bD��$h@�R��.e��+�a?=r�Ɗ#mԂ���b�3Q� @�ቃu�h���U���p��_�AC�%���S�΄R��u1�_���$�&( QC�h�-T��0�0�ـT���(��cPi��A)ʤ��*���ɕ��2��'A��|�F��u%���!�d�*4@Z�'�~�I��JײpNvЪF����c�i�Z�X����''���T-I�	}D�ib��ڎoFnq��OT,K�aŦh��!(��Jx����aU�Vm�J�@a���~bc��Lq���dZ�DF��H�(ԕ:iч[Tax2��e�zD���>ݠ6�S!b��a9�fW�HA0�P�U/c^��'m���C�M�XD�6�'t�A���C�!д�[DHX�O�<A�aQ�d��������xJi�?OJUpPĬp$�`!kʔ~M�쩳�$4���P���֬WD�����1+L �R��|��<�c���w��bf�xT��A�V��[�'c����
�G�,x�S�D����M#PW����*���~Zw��yPÒ>�Z�1�O:�� �8�����G�z�~u{P�'�p?�<*W!��C�5�	Ô9;��HG#�<<�t�r�O���eUZ1��S��ӵ��O��ABj�9r 4���-��@�"Q(�|ˇ�Ĳg��`\5�0� �d�P�Q�{�2�"G�
��n�@�,��?9���=���cE�C4`�Ƞhc�ܮCY�	ӷ��.eA��v6���',(}�T>�]�&�:���.Y���١b7Rh�B�C��1��͌u����'�Ȕ���2�@+?9�O��-�j�'���s�掵3=�.O�3�N�NحzC�ձ/�rl2��'-�|��k�����Y� ,I5� 7�x������/B���4�
q!u��I����*Ĺ*�,�?�4D�y��e ��ј������ܓ�h^��]���[�,\�0L>�&Y4��q��-"���d� ��`�M�)��?9�JK��9��A�q��E �#,�U���'�D"��ȼ� c(cG
�2,��*�N�J��Z�'s@9V G�!�\U�s
F�H$�A�ݴ{P���SƘ���@b�iV-7 �Fyr	Ќ;Ю��WΈ�F�A`�aF���>�ҌjAa�_\��C�ȁI��I+J���&�P�M��n��F"=ᥪ^�P��+m�:���4�(�RQ'_	Ë��8@x�O�*x�?1և�<fB pH�S$?���!"��#���a"���>sCޟ~U�����
F(; c��q�����en�ދ>{Z8��j�=To� d�dcQ���3������A��� �.pB2Ϋ~��A��a�y����W�'�����	�I�C�/Z��x�z�BK~����oV���ȕ�wш��#�2���F�C�����,>l�z�N�w+hd{�B؛(D�OPijqI�MaaJ����$ڂ�!@�O�i� C�_�4%��!Z(4����=<���%Z	g�\1��_���ȃ)ݢ�r&��2wc���˓b�z%z6R�D�$E:��R2=���)�G�'� $J�C"O���æɍ %��
)����E`Z\��Q`H<Q��ھ[�t��"B�5�x������O~T�O�H����A�F���n8F7q��ׁ�"�r@��.F��}B��Vրap��l
)i�/�26��-��#�1R󤠟���dI^A���փJ�K�ў,�0��
� �2�ȑ��ŢW$9�O�%YTi\#aφ jsOY�n$lU1�썰h�L��d�vw��
���-�5�A�j� �Ʃ3"E~f��9\	@QK�'	�N��O�Ȱ��ϕBe�4)�i��R�\e@	�'y���%�z�CA��5qfmb�O��9�l*z��7c������Q̎&���E�af�HZ�"O��۠Ě�__��x��@�Z�j�PE�M��I7C5jH�1Jy�3�	�I`�<K!�$^>\|��E�I��C�>uR�16��6��Ij"7!QrB�ɍA��鱀�8
������nw�B�	&vR���G�E����` �ͮ
Z�B�I�?vP����ӌ+��u���'�FC�ɵ_z ��ԈQ�m���BrJN�%T8C��\����a�<8v�"`̟�*��C�ɧ �a��U!it�@䑾q��C�ɫ.�6�Oɭ)bM2�OQkʹC�I	>^l��,��a�Bf�7�C�	nAn��G� 0@����ZC�	AF�=���#I�,�?� E�g�<��I�,'}h}�v!�r��ȉ�i|�<Ye��<l��,)#�C�B��Z$�}�<���C�`�W���9���B�I�Yκa2R��~�v�e���C䉨.��\����\��Ac E�!9`C�[���KF�R�:��HB�Sf�>C�I����BsK�"ʎ!'��8� C䉽�Y2�K�"zvn �9c�,B�I�M���7iߵDNm�ׄ��X��C�-\R:����Ӏ9�����M+v��C�*:����w�3]� [�ʃ)D�C�Ƀ�ʕ �׊t���rb�9U��B�BS>DZbMI�������0&��B�ɢ 8[cJA
�J0c׫]�T@bB�9����<� 2�XzC�I|� eeY9O��A�D6RC�I�%?�`v��q2���n"r�`B�ɀO�6�@�x�کRP��p��B�	�x^&���V)p@�5���(B�	����˄�čzA$A�RA:<�C䉏X*je�5bb��3c�,7Q(ن�H[��!hI�b�N����ܑS�؆ȓ}���a�E.J�[���I%I�<�3�zΜ<y��$�tT�s�Fh�<cś�HZ�{#�N}VDbB��Y�<� ٙ�g	����),z�-q"O�j�������b�Ãg�\;"O�DRlM�vxvQX�F҇`亼��"O������gt�Y1E��(mq"O0��ҮAw�"��k�R�
%"O^�0G�RITɪ�C"u�D��"O�8b�A��)ބ��a�pn��k%"O��;`ƏDl�x[t@��*_���r"O����#��pH E"	�,Fx��"O�TB5nۖl�f�!`�"6�l�%"O<�uG͘2��gE�o� k�"Od��G�)��TC�!�kR)qA"O��j���"U��!��U&"�&��@"Ol��P��9 C"t)kV:s��K�"O�]2�e�6b��L���6sn�e�"O��3��/�l��(�	=�,���"O@<c�J ~�6��w�.�T a"O =A�e0lT����n�^�x�"O����"��j��T����%7p�´"O� �3��)CY�����<>`.tӡ"O���KЙk$8HU�
_Y	c"Or4������je�V�t���"O�顴G�8@DY�f�WW���q�"O��#�n	c�:�s�!*� ���'D�+4�ߔ'L�%IE%<x��'��X�rf�PT��U-H�/�%�'p��(c�A��*/��3
�'f:���_E�cV[�~I�q[�'3� pg��h��U�v�1e�N���'��!tN\f�s$�*},�	�'����PiT7��L�E��Q����'���sk �BQ�5eЈ^���Q�'���zUڀ9-H�/]�T��m �'h���W�����ᓑM_�~PRh��'���L�{�pA��c��
�С�'��]���XU��	!�M��q*�'jR�z��ѻu����'�V�⠀�'�<�/N�zUCG�)v����'Z����	�o�2��-po\�9�'�X��넾��(�k�o�*�:�'<6$����t�&Y�#c�r$L���'nK��!�2���"U��0�S�c�n�<��bUXJ��>X��MC� j�<A� f����f(� ,c�U�Ld�<�#��95@B�Y�����(��ǛK�<!a�%m�^��g�o�BD��H�<#�
�}�z�ie�_��VQ�Q�k�<��3ǖ��נ�*��Itg�k�<�Rf_.a`� �>8�E��{�<����m��	��.���L�<� Ș7����&&Ke걚�N�E�<)t �Bg�8j�
��r�*:�&���|�l�t�bd�h��D�A�%LM�ȓl[}�oƋ[w05���D�-h
F}���81�|(I%��l�����ì4c8B�	�|(�S3�q�682Q��C��`]"�ǿj��,���UG��C�	e�e 0��(��j��}�C�I11z���V�c�܅��+�v��C�ɻ	V�0�ŗ(�������2��B�	�-�E������� ֩Ʒe�B�	0�%�B	=Y>��h�=;u$C�	�DFdA�g�r݂%��g�
S'�C�I�g���2MЁv�@�i ��&A�C�)� �hqe AJf� ��	8+�~�Z�"O���6i�]����qIA#0��y�"OnX8�	8��"JOCL!q�"O�`Y��Hjxp��H�y�E��"O�UQ!����Z��'��d�(�V[��D{��)��3�ex�J�lsΉi��2�!�DǼl�2A��+T�A��2;�!򤔄.qİ)T&ڍAZNa{VH��J�!��9H�9���CcxР�U�V	J1!�Ě�d�~���X�����Fp�!�$H�  �a#J&��J"n{!�$�[���Q�.,�=(F���!�d�;�t%uF�%�b�#7/��@�f4G{���'̴�������m_�8�@�Q�.D� Ȧ��`R���� .p�TM+D�ࡁG
�$&<3⩞8I��=��+D�̰0�����@�0��e	r�@�`'D�x�4c�&e!މ��� D(f�lG�<�g �m<�ź��T�Bv�г��}X�<�O��9"��:SԢ��B&ȶk���*%"O�0��gA@��Z>o-T�3�"OXxp��ۇj.f"5�'����"O �0���8xJ5�W�G�0�A�2"OfẶ �!�.Qk��1#s� T"OP��I�%� �{���WI���"O�mX��\�|0X��I��|�2"O@U���0R��*�$L�"Onɂ%�a$�ջ�ʏ�6��z@"O����?sX*踤
̾Y����e"O2�Z�@
#%��rԩLTu�yA$"O�0+�dW�a��lh���X��"Oz��F㝞o׶�Z�ꏢ]���(�"O+o��]碡ځb���b9�%Ch�<�$#�	@����h�0̞�@u.K�<��/�xք��&� ��F�G�<��̓�t#�=⣇�C�$�i�Z�<�2m�4� ]��f� )�c��{}B�
_��H�0��A��|@r���c����"Ot��Fy��=}��A"O���������Q���8:z���"O@ًîe	��Jb���~I¡�t"Od1�'F�P�T�a����p1����"O�Y�� ɚjrvx"��-a��{�"O�	4)K&.�~���E�C&��"O(���
kb�!��2�"Ou@�A� J�Э@�fD	���1"O�	��d?I��=Zg&��ml<r&"O<9 6��60W�Ɉ��΄t>�Y�"O`|�#�"A~��ŉ��6�TA�%�Im����D?ڦ!q�
<4�yI�+u�!�E�d���H $ �3�B��!�d��]���(�n�x��pQ#�L�!�d	-rU	p��	��պb�K&!�dҧ|�pX2���`����%��i
!�D�\�A��c�����g�	X�!��f4��[���>o�֕XvDɕp!�� >b ���%�`:6�b%d�X�!�fa@�k7��3&�����!��ט��B*�6L����F�[#L�!�Ē�I�.�j�lϖU���a�7H�!�DY�n����P�$�Tpb�oԅ{!�J80 ���p-�(�u� �D�ȓ3�f�8�힓X8�z�"Ӎ rņ�|�I�^6TH�8u��KO���S�? �՚G�2��� �|��eɓ"O�U��o]�""�!�di��LYd"O�mruN���-��(�!{�.���"O�!��݄0/
�8�K�n`B�:�"O(9���x]ʀ�E�!I��S"OhA{���$U>]2r��wGjĪ�"OP��$Fj��P�^�tȈ��"Ov]�b� �>�` B-R�J��56S��
�k�
� D���R�i�F�&:�܀���}pr�
?�:�R�Ӛ�I��"O����#׋�\��b�t
҂��#�S��-H�|��r�ۥ;���to��)�!��zF����W!��a%��{���6�S�O��1�i�!��
���	8�.���'5������+�z�0Í��2J����t'���of�'~%1D�N���0�[5T�r���'D&�i�a/}_4 )c	�h@��'� aBM?Q�( �g�	�8�'7VT�G�E�3}�! �-���t��'�b-a4!ŷ3�" �1y~|���'T��vF�	^�@ĚҪ ���	�'��t)�NA�	�~ �!�Q+��x
�'�81i��p�ы�
 �P�'y�hE.	*d���`h�z�D�
�']蔰���T��`�����l�<�
�'<0��祜a#��!)ܝ/?6L@
�'�N�Y4劢+{8!��*
'4b�s	�'liB*5���:�޺%�]��'O<T��,��b�����$�r�
�'NЈ�D�SÐ����[�+��+	�'l�[����g0*0�䯈�'����	�'�,TA�鏍Qe2��S�E7�DL	�'�R�+B�E k����aä	 ��:�'1�}1��}+VX+r�X�K>nh��'+l\�F����}��k %S����
�'FLha*�4����WIk�P�	�']���CI�$��+�i��!��'�2 �ɟ1��獔�d�t@��'�!Äc��2��	�� ��(�'�4�RPB�3}V!zu�ҁ,��'�H#�
�]V�����ӆr^��k�'Lr�&�l����]����'�L�C஁�pC�Y���"?;�`�'T|@[���"_��QI�$Q1� x+�'N�1��S<��r��,����'�]�`�� f��x��
B16k���'K�I��"��RK�)>0N��' �C�k&��@���?EO�1S�'e�	�eaA��%�M�'my�D.Mq�<��H�%�y�Š\����a��o�<���$S'@q�%��T�ȥE�@�<DnA�8���ʢ�Y���[x�<Ѧ�U�lܹy�NU�6� UHy�<A�oW�9,�r�QwP$[�jQt�<���Z!*\y��IO�'�,�R3�H�<ц�U�?�n����&Y]��XB�<!���-��5R/�<D�49���V�<	��Ղ0�1��-��D�V`���k�<�ᓅT��iV#�1�rͩL�L�<A�� dl�GgǊ�d�y���K�<Q@��n�,iG��?����t��K�<�q"M
UW � �,�-I�L�T�D�<���E�
�QJæA�.X�gkRZ�<�%��3���Z����^�$ J�ϏX�<� P��FB[�f�
�!��I/d2]�%"Ov�zD��U0vb��
�\\.���"O�(b����T���(�4IV �"O�1B苶'ʤ=����8E����"O
����P�͠���yC��xc"O��+ &�W��PsU�E8�=´"O
-���aEH�;� 2��8[�!�ds� �"�d���3ȑw�!���d��BE0k� Š�j��"O���Ҏ��{]�ಗǀ�e�p��"O�!bshs�Q�`�^�[�4�PQ"O ���Q�x�6|9סF
]����"O���$��r)�Kda"��q�"O��F�W��������,�<�v"O&�cř���pWE^���y�"O`�A�K��DNj�`d@K��0�"O(��W��	\�4Y*#���B�����"O����Y J9rHf���|�"OȻ"�ӀQ�؍�����o�bQ�S"Oz,��A�25���P��9���"�"O:�������ը�^�"�0�"O���h��Q��Vf�A
u"O�qaI��0�V�B�[~���"O:uR�	�7;2܁2e�I��Ep�"O���TL�$,6�+�i	8\�z"OL a�U�a�șK��I=58y�B"O�i��fq�p�ҩO�)���w"O� ҅��~���ñf�^"2)�d"O�h���R�h�����(4�j�"OV�P�M�4(�@��&�?`ղ�"On�C��ߺR����������"OV��B�o���eO�"=�c"Oе���P�&�y��(�(�,r�"O5�떋FS$��#��Ăǜ#!�!�1� Yb�M�F~p5J�yU!���T:$�A=N�� hE	*N!�
/|3p�[��D U5�u)t$D�x�!�DYez<��!H��9�D('����!�D�=T���'��6t���⃕Y!�$[9�X�J���	sq���6�ƌv !�D�SX)�If2���֦ӻR!��U�'�h4��I߄y��x;�+-[&!�d�%;��1�g��;~������
<0h!�$N��ެ�c�B$�����0p]!�$չOw�iS��Hlt�	�C��.!h!��S	5ՂP�viH��4��#.�!�$C'c��(A�(ޣGN�q��"�!�Յn�@{�F�S/��y2���-�!�$�;{��&�K�>q&��bㅈy!�O�8�L���'�yi�$���^n!��)B�nL�\�wyX]ؑ�ٷl!�$T��(�����f(QP�K�!�^/+dV���n�a0��I�� C�	x*�Zw�A���)�/ɘ8@C�I�Bs�)�� �-	��{$Z&a�C�I�8(�� �@��$Ȱu��W
��B�	�O��ePdA�1~�Ƞ�C�(#xB�I0x� �@c���~� �1�A8S�HB�ɨS������$=��uk��!�$B�	*���'�<��is0���sB�I��T=��o��@�CNŸ6�B�*P_D 0��ERf�sI�ΚC��5?�<X�j��V[���@�*G@pC�	&2,�W�B��	#���o��C�)� 4�T)��)�DѲ�\&K&`�ha"OFD�$3da0e3�H��{21!�"O�A�2O�5KO.
B�6+@t��""O8\PħI-Q��Mڳ�R 	@B"OԔ �\$oze1q�)X���"O�6��11hňa�F5"��iq"Ot� �&ʒs�h��EC�7����"Oh��'+;P�ٚ�DL�0	�3�"O,�z��̬w�\�ף��c�V�K�"O̘�(\�2���4$ͦ�lu �"Oȭr�o\�x&	K�Ψs�`|`�"Ol�%�X�c���9rO@�}���R"O����g0LӴ������{�"OT�ZScQ11&kK9>�8dP%"Oƭ��m�#uZ�@�����[�y2�]$�<MI �ɰQ&\�X��	�y��A`z��S`� f���"a� �yR������4�2p}����^��yB/�O�.��Sc�37��� �_��y���<x�Ș�C�[Ē�S3�Ă�y��/O`<h�+�I9Br�OG��y�`P�
H��;�jF�L
��bD���yB�5#�(�@#�ўp�BhC&���yd�0x�����!ih���y��]9&����S�K|�=��B�yr-�1 �I'`t��L�y�G̽To�� 7EO�24
|TW��y�m'V44��Tʸ)v����y�,(��	y�
�, ώ����y2'J��l���V'e2��#��*�yb$�N!����S��(��Ĉ�yϘ|��!1��I�ѲR)8�y�J�ks�pb�-Ҵ@���AI��y�Ţ/��d;2Iݎ(^}s�(�y����!锹	��5�L��'��y���g*�U���,^���P��5�PyR��TQ��nΪc�Ac��X�<)�)��j���F�=X\�@3� OW�<���&u�5�S���\�����$�W�<y��r8$<�e�ߛl>�e#�i}�<��C�Q��]�#�-|�L1C#��C�<�c�Q���b�m�(l�J�Fz�<q�g��l�;a �	�Le�7�Cy�<A�'��G		6�EҴ�;��y�<Q`�2Md�|b ��t_��+�O�P�<�T��70�d(s�� [)��8 6B�ɺ����tOC�BM�\��5%n2B�	�T  � ̊�-t!���t;B�	�vW,��׍3(��a"qƤB�I��vx�J��/����nu��C�I�35vai����Z�4�c���B䉵����@�>�B���dM8w�B�	�*Vz-���I�'���`��Q4�B�	�$ܖ��A̳�L�Xq� $�B�;J�@����I�=�"h�����Dj�B�	X	l�{���d�[׀�(QN�B�	 Zv� c<�������C�<aZ%�v�;mA�m�DM���B��"�X�H�R>^a�]�
L�C� H��#�]�ux��k���-{fC�I�]��@�U�r}ҙ�lطH��B�	�`0�0��%����f�.HEBB�Ʌ(8��	�(�܌[�',dHB�	�~�d)���"Gָ�6��(1	�C�)� I�p#QA��(_-�䍛�"O�9ە CY �C�fƟ;����"O^����A�\�8�c@�a��;C"O��XT�Îu��a��(@�P[��qa"O�@Pc�\�t�d���v^=��"O�`�H����H�1N��s%"Oֹ���R�jI�-���E���"O$M�ʉ$ ���ԈY�ni����"O�d�rHJ�p��r'�7�b�D'�S��(K���c"	,a|e�H�.b!� o����FP
M�4��(@�M!��
������Zڦ���۟8H!�d�%~�Q!&��Z$Y�Ǒ2)!�F�S0]�r��/Tp��GD=~!��Z�_
����cѺH�
mC����!�$Ky�~M0�	�#�t�9ƭ[��!��K"1�h�! �ٵw�!�gȩ1�!� D,�c���x{t�qTA]��O���ĉ����v�6IpL1����vk!�O�4�v<�g��'B�0	Hw#]�nL!�΅�L	�E� T�M��Ꮗc:!�*7��PFaH.:�H)  8WHO��4-$7�4�@�_��`�"OP``���&P)��q,���"O&����2fX+w!�:N���"OV�aǪ٥c.��#�/�>!:^���"O�٩����lH~u a�  :5�"O�-Q��@�F�� �7���By[0"O>es��L,U��!T;_����B"O�ey��ˋ:(*�@7� =�t}���'�ў"~����(����d�t��QR���>�O��ä�'���g��/a�x��"O��a��M`DiWnW �F��"O蝁sA�?
l���.K���@�P"OB0�ѵ+܀V��%�����"O��1�Ϝ�� �MҬ,�6`gOf���'�4�]���K)@�a  +D��Q2ķ��Ty5�գ%L��[�%D��x�
�$n��Yc��yQ�BD�"D�,ȅ�*%�>5" �<+f�P��&D��p�i�jxM�S��5)�`�Q/D�@Д����3,c�l��1K,D�P٤�Ȕ�^�b�QsTT��&4��� hF/���� �.EB�50�L�^yB��`�'E�*0�������l}8h��
�'>%0����J���Uf��e������hO?�@���x��Qd�!bU2�ʰ�Gv�<@Ε3'���14HG�>��UB��t�<�#T���i
�z��H�"Y)�!���0K���2�1p�T ��o�4/�ў,�?�͟"���n��;,�;2�э�4�[`"OI ���=L�$ ��,��UbU"O�v'ŧ~L`�Z�풪a�0��g�d0LO�9`Ҡ�9�꽲�Ln|f�@�"Ob<����^_Z�*T�LC�q�"O�I(�	�| �`�I=y5���"O��{���]�*�V�P�ֱ�'"Oj*���U	�#DE�ع�`"O�Xp�_	5�`]� ��(|
B�'X�$лk�|��2͛�<�6��-��'fў�>IP�H�7i˴h�bm
�{�ę��
;D��r@%@�0\�f%�����AE�7D���$'432��3E"���F7D�ѦA�|$����L�Y�0���A5D�� ��"ș�mi ���� H���!��|��'{Đs ��>�p����0ԙ�'�g�^0Z�P�m5zaX��
�'�`�"�e�
!�5 �K7Z�P�X�'��¥�4?��pFF!U����
�' b)Ѷ��ERAR���S�ɸ�'���c��5�M���Q�a�X���'e�x�#��'D`Q���.�h�3	�'�=�w�p��ɀd`�. ߒ�Y�'T��	��S�|3�XԡU����{��D+���
 :Axl�A�_e4��E"O,�8��\ f����
2�a�"O�X�"�"B���0A(p�؉"O�պ�B�m�� ��.�Խ�1�	X>�y���K��!B�y�pQ�"D��dHG#f3\�2���/<���K#��0<�fǂt�"CqdW Sn�R�B�'B�'-1�@����W��I�0+��z���x"OD�(��$�\-3`˝�x��Iy�"O���j'��d��0Xx�b�"O����S�k�N��*�L:	R�"O�Ũ�J�A"fq��1I6 �r�'�IU~ҥ�&����f�+�x�)禅��y�皤qLdPz#��|9��+V;�y�MO !�vA#L��Q�F�yR�B�;7�7[��J����y2�Zy��bB 2�`%���y�(�Z�x#��2��X���/��=��y�ѷ]SRi� ��v.䈀ʘ�y��'�N��ƣ�0v�����4���'thA���JQ��U��m�6F!��'�`���C�"�xqx��ځA粬��'�R ����x>��3@	�=� �I�'?�IW��l\p��#&	.���'������D�5j@p���-GD�C���'6�,�F@�DD8�D�t��
�'%�K0iS�bQ.0ɥJ� P�'s�])�[�d����t<4�
�'Af�I�,^	*�t��d��w'>H
�'1D�k�hY�g~2���W��<�(	�'��3�D01��)0�Ϋv�rMQ�'��p�gi�7Fܹ6�s����	�'q�h�s%͢o�>4����}.���	�'���E��|Q(�!7Bq4Q��$7���|*r�T�S7��jÆ
&)�!
E�H�<�D(%h���`ª͹4U(��R|�<AC.Ӳls\�����K���l�<y�C��5����'�#�4���R�<ͨ �2]���W,�� ��V�<)��O�3-N��'
?l���Q�Zџ4D{����ʤ��
����� "��*�?���igL��zԁ�@�&@�u"�PD�O��D"�g?�� F\�4J��Vrb�l�<!QLQ��s��!H5*��`�<)(3~�\y�s��1v(�@�<�'k�sKA����H�Rԡ1��<�gm��^��Lz�#ȕsҸE�C�w�<駦��aX��k�d�)H1��w�<9�c�>qZ:|��N�\�BU��e�g�<qWe�/���r�%B�\���2g�<I����ǭC J@h�d�ˮrU��Q�z���
H���`��yԌ��l
b��0���Q�� dH�$UЅ�Iٟ��'��%��/��E.�t��:Kp=3��� :	aӈK"2gN��B�]>�T�"O�d2�.�z���(�?��t��"O`�󈅬^�@
��F�'y�l�"O��#	qox��1h0�A"O-A1���h)�*]-��{�"O�|�'�+���kg�S�)t����'�!��5}m�d@SF�X��u�P�ʛAJ!���E�JPq�i']ج����tߡ�$�#ZQ[s����>L$��<#��C�I�Z-�!�OV����
Ɔ��C���Pq&�:�* �0,�3$�C�I�$�M�R����X� ÆEnC�	I��:#��f���6���|�O����8��H�È4I�`p�� 05Y!���'��9CT�X�p�h��OE�eO�Ih��(�����L'D���j�@&O�Z�����<LO6�˒�n{^�B$�H�@q��3w"Or��OZ�=�y��ܝo�T�u"Oh1Q����\LZ�䒱<R����"O|q�.ҕ�����A�j�vș��|R�)J��4�Ì�BUR�����8j�B�	�"sZТ�_�k�����ɜ>(+rB�	>=�j��̴f��p����1��N�b ��®&'𜸋g�T�j !���fV�����<G�6(���L�!�D˘u��ʲ"[�6-�{�j/2!�d��T�8��o	�"�&iC�]�}��'�d�>n����޴h����,!�	$*�b3��K�e��}b����񄚦*��*�$��`�|���L>q��$5?��H�$�]�%�Y/=l��D��h�<�1dZ�@����F�ͳg�>��wɐb�<a
�5��J
��$8��`�bx�xExR��P����@��|u$\;voT���=����dU	^��0�F���YHpL�3�!�]�8u(ffE�'t�	˵J�F�!��?G���iC���qH�J��ވB9�'ga|BLѯB�v����Ϛ �-91�@��y"H�f5ld��[6%�<�@�
��y���3��d�,G��a��X�y�n˥���s���2O^�[wn���y�D�c,-��]�1^��ڶ���yBl��"Ӏ�����?��}�����yrc�	!!���զ��aٔzSjT��y�/��v��!݂Zl��Qm·�y�F#�8���WЌxA�G��y2��A�,|��h֧~;���p≍�yҩ�/@��5��bZ�K_0պ7�ճ��>��O\m'Û�%b(�uF��ܒ��"O@yt�_���)C,.�P��"O� �� ^�6W�s4�uZ��"OlY�6h�`��a�Q6f�ۆ"OF����P�ri���r蔇} "q�"O��À	H?a��d�h�P���"O@E���h���y���:|�����'���(�CD޴z�T �W#��]���#?D���Ϋ_/�ݓ��3�R壧+?D����T�X����w���`�8D��2d���j�A�-)I�xQ�8T�P��f[�{ErD�"#C'e^4��"O��rg�V'�Dܹ��5\J R�"O�U���1.x���$h�jdR�"O������>��M�Y�.4�P"O�T�A�3?$Ph�'ݐ	ɾ���"O� 4@�+M�y�E�A(SH-Qq"Ox5`ㄆ�c���r C0D�Yu"O,�(%Ȧ.��, ඉ�"O��'^#*��ؘ#��B�p�P�"O$�����'�(�{�����l��'�ў"~�f��>@C�tp��w>T���� �y��
���4C6��X���c�h�)�y��A�	Q(�Qb ����n�"�y��N���0�V)I6�指�yҦ��uO�hP��GeH���,��y��\?�����<Jk�9C��ֶ���hOq�R|��."�>d�$�#�|��|�)����0�G�M�E�񏃈K�C�	�U6�̛��mFp���0��C�	�j�p�W�(ٲ��qU ��$�hD{��4_��(�%��L���ɤB[!�y2�ɭ����F 9�]7JT�y��?�l*�)փ2ü��&c��ybdΘ_� ���n�75��	�DF����0>�K�{J��B-׆<��Rr$	^�<-=N��膕*h�m�`Dl�B䉠n�Q�mٮy���;E����lC�I�G{pArv�|�Y!!bK��5D��c o�*K��3�N���d��/D��3��G�6����-�J.��
8D���-�m#F<��MӸxeL-qi7D��b��O�h���#��<a�i�	7D����M5LEp� ���e����6��9�S�'n�$�� ޘU�Ll[���;MZrm��k�.U��j�<F�����Y:F�|a�ȓ&}f9�����1p��/���ȓ~�Z!q�v0A����!�ȓ_y%Y��;p����U:΀хȓ*�.Hۦ(^fɈ�0Vm�	U:� �ȓw���N�.d<@�N�0w%�1��Ig�'�b��W ���
�y��׿`�6�эr�)��NR�,�-B	`ltD������yg�,�d��U���\1dapuj  �yT�i(����� \�0�$+���y��E&D8C�ֽ F䠣��y��>Hv$�v͘�s���It�V��y��"k�4lc��T*r1���C$�?��?�'��0��1F��ЖN�)z���
�'@�|A@áԨ�5a��J��b
�'Me��l��.��աd�	�+��ؙ	�'�fpy6d�#E?�\kc��&�~�2���yR�Ո~U���Dͷ�sp��yBa 8#8q���A���1�B��(�yR퍮0T��L���B����Չ�yrh�1�*����`�abܒ�yR��M�i��㍭ќ����y�d��^$�e��	���`j��Y��y��0M����GF*��ѵ���y���`�㴥F�Db2���F��y2]�x��0atJڅE���悿�y��ا&�HHB1Ƃ16d�z��Y2�yb��;UHA��L�+{^�ۇ`Τ��'�az���M�p�j 
Y�4R�r�E��y")^�mq2Ĉ�e"���.E��y>AF�d� b8�$�rfZ��yr�	&5��-� d
��
�m�0�?�
�'Qu�u�ΰ�B�'��ap*y��'H0Ex ���R�P�/��^��J>����)B�?N|�e(_:>A�`e�!IJ!�� ڔ�a§�̨����}��5��"O�q�ԁN%0���C۰s����S"O�1X!�^"�,P�C�X*r���"O���e��x�言d�<6�؉A"O�PÂ&�,H�L�HƆU�Q��5Hp"O�4����E񲁐UF@�x�d��G��5�S�i[�J 9���, O�����%ў��ӣe�B�8�
�*tШ��R�B�	�:����o.r���GߨE8B��%q9�y���
�%�Z4��F�&�T��p�d@���?\?X�)E�Đ*G�!i�I7D��sV�.�92c�ě�b5�V`)D��c�Q�$dM�@X�$U��+3D��� ��GD�uK��U���q��2D�p�4�B<ʥ�����U�!Z�!�G�}V*� 3H�4l�ܐ��̦_~!��8G_�� �$�(����	3?~��W��(� 1��U2�!�Ɗ�X��5��V������\d]�lP�VP�ɨ��'p�B�I�9�$:�/ͫU��eH��X�a^����;�	&8w����5d���Α�Z��B��;r�\9��(ܾ�i
�.�4:�B��=Y�b)�W��?L:h�Zv	��4�xB�%�ti@ulϲ
$ 3f�ږS�\B�I�j'v�P E[q�މJ"���2����0� �0D
)�|A���/澸8�&!D��X�P�Czԙf�la�b=D�T8t@�Yb<I�Î�.�@�aF¹<1��品e ����F4�����g^�-�bC��;R�b�ҀfQ��a{��ې[ؖB�I8�~ۤ�*O��C1���A�:B䉴` ���Q&�#�V�Q�#Y2o��C�	�J�qS�)_##޹{�n~!��E��L�
"bX e���y���:Ro!�$ŉoR��RN_/(�$��UFPP!��	�G���r,��-�����sI!�dX�O�N8�&Ĝ�gl�뵌A]P!��۽5�f�ь=���,��7�!�d��&Ut��㌋b�H|q��;m�Ib��Թ��Ӏ�i���.0�u��H8D�t�E0�n��C�����Sk*D��`w�Y�
��'�&�|\�!�Ą�ZeƉ	��
�@��Y���\/!U!�䍆iy2)C�����c�m��LO!����y���
�Jp0�W��$E!�$ȃ*!ؠ�'Xh����N�4C!�ׇm�U����jNP|zw�d8!��Q� mf̓�瀻_�Z�	'�^�!򤏙l�]��If�x��!��2!��$?�Z�L��)��#�]�I!�$�$�Z�{�Fz���:1!�dv�%Ac��P���S0�Z�`�}"[��be�3g6`�%��{���"O4{�*Մd�t��̶
\�m"O��.�p�ƀs��P�:�j��%�'���G!8e: Fۍ#�x@
�+Kw�B�	�:�X�0@		�_��'�W2zZB�	�tR�
�N\ @K�o�B�!�B��C��c���υ>n�C�	�\򰱓W�����A2��H4{:ڣ=��'i(�\� -"�SM��z�,�����X�A	BGڔ�Q�f��=K �kc��FR�3(�7'8���ȓ'� 
pd@8��u��%^(9o�U��S�? �\*(2k�j�"Ŏ�Z��Q��"O2��
U���H�MB*T��K�"OD����D�m�4X0��:QE<���"OLUPO�O�r0#F-U$:�}R "O�ISU ��w����V��!94�#3"O��ӣ�NW�t��,ڰA(�B�"O�� ��K���ӱf�n=2C"O6�0�gpvl���L�'N�ų"OP�Y���)>�dyT�6QO�SS�'S�D� hIC$	a>p�rH!�F�CcҘ��j��#��Т�"Ot����,�����*�9_�J�"OP؋T)��F�qK#fP��b�"O�zdIM�J!��0�F�X>�|S�"O �sǤ�}�N��P��t��$]�!�d�e�t�����&|kl�
@�9u���i>Gx2K�+ Z=b��
*�V�Ӕ�]��hO����O8lآ��g%�8';�ȑ�ОO!�dD�J�t�����(�
Xb�&��!�$�>n\��8�@��$�~u��ܢ\�!��(E&�*���@M�����9s�!��$�d 8�	�7(�k�e}�!�)L����5
Ր���A!�D	�2��0���&�X�bξ!2!�Dδ2�4@b	t��D)�?'!�d_�[T��!DK,J���Ƅ��!���Lʄ��B2>$���ϒK!�D�5<�(�taʿ&h�w��!��� 
�(D�aHU�D�ґ// "!򤉟T-^��G,PK�Z�+²@!�ЁG���%KY"�r끋_!�*h��İˀC��#a�^!�䁌_���N�5����E-7Z!�D�ӊ4A���\6�I(�e��T'!�d 8u������X)�,1��x�!�Ě�N�蠛a쁛9B�3R�^�!�!��ڗg~=8�C�,0�y��,�J�!�$K=6��4�be�0v��!ֻJ!��$l��UW���i+��c��Ӏ!���@o���ȃ�/+
��%!��\-t������(�L��"�4x�!��sj��!���++��a�� �~�!�5��
��t��e�I�B�B�I ;	��3���8M��E;qG��mvC�	2����/�&J\v�STlۖ�NC�	�R�� 頩-�Z�2���9:C�ɶY�hY����d���,F��B�	++����fA
���ÔCQ�
q�B�	?a� I�-	Kx��%@�;�ZB�I� j��cc�ɬe�nH�q�B3�B�ɦA��A��4f�|���)���FB��3]�=�˒�Py$)D�B#X��B�	�+ӌ|S�K-a�3�L�:��B�I0�H�5� �^�|h�
]�M.vB�FX�	��H�ĢF�ݴ_�6B�Ʌ=DJX � O�˾�	0.]�(:�B�I�u�|�gi�"H�Eΐ���B�I'SfR��B`ߤ�x�����K��B�	�!)H i D	T{1�J ߖB��1��,;W+�������1vB�I�^���33M�4nm� `�!5/PB䉩0qj�B )�R��z-˺JmB䉫7т�ɗ���8��u�h��B�	[�.���IY�s�)21&�y
� Πp� o���a,Q���{�"O>��@.T�hz�Ś�L��O��
�"O8��&j���f@&aF5]L�"Oȭ���"h���[⏋�.��q�A"Of��ʇO9��H�.�;k�>�PE"O
�C��yc*HR�K�K����"O�=��n��k��++Q�ah��@"O�D2��6�b�D�ROj��r"O ��F��"������H����"OB!r
4�@-���Jl9�͑2"O��K��^�l���� �D��"O��񄆍�<�Vp0 \Ϻ�!g"O>�{�e��B\��@�9b�� �2"OqI�2����0�;� �`r"Oڤ�f�K�Bc{�����.��!�$O56F!)��s��8��c� v!�$[?<��e���O#"L%��B��oo!�$�%;J��%/��0c,ĪU!�䃞9��I#E��l��q�A�f?!�ă�l�Lm��E��k���;��&"!�D��`0ֱ�ʋ颅�@IJ(!�d�~ޤ=��nV�1�IX�	��Uy!����s�Z��sJ�k�`�i��?np!򤔊���Ce"�h���'68_!�B�][�LS�`�\��A��^�!�G�9�x@J��,���ӤS�.�!�D�,�j�����qB�����!�I�x�Z8�S�vc$%[�G�@�!��UB���IJ*���'��	}!�Ḏ"�	c��Ěe�~"gf�2!�`��FH� 93V�Z媘6W
!�$�OL�iU��21|P %�@!�dH`�X@qP)ݒS$b����G�!��*flJ��fL"?	��[@�<u�!��X�
o��7-�\��@s5�ݺ�!�D�PCh*���(�v9�a�à_p!�1yQj��1�-0�TMr�"&_!�DT�Jh ��@{�F)
�N�8U$!�d�]�>�*�g�.:+����X!�D��~ɢ��Ņ#1rq��`�>P!򄞽(��t�߬#����x�!�d�C�D�oVRAq{T��$�!�@J!���E8<>�Ѵ ěd�!��,*�]�4�'LV��p���)W!���) "��6G��&RusF�F�j�!�H2����)I�P��y�-�=L�!�D���y�u�ӟ����_�s�!�$�"<q��	��=kn�
�#C�h�!��1:�Ҭ}k�)!(ך$�!�d�)EڠP�J́wg��=�!�䎠K����1���SsƵ�FR%�!�D�R|�p��%�Wfa���<!�D�+@�B���_�
Q�����!�d��+JE�#�R��d�/�b�!�$Z�:�1Ţ��!{v�0�$�d !�D�?x0Q�'�:B͎)`BdʇA!���!���7�<��C��!��Hl�e�`Ҩe��-�q���!�Da����@��D�ো&?�!�d�b*���I�UlP�kGeQH!��Z�&l�Q��6y� 9�'Ì@b!�G6����G%�a�,SZI!��~�X��E,�Av���M�y=!���,(n�ոv�Z<'�t�P��k��OX�=��� �={ 
ظ�B�Aƫ��7�J�"Oz�Y���(&/�X��ٴ�k2"OF<�F �a$X�p�i��Y�b"O�@q�@=؊	��H�:G�����"O��!Ӫ^G���1c	�]uFxp"O� �
3k�h�rf˱X(1
"O�Á[P��A�T�k��2�"O)1&KF(�NI;6�[6XN@Iб"O"\���ޱ-,��tU2l�DQ��"O�=KS�\�U���%���̦��0"O���$ΌE�����V�M����"O�$��.*7��3gV�@��3�"O���M]%�V� �f�z/��3"Oxi�&n[�t؃�E72�έi2"Ot48��� �V��E�E�&��P�w"O\Tkr8��Hǩ^�Qw���"O�X��i�e�v���E�kaȝ1e"O }8��/@D���[�fй3"O4���B��SCR1�l`"OB�Bq!��{{�)`G�f�����"Oj��\��B��>��E��H��l��'�ў�>9�v`�/�x9K2U�� �m/D��J3mT�>��h"`��5�P�h3D�h��L�M��@��gt�(0�%D���G@�<�XyBc��&`:��"D�d�D�>J.T8�G�!v����4H6D��aU�ɧ	PtI�na�	�qg6D�<�elAR�ɔρ%Y9�ݳrN0D�h¶�ӿ~\�eʑ	^�F��$D��Ni���������'6��C�	�$D���%�̥c�E� #�C�ɉ)(
�kU%�'F�!{A��Pn�C�	�D�Υf���>	v U�X3�PC䉹?*b���ٵj$��刔5�C䉋{�4!7,��JA����y�C�*b<�\��Å+'7:@bAZ K��C�"<��	�j��*m����'��C䉭u�<�G��S�$�I���40x~C�ɏ�fqk�	I�Lv��W#[m(B�I���H �D���&G��TB��=V���q��I�~���#p.�4[�B�I�<ԘXD'ފ���$��8��C��-c�����	ɽ6��	0����4C�ɍ,N~%yV+U�ʼ�"���NB4C�I�
����U���&�J��FAу:+`C�I�4�a�cT�6�(X�'�=)�`C�I�|��D�@���9��;�fɷ�2C�%FI��醇�֍�Js.C�I�r��0�e��2;�����~)��D{J?��2�J�wK��BOڄix�i�v/4D�hB')����F�14����.D� �@�2;����H��mǈ���++D�|�S�^�[��ɓw��-@�X�`��'D� C3��6 ���#�+)�
��R&'D��񅒒5���Ǐ�t҈�%�1D�9I5�0�;�!L.e��4���0T��y�F�%v�r$$�($"#"O@\�a%W�<j��v#��:�	�Q"O��1�(�X���a��T�R��U�#"O�x3AfL�nR�q��B��Q�G"Ol�ؠ!��,��iCp%=%Ot���"O���V(R�@��<����k�|bc"O1bwn�+�q`$�0q��E:�"Oz�+F!թyY�T�g�Ie2h��"O� J\���ՀsuD����@e: ��"O8EA!aW?B���V@')�L�1"O4�&ûi����3����4��"OHA����V�F�L?^����"O���GmO�}��I�B#Ğ,x��2 "O�0S"���D��T`R��(��%��"O�l+�/��{SPYe�)-���d"O:[3-�.L�
�p��N�Z<��3W"O6�a��BHZRϔ�5H��G"OX3AL�,Gw��#ӍZ�d2j�&"OV * (P1�&4�i��Z~�|��"O���T?���z��4%����"Ov��1�\j~�Ï_m�H�u"O�T�!Ί�]�0}(P�v|\��b"OlLj��ؓM�DȂ�K9=x-�"O��XǋZ?$�B�`H/q*Zp{�"O��GШ�Ѫ�Nu
�j�"O�
a�),�n�ѣ�0h���I�"O��/�
1"���F<��0�+!���!ۜœ@ϛ�n$�Xу�'-@!��7��]��d\l(��19!�ė�e"L�`��+�<��)!�Y	F�|��Po�m�`P �(D�w !��?WW�ա�d�G芩��(�_�!�Z<Q5ū�X��^0�T�ѥa�!�Ě0��=��Kլ%ְPk%i���Py�D[�H7`ŐH�a"�ٳC ��y���
^���s���40tzQPC T?�y��'����ո9������y���	���
ڷ�(�R�1�yR�N!Vo�Ӈb��qSV��r\��y�&�\t4���W g)�*/���yҌB}X����R�H"��{���?�y�%�(g�,��I�@�$u[�d4�y���}�7�7?ƄI��[>�yR��)s掄z�J�;�V9Â�ߍ�y��H9�Xck��N�c"�&�y� R�}/� ���(��!��k&�y��""�R�[��bh>mJ6�%�y�M7,S�H�#US ����1�!��ФZ�XT:v!¶6�F�i��H�ko!��%(�8��щԏw��u3��;mP!�D�.Tj@���b�@0$Y4È.!�$�Xb6(Z��HL��bB�PQ!�$H�[n"�uIA� ������8h!�䊃c~�e��F�#�:��ӊ>0!��y���!�c�{� ��EG�!�B9�%G��0{�9ׁБ:�!�䃡Y�\�#�/"la�E ��!�D�.)���z���}v���6%�!��T4x��B��r:E�I��!�d�W�&I!d�=v�P�JÏ���!�d�z�z���(D�X�|y���2-�!�䆽}z�T`����c���E�N0Ag!�đ=[E����(L�� ��B3J!�dZ�B-(�� �0�g���7J!��>@Q��`�A�$��"��
F�!��Y�6QJ�G�;ȃ���$-!�$��
�( �H��;Y���w���!�D�$n֒ ����')>����h�2}�!��j��)y���C�fm�(�:T�!��T�Qe��Gj��{�f�)�!�=TՌ|@vE#Z	�=���R��!�
�!)X�똁{Rݪ��/-�!�� �`�F�W���/V�Z����"O8�!��t��1s��ׯ���e"O��ұ؁Xr��,<Ǿ���"O�E��$�L"��Q�ڶ\Ÿ�"O��Ҕ�ݍ�:D�B��?A
�E��"O2�ʥ���J��XrW �3��h�"O�	���~Q�WOҹ]��,A�"O�p�Pk6V2�D�6� �3ऩ�"O��Qr�ק �1!g�'�4�g"O��It�S�( c�G�H�iG"O��8T��b���Y5�V>,>�Z�"O�H��Ŏ?3�\��ւ&/m�#"O԰�ĭ 1�֕���|�,�"O��Z�J�1�&T�1�]�Q�L��B"O8DZ1#�->�8�S��+����V"O����	B	��X h�54t�d��"O�p�scúe7t���͞e���"O� �#
T�@���pt���3\LU �"O��БȌ�^#�a�g�/�^�E"O�j�@��a�@����VǞ�""O|ݢ�`�i����@��Zs"O8-�aBGN��y�q,_�F�"O txA�t"��s�_3d(82'"O����GɫJP�TK�?��0��"ODQrWÝ�gE�AE�Έ3��19�"OF��`�Y�nL�JqA�#2TZ��d"O��B!Y�=.�0[��8-c��pV"O�M��9G�P�ӴA��\&��a"O�͓��S6e�ti7�.h����"OR$(�L	6 ��`@��5�=F"O8yB���Ё����2�k�"O��bc$ʹ,�@l����)�. �R"O��PѬ�+I�P�f�Tz����"O����HS�dT�1��L�0��U�5"O�S��	�h;ĥ����s��-�c"O6͘�I�?s60�3�#h�ƙa""OکC���_3
=�v�A�w��]��"Ojы'-�	~�p2�K�#;8�R�"On����L	-xâ@��/�8�"O�MPCF��S`�Q��$M�LV��"O��f��9�*�DT�>n�x s"O���L�ha�- �{����"O��ڕΓ�I��۔Ε�g�e�p"O��BL�	��8p�I!N����"O��Scd	0n�
���J=p�`"O��
���Tf��"�"Od,�0!�$d^�	��/H���`�f"O�8�#*��T�|��n��ii&�[""O���:j�P1c�*�:��"O}�1�J�"~05b�,��$*�W"O�%�+,&���eJ��Av��T"O���ǂ�;������
�.q�u)�"O`���c�	gy�8���0c���2"O�أIQ.g����IzK`�k "Ol��팷.Kp�	��\&x����p"O�թ�#�,wF��P�	x/����"O�-I�������C�y�`�_��y�ўYlX�!܂ql�x ���!�yB�O�8ü�°L�z��s���y�o�"�cV�B%p{b [�L��yr�I�5N	����n���C�y��J�NĢm9A&�'$�Ȗo�>�y�^%�:��P(�j��%���yb�cʮ��̔�\�"\X� �y
� 6X�djˮS��}(��A�KY��c�"O��Ƅ�>4���b�	�n�a� "O�9ZUk��hcd�`�9t�8�P�"Oh�H&I�0k&��B�ʔd�I"O�-
4�4^��(�@�Y���#�"O&�hC��4��=����a(��'"O.�I�g�� ��7hߩ9�D�"O����B�)f
z�(�F�!|,���"O*(r�o]�:��,:�� #I&,JS"O
!�r,S�>�����e@�fj}@�"O��)ӴS3���Sd�pbjd��"O8���	:��0��R7��1"O~(3��$yFH0c\�G5мC@"Oh��fzQ�,��z2��5"O9!4)enh��@!�z%<�
�"O��	�E�֐�!"�1��\�"O�<�* ��a8��8l� RB"O��(����^8F Z�-|�MA�"O��A����pk|�XbEļv�a	"Olm�3�L�1��l�s��2gt�ܸ�"ORհ�[�C�p�1���B�����"O؀��%i�I���	�r���"O^!c�k%[����g�S�ι��"O�(��	����%��I�le�\�U"OP�kEL�a��a��ͅlQ��C�"O$1�rGCR��Ԇ�1�:��"O�I��8&P�yj��žz�x�7�?D��rD�L	6H"ID��p��HC#>D���o�-%'�LA'������9D�ȣ��Q+��tѢ�ÜQ���7D�z�'ۊ����r녔g^����4D��QåK�hB�zC��-А ��4D�0��A!r6:��Ӌ�.sIXH1�0D����%߄d^,%��E/�
�HSH*D��(Ӫ�A��Jt6%O:e�'D�܈𪌙�n(�0 ̙.�����1D�P���0=m���i�!-��g�/D��j�jĚG�ٺdb��R��h�:D� �G*�su��*\�wD� �9D�pk���&�����TBx�;S-D����2%?�m��))lb�
-D�� 5	g���ՃCA#&x �i-D�(k%�%*�0���I����@)D�<s��'e��t8Ą�$,Qa��;D�,�&CG�e��P�/��x �y7D�8�S�C�E�D��$Q��1�R�6D����A
'��q�ȌjX4y!��3D� �w����� �#�L�o���f6D�P�r',Ev�Z��˨63�ճ�M3D��`��
�>>6�	3�
�|ћ�a-D�x[�{���YB�	x^9p�+D��Q�MI}׊�J��J�d����(D��
f`@���̱��U<*+p�&D�ĩ�67+
80�Ӛ	��
��'D�\k��%h��h��Q�f��<��2D� В�X�J�l��h�)u����+D��1���`�b�鑏8=2�)	$M/D��QBɯ3�l����F%�ah6�,��p<9�#�Q�4P$o�� �`�R�S���?�!A�3��y�U*�CO`!ȐCR�<�%!_�z:>�6
P7kV�C$�L̓�hO1��l{`�˱.�4ű��23�j�
�"OR��"��gEĈ`O�=V�8����t8�|��E�n6�l+WG ��Y�j.D�� �i�KG�-/l\�s��$��a��'��'���r@�ߪ���K@oi�)!�'��l��f�h�*ЄSrB����:�S��d�V��9A���M�@�A���.�y�ω(By�� �]�1~~��#��yR�:a��ASe��7/>�K��ֳ�y"h��tr��?@�TcR돳��;�O�L��R�:��@i�&Ġu5N}!�x^��yCe&�S���*D�ĠT%0(HQ*��[7��?I�'!\�����xR��#bA��E�\}!��7���"~��@	&U�m���l�1�NW��y�e�?�XD��#Bъez@
����<y
�3�d��D�B"N�C��K�QВ��<:�����P���*�G�/AX���ȓZ�N�{���&���z���w�ԹEz��'����peY�LS(���.��/3p�1���	p���*��9���k�JU���1�S�Op����G2��]��E�u��h��I}���I�7!c�4�#I �P΢���5f��d���	7�I?qؐZ�	R38Ő h�# D����e�>����T1#�>��*�O�}�'ٛ��s�h�� �ݭC}"��TN��y��dMF�CIM+���#�ގ�y�A�|��`cT��n���BVd���y�=|8� (Ҕa�<����N��y�i�l2e8���'EM�\؆$��y򃚵#�	 a6�����I'�ybKD���1�Ƭ��;:t���'1�yr'�u��%�S�L�+����Pŝ>��D>�O(`zPc�>�|�js�hc�h@'�'�	�n�<ӆ
�DZ�8�:k3�C�I3kP�C�B��f����#<���?U� Kת�"(���Z����k8D�|0���w�D��栞�~�L�2�<Q����K�aA��+����ˎ�!C�z��I��ؿ*����P�
a0C�I�l�2��2�M�/�|��f�#7i:C�I�!��]q�LY�GD4�QE��%��'�a}�eEl<�����P�쐪3�ƕv]��=�~"1K�>QȜ�%�  ��㍾-t�!F�n�<���<h�����j-b\��-�y�����(On�0f��4�FFf�`�f�)Em$�Ұ<4�>�Qj��|��$������v�U��E{���'��mg/J�w����`-��M:C�I� Z��p�	[#��DJ�&[���x���Ox�=�OD���A��ex}h��^s|(��s*��;�`��$ H�J��K�sl��O@���\w:(� ���9h���A���0���Fz�<�Za��ئ�����隋���x "O��pƭV`��Q�)կ3��	��S�'��>��- _���@F�9�p�ٱ
�
��B�	�Z�=����"7e�H )C�z��ד�?�TNS�-�x�R������UI����<�]9R�R0�JC�qsEE�<%�2 �4�q.ĴzP�e#�gVCX��Gyr���c����j��$��en��p>�N<!�lIr�j	�D�Ù���b#Mc�<A��_�<�8�{�&��LA�����\�<��M�3�&��#��~��� �Z�	|��J�<I���]�Ba��n,�O@�H�q��,�<��#Fѩ���ȓm,
�+ηKe�!˖��#�% )ړ�0|B��H�����i��U��Y��J�<�D��2�4��Px��9�Rl�<� ̔P�hC)����#�>[�ʸ��Oj)�Ɨ+�m��6ڐ��|[��_�<Ac�Q$`#�i7��' �
�k��@�<���	�FzHxr�L�!~[~u;�e�V�<iS$Ɩ\ ܡ�d��i{�,OR��hO1�(!@j^#*`0��(�1a�U�r"O�,�E��&ިT���U0PF���"Oڍ;Å�s�6��D,ȻT/���"O��7��0���kE67�"8Pc"O���	!
�̰�)D~����"O4Ȱ��U=T,�����O��l�"O����@s��T� �	> �#��IT>i8tDG�e����Oڲ;DHV��yR�\�d"�iB���4���Oʵ�y2��/UZM8��ϐ;ʤ�R�D���y2
�p�`<(����: �t���L�yB�d�8AH�=I�������yDB%�Ѡ���!AIh�����'��zr���X0�fF�fgj�;U����O��~�Ӏ3�j��������&ԕ:�!�Dӵl��@����=L�"93V���R�!�dC�W�N�z�D�����X�!�$K\��@Y��j��
e�Ǿ�!�� �D���j������E�9t!�b��]H��^7D'8|j��FU�!�$"g
�AJ�����i� j16�!��O*X�����Pa:�jդ�h�d"OV��u�I��J+#��XA�'lў�S:Ŝ0���R.�|R�*D��д�J7*ɤ �R��(�h��A-'D�\JQn) ����X6y�B$�d%D�d�q뇼��m��@�o$x� �$D��+�� �2&i�	 �� F� OH��ē7H���$�ҸV�����
	�w�BYZ��?Y��
R(sbgO�f�����5<��-Gxb�)���)x��P�ŪW�t��ΟW��D{�P�,V,q�1��*Tv�l����."�C�)Fxc��Q*a�&��R��ٶ�ՠ�yB"U*V��C�eZ!JwdI3Q����~�kI����0,�+W��'�Qtz(��r�5D�8Zt�W�%�����P8���gC D�<񵧃�L���G�M-;ȁ��O;D�(Q
йzu�Ђ�l�!\`�;s�9D�h
���:�ڡ�"IJ�č��9��D؞P�LM�X4�O-\����w���=E�d�i��sT���	�8LxlHW/����'����ӦO%Y�ّă�K��3�'�kE�[��&�>@θ��
�'.�@�.��Z$�/5$#
�'���Rb	ѓF��J� �.vgH�	�'O�sd́���4�Fe��2 C�'�����C�d򆀑{�I+�'޼�U$�3O��bȕkn4D��'�P��^�X�z�N��/���[�'1�Œ�b��M�B��TCH�-�p�'��h�Č�wJFQ9��U�:uB�'����.W#k��C�D[�r�c�'��؄�ʓo���rC�=�����'֤xz��ʨOp�5 2�DBx�i)�'���%!��T�l)���Ż7�^���'Y$��	Ȼt��D8�ɹF����'�� a��
�8XČE�E
� b�'rr���D�G� �$]����'1����Ib��|8�f��g��=�
��� ܝ;��:�*d��J�F'P�p"O���&����Lk�%��&��w"O8}��ˏc��s6�	�8�$�r"O��`��8��E� ]�V�)g"O6���O�ߎ�B ��9er廃"O����%L����`�::H�`A�"O�X�jT2�b��c��3_ ��'"O�P�s�J�KoH�m�8��R�"OA��LX2V�Fݰւ�/�ɱ"O���b*^�L�.�3�h�8�)�"O�5B�Kկ4��5�t  e�R�bF"Ot�j�����BRE��M�}��"O����
Q40�{�	�E�BxD"O��6$�'ƊJ��V�g� �a�"O.��%�V?<�p�d����Mj"O����%��0�\%�RfS����"O� �s앛Yg�����)�AC"O�x�A�G(��斢%T��`"OB��@���a�ꉠ���?���"O
�
��!AP`�fƍ� ���z�"O�4ɴA��
H���$ h�؜s"O
�xD�ڻv�Ne
W�aP���"O���4%Q�ФJ'��rF�MH�<A3ȁ
�6��C�.J ��g�I�<A��t�"I����;��Tz�@KC�<���H�z�q�V�F�[$��)�/P}�<q�����F�p��01����M�<�U��s���F��S�5��]Zf}3��N�h[�-C%!Z���`�M�Q�TqA��[	>B ��G,D�8ő�#rY גZ�>�HÆ&D�|��B;8��*Q��K�P��J)D�pS�K��9�dl*kP���0D���aF@��ը��Q�4���" 
1D����M�J���8��C@i�h"g�"D��"�]��z�f���jp�!D�̒ס��}� ��E�8];���A<D�˔*�HnX���mZ�p��8B��0D�$�0����&��Gخ^�9�$D��i�5�����*١?T���#&D�8�
�Y��5��W�*QnDAS�)D��R���'$}-��FH�$\���'D��)�@93�f
�C�-|&"a7D�P�ǉ�>[�B1k�
-e�
ЙƄ(D�4:�C,;WPt����u��k��&D�p��,��(���f�;]Z�ۤ(D����JC0%ӱ��;)_<Q ��#D��%�{���A��G�F^*\�`�;D��X�D�}H�[u�ŹM� �y��9D�X�D��\J���6-�/D��v� D��aO �4��S!Jj1�lh��<D����K�2;~�cP��b�� O;D�0(��5 ��K���F/�1���;D��˱!E�%�\bP�ު�bYB7�'D�p��BI�� y�	6�؊ OB�	FH��*ݻ{N�9�䄕���B�	!d� ��#G���zu��Q7��D�	�2�b��4����fR`t!��J�d�28:�#�0afX8�� 2!�L�8NУ�i�:�0yХ@vp!�䕮6\��t�	�4<&���<i!�Ċ�y��uz�	�@�nm��G�=l!�Ā�_"AhC�ʃXh����}*!��	+-��Aۇᆀ?SX�U��Y-!�$��lHaf	ΕB��x6+V�~�!�� ^d��nK}��@��c$|��a�"O���-ͻY*�#���?��m{�"O��8 D��N���Д��
Z"�R""OD (�&N1|¬P�D�Ǯ1KJh�"Oj�9�K^41�"�pR���R�3""O��;��W�(r��ZjN�w�B�`"OR��'����Rv��'�z��u"O0��1����2�Ԭ�"O"��`�\�(���Y��K���"Ol�C��Á'V���
�@�A�"O��ǉ@�_#2�+���7 �"O)"�CA �Q���;Z�0�"Obx)T%.p!^��S������"Oi)Ƈ5m���bh%��PS"O���C��5X�����W���k0"O�	��ע��¤�1_�=+�"O$�y�
2*M. (Vb�'w�<1��"O�a�7CxW��5�J�����"O�$	�����3J�r�<Q�"O��$ D"G"�\ȅ��vM�R�"O(��(Ӏ����Fb�f=����"O-�Fl�E���hR�.Iv Bf"O4�B`�,بM"B�DQo:�*t"O���ӫ��`x���g�&*���)T"Ov9J�P�/l&����ţW�T|��"O��i����1�@�23�Ic��h5"O�I�Eҕ
'L\x�%�<f��J"O�T�iF�1(L鳃R�u��{�"O���`�y)���⃷#��@S�"O�y8խ�S�� 8�!.}��`i0"O�҃�-�,Z���)��d�x��;S�1�=�~J�d��)�r����ыE�8s!COj�<1S*�!��
��؄@M�8����"2� �'���i-C=ĘϘ'6,����0��ti5/�8��3��v�hT0�܍B���ˆ�5���:��
 j{��l 8Vv݄���(逡�a��g�<IS�@M$���>��n�*c�5Q�j�5
�LJ��V�j%K�b�~����LJAX�"թW� ��=y���O��
W�%�eZEP������O,@P�S�+�L���T�N#r�Q<��z6�&J2�bYæ9z��[=A�⤇�ɪE�ؼ`�O��	]�Y�g��|'��jg�@5���۴x�J��b(z�K�j�,��G���<�B�"*����ݦ/�9�gCOS��Ы�ɔq髧��of$=2���70ft������a��Ңq�YqS�F.�K_>Z���61�'��ጇN��,��N_�^2�EF{	�"B�h�A�?;����cW�p�0���kL:��pO��5eN�)4]�	����(��u`* ��O�##f
�I�D��CE�?}�mP��'c���TJՙ?_L��a'Y`��<s�f��K���܋`�C:s�pI�h	�&1yC��ڼ�.\���o�()�OV���. %b޸���V�hc�@C��(�`���L�|������B��S�4� D�u��'� ��6���1Gݨs�B�S�O5�����I�4���"�[5䐍�����y�������J ���+/�4)�HIIN.ɱ�U6턵�'7.%�Ĕ?}(Wa�3O��%A�/�t(�RF!ړ�A�2� �n=# i�%���1PA�,J�a�5G �հ�#�-�[F�o'P{,O(�H������	�
j�:�鐀t��b6���9QB����Q�) 		"`_tʳe�	 ~�
�I��u�1�n5�VH�s���CmP�pЁ�DN2i� Ii���*9��|�lSuI�1X�kK.�$������]�&ii��ނ��L���ӛ}��D�M?u�ҥ]�5� =�'D���I��g�h]��(��s.�9�
��x������[��PEX(h6��6QT�=!��]aq�!b�P{u�i!�'��y��J�����J@)0��[bDr5¹!v����O^0E0y�P���Nƹ5�h�@���TlHx� � )�6�Ap�܈+ɸ)k �ŶqO�=�"ێ��O���qA_�[�Zq�3�����8��OX���*K��2y(�gYLo�� /�K���	��t��%)���x�& a�Q4l��yb��*������(�\��I�=㐠JpQ	<�:��-��=�n�[I?E�%%�)y�I�Lq0l���H�1 Bɫ�L�s{��D����p �&�/[0���bK�"u��8!��<j��5���-��5�V�8���I<|ʑzw�_ulҜ��#FP����T�R�4�{���5�M��ڃ?{�� H(p��Qm�K�L�L+��A�K�!�dT�Lt��8pM�+S]8�c*u��ɠV���!z��1=H3��4�ӮOI6�J�+�}	 EX�DҜC�ZC�I,�X1ؒ�Zr��(�m�o͊�'�v���GQ�k�zd�p���n≉g��	��ŗm���xMOK������d��ٻ�g\hd��J��>��4b`b�q�U��F�� O�.�Д���$���D@�=@R��#f�j��@���j��_2���ca�2)<�C����0!F &y\��4)��)r|���Y)W�Q&O�ҧ(�HQ�tbK�� �!P+V6J�$��F"O���@�\�(�6�P�&�^��0)�Y�䈬N �� Ӂ2��$ЉyV�QyTO�(&����"��P�}\(`�$� Ʃ8f�R�
|�2�˃�mF�u��	cG�scƙ�:`�=j҉ ����?9Cl�d�䘩׈�'�&�j�O��DB��sIs9��-(D�`jA��W8l�1#%^e+ ���h"?�C�
=�^H�A��N(�蹋�)�"y���r�[]��
� �30!�Lɼd��J�m�n�C����z^����,�'c~���I<�ѹ���|n'x଑c5m��uᬀ�g���yr� �F�~�����?�|�Q&����?yD*�8Yvz���7lO� r��Z��^`jGE�,Tl��q�'V�Ђ�E: �(n��C�.��4C�����6ND�&��B�h_��`��V'�����,&��������2ܪL���ӛk RD��͈�*s�Q�wK`B�	W�$�!^+DJ��Ŏ7ADtI5�Ix��H��D��'����D	C�Fi$� �76Ly��'yy�2 �<Q���#�ҵ=�X���+~�C�_�<�(���܁�*HJ�ݔ@
Y[�e�T�{�@Ѵ&Y��pu������D��X-����+,n��4D�����):?��v��0��q�N6#l��z�)�h�n��TL�"e�� f�A�Q�aY�"Op��P�J�2hp���@w0,
G.�
ݹ����O�#Ȉ�Ey�T��oB��j1"O}z��V	V9z2]�}��%z�"O�0�2��Zc.���$��P��\�v"O�wnB�@x�2ǉ�1;��"O���!mM
�䓢Ǐ����"O�+���u���
FF�%Q��*�"O��S�%�l`�I��G�0�d,�7"OP:7��E�LA�p��`�~l��"O&u�@%��i�0衤Ր�a�"Ov8��m�����c\�r��]�f"O��u�M�
	6�bg��s���Z�"O�582.�/s�ujvLH5u� [�"O(T�R��;�"q( ���ײ�y��W�RNxY򴏌�V���S��=�yBh�@{�8�7�Ż{�
9h��&�y�/&��ݩ�@́j�*�Y��	�y�/
6�b`�[�1yp(Qn��y�/���I�" �>��U��;�y��Dl���	�?d�@�	�DH+�y� .�:Xe�@�e�uH��޾�y�aАn�`�£lE3 ŐAL^�y҈��q�D}�	U���Y�K��yR�Nk(���Z&rp3�aɋ�y�[��(! <K�X�����y�΍�\�h+�l�� I�0/��y��^2>|����ͺ	r��@���y/��tl|��e�݈
�� ��2�yҮT�Va=J�AȑJ��)p  ��y�7[��}z#�
�%��:�y"��d[zX��K�x���Ÿ�yB�O-� p�W,r~�	ӑ���y��_�5[���FU�m�(̝�y
� \%�-�=p����a�?z%0�"O���@k=Dp��@��Z�j���"O^x�cNo-��fe��f��E"O�$�4�ݣC��xb�D[�x|",��"OX�H�J?aW�PS��X�c1"O�	b�MI$K�PQ	"e��tU(l{"O�9Q�` �h���MO�=�$"O
(*4�&\gH��NJ�Ղ�"O�E!�	#��it,Ё-X��R"O�uÀ*�9V�t��`�� a��	g"On!i�M�.ќ|�u%\.eT���0"O�u���2 6��'Wucʄ��"ON�샿vl�zTo�<WPtt��"O�rF
T��t�^,Pxx4`"O��r(�[�(aN��'Zt}�u"O�A$h�� h�,���9m�6�� "O���E՟#�<�0�}����P"O���wA��/(�x��ݑj�|PQ�"O���Űw]��iB�'N 0�"O��pm��:��Q,d���&"OR�ZC拿6uL i�`٘|�X�y0"O&��1�B�;����ca�8�����"Ob��'�G�R����1��*F"O��3&��(~5TԠū��|�%�v"O�\��B%7�s��H&a��W"O�gD]�2\x1��
�h����q"O4Jb��4�������.�t5�"Ob�BdʒP��R�c�8��""O��:��A�>o���U�S�R\���"O�Ti7�U/��J"���T pH��"O��Q�H
egZ*C	S�$�hY��"O&u��	�>�0��`�r	�(""O���0k��(�L�+!�T�X"O�2���.B����+�2^�Y�"O&]���Dds�K�J��@�"OH���R�pZ���Rߊ�#"O�I��@*F���z�iB����"O&EK�M�hW��;��H;$�{2"O�(h%JN2[�D�"U���5z�"Oi�qH�?7��+DG*6��1"Ov�{�ƚ�{�>p`�H��S�2�K�"O��k􈅡j��}+�	[)M�r�zU"O�L�Q���<x03�\�wӢA$"O,C�`�.�:Y��EW�fozx��"OP��"S**ȱ;���)Wh���"ON)�)����X�����	5�p�"Oh]J�D�.b1J@�O�5�+�y�<�5��)��D:,C�}R�!�5mw�<Qԯ��p��XU��A�D]�0eCF�<iE� �3i��7�H�Z�"j�B�<�G��R%n�z��YP޵:`�}�<a3MCq��ɀ�nS	U�$T���TQ�<��ʀ#��WO�p������GR�<��d�;yW
��-E�ܖs�`@N�<QD���]�<�y�F*:(��9%�FB�<Q�M7f��xʵ���9���Я�D�<�C長[�D8��(ם(nT<��	X�<rb$��)F,J`�Dي�/�s�<!�H�R�ݫ�"�3e(� ��]R�<��"�[=��'���P6��9 �p�<A��& ��jS�^^|a끅m�<ɷf��
��S��n#:�B�i�<�@�
��A�I%RK�Qׯn�<Ag�J�N��is6G�'����U�d�<� f�@5���K� s.ۛH< ��"OV *�h�'Sp���/Q�Oj���"O���!�!F�^YeCZ-����*OH�@2+V)#8%��'_�24R4�
�'a�̣���Z���X� ^�+êp�	�'�$�y"L��F8(�Q6(���A	�'��|�� ,I	1M�WzA��'�6p�5�W�&Gn�sf$A����'D6�g~�t9#/��w�Bٰ�'�^�2��3\�z�c#@G�Z1y�'
�<0���DYcϊf}�q*
�'6t�C �|o��R�X_d<`��'� �2hA'��`��l�=Q|�){	�'pF��j�w �P6�P�_�~!��'�T`�%
�\0��5��WA4���'��2��ÐI�:q�dǂÔ���'R���a����I$ċ�����',�|&�T}s�-C�{����'2��
��Lit��1m��lI�'�q{S&]�a����X8>��'_�eǟ�|����#�	i
�8R�'uX�Z�'Y�Y����k��di�'`�\;FeU�{J��ف �`lЂ	�'`2!R�a� k(	�p#Չ@�L�S	�'��Cʋ�5EV��cfEC��:�'U��&�&:�!�5�?�e�'$�[�h�-?����EV�ܡ�'��(�C�<:t6�c�M�v�S�'n��3U�6I@:Q���<90���'i`��.�c��12	|*�݊
�'��%�mM�\�8�!�� /�P�
�'�����o�;�r��c�V���Z
�'�8�bf#��p��"R
y�\���'
N��OۼN0�Qf�i�!��'�x-�F�\�t�
� ��q5^���'� ��Q��� ��@��m(�аr�'�
,ҡ��*6��aD�\�b���'WL�
���0��	���!C���M��^�{Ò\���՞bXC�ɀj�p�1�E?D<8cU �6��B�I�e�� DFʴx� �&e�&
f�,H,�2��'f�>�I�_?4)a��\�3�8���f�>p;�B�	)!$�Z��ݿ|�!�'��!"?�6�\���۷2�O~��%��94h����?3ۤ�W*[0T��cÖ�d+��d��,��<)��� ��ya��ŔBe� �k�M�<g �_�X�ɤfu��ZȀlZ7�����鍥*�& %<� ta�O�E`N?���<�4�D�������#\O(��W"_-8�6Y� ���:�D��B��@H��{T�3<߼5:'�U�->dY,O�t۶<�3}��֝gT��A�O�4�T P��8�'(0gM�x���b��B��f����q����las([�F����鈺]��@��0>�B#B�8��A��e�n�	PG�)/8:t��lQ ��;�@˧140b��.3�H�'h�I�6 �r��&�r���1
�'��x��j�6T�Ƥ��*� l��m�f��&}��P#�9�"0�6�\n��|�/Ot��`@;�aK޺\$���L�c�xT��Fr��8+�+~�qF�F�{�t���:N��h@�	D,=�tH�I
�}���Y�`��a%/�q��Q�1&�r��� �Nb�	�=Q� %4����O�2j��t�IX�f��T��!� 9b)�l��x�!��I�����'A^�	�mœ^�Bxz��.1$�͒r��X ѕ�D&4�0�CBX���W+�д��댉��$��J�%����T��-�P&��L)!�dB�š�)f��$Ql�"�V� !�2D�L��`.����4��7�T<��+�|�c��8��@���D�|���w�|���ط
��x%��ۣK�"qN��f�8V͌d�PNQ"!p�kBTX���=�#
,�Y.҈�%�� ]�%p�B7LҖ�E}M�[�FQ���B̧p�RA�c���W��s����t��S�? .�Y�-�458������Xv�O���a�Q�s�|�N��}���ѭ?�n<�5-Y�͚Ԋ�j�<y�]S��i�CCX�	N�LS%�f�Ć�{�X�&��0<)D���J��+�4���qň\8�,��#��q���
�;�&��)_!8�"]:%���>�3�\�6����'1x=p�䐃s9���ɱ0@ �Op@U�ǒac>��VI-׃@kܧ'�|
�K]Kl�B�\lɄȓ	�tHT�֒?Z<�y���E�����O�����3m���%�IM��ē`6�P����H܈Ȑ+�,��I�b0�PHͦ�.�i#�"e�,��f�[$���?�v�ϼ7�����H(Bl�A�'��x��I6{(�$>��0մtv���J{3*���:D�x��#ӰoS|�p�dݟP6�VC�<��#őspZ�@ ;}��	�x�9q C�p�qR �y�!��(�6a{"GN9*̒��v+*��O�1փ�"�X��qO����-~�pZ3�V49 �YQ1�'��4�̸D����m��@0v@�8!ؤT�h؟dj��>ieʕ ���@�X$���;�r���'�T�� �s�,[#���Ԡ+ff%��"�	���\4�y���B���b�O���6舀���<o4� LP�R��r�1ڧ
�I[¥���X��]-
���ȓM�dI�O�	e'�P�b�/S���Č��(�@f�'-��"5��^�g�	�I"��;aO��F��AE��
jB�I;#c�}˲��3��m�0Ba� ��ܶ/�^#�ا��=��#��F��
1���2�i�}���8#/-5���릳i��|��(	�0�`�ߞSe�	�	�'��Ig1=��A�g�CB�`�Bȃ� ��#�N~�O�|Y	 �X�|�Fl�a?�q��',tU1�/�9c|���K_4X&R������*$�c�'}�<#fڇ��[d%"K����'0D���MF���ܡڶ:�������O`�`�OO9�}�ۓ>��.[�ިzvi�0����ɪf�z��w��?���C8 ���
�GB:f���cU�y�Ƣs�y���!S#ԠI�%���O��S����G�}���,S�N0��N(r({��N�<�#EN�l���8��U�7B�=S�Lqс�v�S��?rAٍ
���x�R##��q�Ҡ�j�<)�M�p0q铀V�g��0�%)Gm�<���+a�~����~0����@d�<Q�N�-I>���o�0~V��RA]�<�qB�
U�Z�E�RT��D	Q��T�<���ݞf<��ZǏ�s����D�<I���X���A����2�B�<��b֔x{�eH�
�*=�(i��q�<�u_q�4mr!.�'_�y��
m�<a��_�:��T�� *#LcS�b�<qf, �;\��C��`��fK�V�<)� �4~�T�c��T�)�Ҙ`)�D�<�$�כ<34ش�S	z6��"�X|�<qV�ͅ��U� p�E`]s�<AT��&w�R���etNN���e�{�<)�4oP�ݩ���uL�[DDr�<Q�GN�\��в�é'�VX�2�Jl�<���<Z�t��V�32��n�<ab=2�>�0���+I�6|a���k�<ɕD��Z�����h�-�VA�a�<Yj�m	"�[��̞,g(|1�T�<yAh̙6���`�9�bY�rL�W�<��b�1"kr!�?;Ӷ��Q�<��c��4�w@��(�z��φU�<��M>q-���� ؍�P ���S�<9����YСC�O/3�E(1��w�<it�E�*�Nɪ��A�̉��@�p�<��e�,��L���<0z�z�&o�<� "�!ST<@QϜ!op�͈U"OL, ̊�(db�!0MU#X҈{�"O��*G�B��P�mN	 .��"O}���B� ����m�(u"O�P�� �bX !Q�B>�p��"O�4xQ듶B�y�8$U�"O�UK@萤RP��¡�J(n&���"O&�yd�4\rYqUZ�,U�ɋ�"O������q�R`Ք@؅)�"Od�[q�Gc��a�J߬UH�8�"Ot��\l���r6��K�^�#�"O����Z�'@>0q��U�wv��"O�l�7�A�N��P�3eg$`*b"O�$��mǾ`�
3փE>V��"Ob!R�m�=,��\1��ߋs�88�U"O�	���I��Db����x���5"Ovd*��R�w;����R�<�6x�C"O�ݳ ��&�n�cH�ki��Xc"OM����8$59�fɱDA��@�"Of4` �_�^�Ҩ���>l7��R�"Od�T.X|�X�صy"�Ls�"O`h��i�G�N��#nك: ��N�<��dÑ��m�L�:
�1 e�B�<	n�h��= #�W� �DQ�lK�<y�h��%/6����qj��@�G�<��q �)G'	�3�LMA�<�bЬBv�$�#Ļ)Y����l�A�<�g!V�o1��[%�
�KiB�R���A�<����go��0"Iޮ>����Jy�<1)N=#�69P��96f�҄�s�<	G�̣0s�<�Q���j�f]��s�<���
\�RAR`E�9)��q���e�<i�#ήDkH�!�K-u���c#�c�<�cbܯ=M�Y���0U4,���-D���vaW�݆�N�9�n��z��B�	i+��R� �?.�P�`�1�L�FBJ�r l���&	������n�f��e��{Y��M	jW!�d]4nP	:�쁖af(0Q�&�7tO!�E�b���Xt(N�H��P*���qc!�۰Z�������Ƞ1@�NY98W!�G�P!E�F�t��B�+��P!�䘻n�t�q�M�Ts���'�+J��z�՝��a�p����!��A��_�SԪ���H���iUs�>��'^�Gbl4V�V��kn��������O�XIe���hC�H[<<�5C���V�$�o��$h��)��	b�S�,���R�#Lo������&GK�5[�'�qZ���%�>)z2�Ory�+�.�  ��I��Y�X;��>�J����\�������<E��Ǝ�-w��8fE�B:�h �A Un��2G��aR�- ��<E���X�5�͑i�6K>܉�SFLm��zS ����0�a��.҈y x����ŐԂ�� A�*��'� ?�EI�4�q������0�\0O����,c�^���O��m��&n)>|�.�M�O����B��a�r-�mY�	��A	�+�� � .[�Uc�i������M�O]��Ww�My��A,cC*5!R��
T�0�Z5g{Ӕ-�%�H�$@�r����H���J�,���S͔
�Z����]����ri�	3�D�$����S�RNh٨�@��/�0����S:%<д��L�ɦvNp��g�)�$N�9� 򁉀�7�P9Pw(����5�X)p7�����	 ���������5_����婌SJ��Ѓ����/F.Ma��rE�`xݥ���OwV�3c���%�Ԩ�Be�uY�F�S~r)Q�-�����|��i�z�j�W�*X?\$��b9z7�$�<r�t���C%|O� ��Q�8��4b�;8E�\`c"OR!e��������3v:�Q��"O���w   ��   �	  �  �  �   (  1  �;  �F  R  J]  6h  /t  l  ��  ��  S�  �  b�  s�  G�  ��  ��  �  R�  ��  ��  8�  y�  ��  k�  � 5	 z � ? �" ) N/ �5 �; nB �H .O �U r\ �b m 6u z{ � p� �� <� �� ��  x�y�C˸��%�RhO5d��p��'l�I�By��@0�'�F��L��|�t���pd��46��-zw�G$�`�	�A��{g�cY�.rA��͇A�BY�G����u�蕦f`�T��V3�$��06��	��d�<x�-c��3d�v=Y�	9mC�����UF}s��^t��֝CB���M�FH�z�e����В.Xe\�����.2H¥В&|ت�)Z��7��	�:���Ot���O.���4r���Z�*�X�#d�څ'P8��O���O
˓����O���O����\�Q�x�tc�#2&���O
��5�$��o2�d��6����?R%�Ȇo ��;�'Y�b�F����d�<�Ф�dAvZ�`�*r��1�Kǟ|���X:�8P�@&ϣ\@u�O9)"0�_#{�(�h�e���������~?�A�!�O$���O��D�Oʓ�?���D��#�$�J��߂��1x�k���?���i)�7m����K�Od�nZ<�?�ߴC��	�jf��E+G+cې\���\�)8,�@��$&���^"̆�Jk {�QY�'��<q7&P+Bt��@�����ⵓ���O�=E�	��=��=p��	�=)�SKհyV�Im�� �B�C���w#��r��L Wk(����8�Ӈ4��u8CMK�AZR%h�-1R���<�S�O���r��C�]���#g�$�%�G�ay�L�c�"7m�d�D�
R^�����th����1U4��<Y���?ћO,,����'���x7i\�\0�����9�\|
�h�*�<¤�.���q��۱=�H��G+PM�dq���O���-?鳫�f	�+`�.;X|��̟T�'�ў�>��EIJ�}~L���_^��h�/$�O����j���J�D��M ��nU��"�d9�ɻ<*�"|��'}!*��!Mk�i���S�Đ(��?Q�Jĥ�6�F�a���ȕ�Y�ks�i�ȓr�>]��J��U���Kd�م�N�`�j��ȕu�v4P�흢m�H���_��"�'E�H�y�2�\��� D�d#�疄m�$
��{�h�@�F�3���	�2]�#<ͧ�?�����קI��,B�'G�%L �`���PyR헴=�Ȍ����4��H3E�ų�y�g��-(��V��5C��#����yRF�0J\mP��� +�C��%�y"��/6�<=y��b,�)�'�.��P��(����r	�1�R�{��	�dy�X@�_�8����d�	z�)����QR�+��RL�B���)b�C�I�	��R�͟
2�V})�.��c�C䉄2����t "jr89�n� i�C䉩k�P��)K7"Fع,�?ON�C�Ir/Ԥ"��B]�Y���Ȉs̓O��>i6Í��V�'��BҼ)HJ�ӧm�'�z�{�J4��U����̟\ϧs�6�rܴ��'�n	��bH8	��Ip��	��0��
Ó7/ �y��C�/����07����ϻ�0<q�dL���޴p`�f�'/`R%��$�b0�$�I�D�ĸ!U�D�	K�S�O��-�(ф_��1Q(����2
��\2�'9#!�t�c��I��QL���?	)O�h�dJE1:�Z�?�	ʟ᱀�4+�P�1#��P�VM�!����I: ,F�qO>Q���ϋ0��3�MA1
p��ꑇ??�5#W�Tq�"|��́[Z����@'=��T��}~")���?����ϘO�X	ZFdN�#zl����*Ⱥ̹M>���0=y�F^mq��F�YT�,�B�i�'���}z�H�3vpA��"�;>D%�2�(�Mӄ)��?i�2|J �'����?�+O��+@M�)/�(�q�şݼH�S�$�	�&�Z���Dd��@�S��D�B��g1O���q�'p�,B7�܍_d�HÕ"˞$|�t����DŖ=�r��'�剻[X�%�ͳ/�=RC��^t̅ȓ-(ȴ��`��^��ze��>���'��"=ͧ�?y.O�1��,�;"'��q#Q2e��*��HR��d�O���O��O�'=˰uX�n@�B�zՀ�B!Ng6dK���q<a6�M�W���
sc�4������͝0�L���T���"����w��C@ܙ}�ĭ�wO��<s�~b��aA��Y��;!#�Pd�!�ȓ�I��@�8�h�냇�8\��'� ܴ���Lt2X���I78�u"�$\y�鋧�F�G���Icyb�' ��'����Y�I�<!��'��� ��Y�i�2
Vf��k�1V{�x��'0D�!q�S�e�j!�I�d������)��R�m�5LU�v��D���ɷ0dJ���O�	o���ā�G�5�������%&��\�ũ�y"�'��OQ>	y���9N8�U����\\�qZ`�>�O�mZ�R�
()S����I��ɒ%�ܠ��Jyk�3�6͂<���|��'�*��3w fi�s�_Lp�?y�0�.����5+��H��?	+�B�'G���Q��V�%��������� �O~���]	 x���B`R�$���Phqԓ����N ˂�K�.\�8��9�5�� ���O���N����Is�O�,�� KC��i�2ǘC-`͐H>Q��0=���;�DE���	�C��Q���KB�':6��O|�O�Kgؤ���(%�B�1�!���`�m���\�Io�|���?���ɟ$�'�4iaA�~H�d@�"aG��ZT��O:�p=A�!��aw���_;�S�[̓`����Dt^��4O�(
,��Ӹ,6���H2G�Orb>�d�O`�P��8�/�^��!dN�sK\B�ɇ[|>ĩVL�0%�prE
	��%U�|���4���/?�IAO �);�]�����]AyRC�	���'ɧ�O��q�cn\3c,�Mca�KJj���'=�0 �	uq�Y9��9;�����'-�\�� &ee^u���^A��b�'��؀�y>�j1k�Pt�}S�'xX�)U�0?0 ��F��$C�h@O>I��I�{���I�?���&�9	\M�2LХ]���3�d�O`�?�'��D�b@!Wa�, %��8-��eQ�'�u0���0����DBW� �''��8bC�!~B҄p$J!O����'π����0B
�,H�(�t%���E0�iЗ%m��r�l��:g���d�hO���oLpL�v/QJ����5儒XS(���̟���I&=5�qѧ�N.Ѝ��Z�1�B�I6�ܡ���Xh�f8F���rB䉯\i��a�.2����]��C�	�yũ�U�G�"U�����\*�?����0pi��I�B7_��Y�$[�,���dQ"[���ş`�Ir~r@��zSr���D�	C���F@
�yN�<��TҲ��d�%� 	�y��ܫND��HĨ�.�p�@��y�%ƔN��y���E�9����	"�y���6��Y��6�f��d���^h��(�l@M2���T�=�0I�S��K�`ٟt��K�)��6떌��Rs¸�aGC�XZC�	�gt�u���Q%+�A�A���,C�I��Z���C�X�Ԏ�C�		,�T��Z��UPƍ\9`�C䉑UK6)3�Y�[Yv��F0"��O�|E~��G��~Rj�?��%固<B��f�	�?qK>�������	+��4�D�<jzh�E˶dZB��u�]� �	�H;��4(ʘOa�C�	������1[�n�Iw��=j�C��9 �� v�ĭjJX��cE�r����Ɵ��c���7��a���g�C6ړ'T�F�TK����`i�eߝD�hH��A��2�'Ha~2�P2 |����Nl�zy�qk[2�ybD����AS:hD^�����y�IH$VX�;�$	$u6b�) b��y�a�p�*(��!A�<kT@k6ƃ���O<LE��-�")� �B�_
-�n�����?i5a�o�����':2������M��AQ� H0_��	�u�.D�|K.O�.\:�w�X�n�B�
�+D�H �L�6�@GڍW���:'D�d��MC�%�ޕ���
�䠑%D���m
2���1,�*G�ր���<1��)ʧ/�i�)��k��|��bW�U�'}Pd1��'R�|���h�*�x �BOW?0�rl1S
Q�y
� 8LHcW�C�4�7�P���]�E���	iB$Q�`�%����8��z7	�5ba�i>bf���r.Bt��m�!P�6�AA'��R%%�D���X�/V���$EX��r�R�^Yr�����U���|��'���z�\pw�L!|&�-yQaM�,�.Y�ȓ�<����M�#_�`� !���5�ȓ5~�-f��@�-�R���7≇�"�U���ԈYd	. i�<��	��?	4A_x�nt�É�?3]��Ed�'o��+���Ɓ�[�B��B�+˴;T���O���d�(=5^Ē���g��"�ɏ3U!�Ġ_U6|���Q��� ��7?!�ϗg�ށ"�A�9���O�%eP!���7qPB`#I;��`��Sџ����	��d�P�����^�d�?N2A�:�O��O^��,?!fe��E���#Ȓ0I4��i�P�<������
�KT\PIC�SL�<!���]qj��͟� :j�p��D�<�q��
��ds�`L4z��:� \~�<�ŉV�P�kV��*:�޴4�xyA&�S�O+@����8r���`�.O�3�G�O<�9��)cs��"f�R�x�{�,H<T�!�d�i�z͹v��#_����+�d!���7F���ί��\�i��!��P-b���Zi@�[�E�!��\�	p*�<�� ��|3�'|�"?��c�A?���֎R߾͂�M-�+��̟�$����T�g����(��gQ
	�s��4@�!�/U9 �4D��Tfh���!�
�Z�fx�EKO;qR��r��.3!�䎣w9Ha�AP�YFތ!������Ob1j%�7g`�:q���6G6p����'s�"~����7�Uӕd�0:��4HY
�?y��0?9bn�Y).l��F�Mr�aU�<��/p�j�s�O����Y�$�Q�<�VO˖>o �Ԉ(PF��D�J�<�O߉�(qj䈎 '�>�$XF�'؈�}�0��8�<p+s�S1�5P� �؟dz4!<��|����?��O:<��� �?l�Y׆�i���!e"O��`�h�!ڮ(�� Bv�rmȣ"O6LK)�h�� �R�z��̉4"O�� ���I.]��,JU� �5�!�䓥T��{��X(=��IA��n)�I0�HOQ>�*���mUL,R��M���P{�ɤ<�F�V1�?I���Sܧ6����.	4�D,������=���δ��Hq� ȃ��E���VfȀ��W�R���d$`�b[�'���c�`	fMd�Ɇ��!AV)r�'�^�p '[�R�c�m�w �ĂJ>��	�����
:�&���G��,� Z8���d0�$�O0�?�'�0�An��T{��rTH��L��$��;D:�	B.�p;Lu��#^V|��Z@���΋�}R4聀jƠ���9h�ph�`Z�^�T1�T'gQ��Ɋ�?��GA�w��t�SA�?�B�Y�[[�'�����	��x�J�@*�-[L&a8A@
�f'h���O���d_�Ln] \��i�R;B��;"O6��ԣ>'(�k��6:����0"O �۠)X�gd�q��<X\j "Oh��G*�������K*�%���h������~G������K?~\��'@nD��4���d�O^�+�е�%��G|Z�Z�.�p�nчȓhB��������82ǂ˾lќ��S�? R����֯G�d@bGٹ*�R�"OB���O.�t,��Gь�Lxc"O�MzG�-Ab\�"d7Y�+�Y��s����A�Đ�5n�9QFPr�N�0H$�B'���?�L>�}
�P,\�d5ʢa�lSL��A�Q�<Aĩ]��Y�LR�Q�x��mL�<�W�X�N�T�5�CC�2�¦�~�<�P�� |I�2��3ӕw�ټ?�!��!F.X�p�=Sb���F�
��'��#?)�L�z?��%�2v�t,j���z�P����̟l'�T��T�g���'~� e�s���[q�D;_�!�dɚ{�\��(k��Y�B�82�!�D@�ŘW��-mjM���0_!�;�����	�5^��%�\un���OJ�BB =�R�M��ar��	%mx#~*э��_d܄��F�O��9�ů�?���0?�bY�D�	��\��$��O�<9d��&Y�
2&� [�\܀���H�<�i�\�HC�&^�if�i�!��F�<�"�$}��$פ�v�Jm�&L�'l
�}��E�0m��:�덦c��Г�ş��&i6��|R��?��O�D�J�nݐT�h!�z<�"O!��H�]<�`�b���o7�p�"O���Yκ|
E$�QzMS�"O�h��)��HhP|b��
v�Ԣ�"Oju��,d�f�BP#�}n��s�Z��a����7�p1W�W�T��]Ȑ�I�4=&˓ �x����?L>�}��H�?��8:"M8X��!�˅Y�<�3N
+�^�CC�1%X(�@��y�<9��%s�8hk4m445^��Us�<�uÞ;X��-QWC�W�F0`�q�<A�f�:PptzP�Hm:���hMX򉫒�O��C�O����G[L�A3f ��A>��'i�'@��>���?��1�6�	3l���@�<��F39�n��r�+&^<͊���{�<AqF����ш�]��+� �ȓ+���	ʏMH�p��n%�N����?	��_�%�V�󠡔�wG�R��O]�'�����	�6>�*b�׽CŃ�	
�NS����O\��DT[E�|���KK��d�$�>�!��7|B ��f���h"P��M�d�!�Dھ��a��^�Lj@A�`͗)�!�䔫$�}@���WR,,{B,�z;џ�؋��K�)¬�'Y,@*Ȧ��$�����O���O@�D+?�Tf �:Q�t�	��p�����iSl�<���P�0"4�t�[j���G�k�<i㋙$t`��N|�`��$�^e�<�#k�!])xcb��d����Hj�<yR�^�r�j�(!�;>�n0Af��Py�M;�S�O�8u�À�.r��n�*2/O�5"���O��>��i�Q*�;Q@[6q�n�I�ď�y�!����8%�ȱfB>��@γ]�!�	7ð������/8a����$ !�X�"���"!<	L�3`��k!�d�v�bL�ݶZ���AS�1�'(�#?!WF g?Q"H�)v����ዎx�	��IMܟ�&��ID�g�Ď*��$I�Iֲ��Q�HW�!��Y�o��ܡ�G>*v��%�:�!���O�,Eq��S�0�=ѰJK�i�!�$H30R̠��(h�䩜,��b��O�8*�E�\ԓe,��.8ٔ퉙Yq�#~�B�^H��]���3�L-I���?����0?AB�W�5�j!%�ȉnI"Â�U�<)�kŲCV���gW;2dq�E�R�<� &")�$ܼA�M��<J�� �"O.���DT�\x��:���-"D���0�I��h���B��J5P�m	0l	:ET�	 !�'sR����4��d�O��@d��3�Q) �B5i4!�4�Ї�F�|(7'ېdIF��G[G2��ȓO
���"��8� �����F1��i�=��m�-j����O�1���ȓ^^2�gG�u���F#Ғvŗ'�("=E�t�)w:��OA*5��D�@M���πzV����OޒOq�D���	z�l�a��|� @�"O�|[��R8bQI��@74�n��p"O4y�e�F�t3�<{�K�Df��[�"O8A�,��s��X�R�D�>I�a"O�]h �P�E^x��J�i�Xj$�|B�"�r����8�E��i��E�xE�'��
|���I@��ʟ`��ON�	�!��Bh����Z�5����"Ou�&f�[�� IX&Z9``��y�NS:R��;���r�	Ip(��yR��'g�:p�Ы8�����˟���?��'_�AE,��$F5�BĩH�$
�����?�
ѩ����S���R��i����x��ȳB��;��A��G�zݼЈ��*D�Đ��sT�z��#.����%�'D�TPׇ�7+�}��jP�5�o1D��{���Lޜ2Ze�9��J%���>���)�
�T��W4$�zkg��O�Q+��i>��	����'dLK�!�F����^����B�'ӐA�핃2���Ӥb��E�B|�<��e�x�8i"�B"4ڢX���~�<ɲeN�WL�:�lL�T���i�j�A�<I@�-�d���X߼H9�nRyb�5�S�O�(�у_?X ����Y�rN&ղb�'4���c��p�ܴ1�i`���?������J�i&i02��5qh����$�O����O"h���Ϭ$N^�[� :G9@��*b>�!��7�x�ڰh���>pq��+����" ܔl;�)�$_�`���qrT�rD.Z#ɤ��3���bz">AN�ʟ�	q̧!��59���Z�Α�Gɂ���'`r�'�t��1ꖰg,A�!ϩ֔t��|)�I��L�#���l�¡�h m���A�\|#��i�v�X��'>�O�D�'m�pz"�D�v���Y���N��M��'���D�ׁUP0��V�ѯqS>�s!Q>��|�C��Hh�(87�d�$J��A�<	v��D��q�l �"�Z ���'��ށyu��o�N�2%���.(�}�T����O��S�Su~�
V�?,A8F�Ùs�b�3�@��y���8�bq5F]�T�.5�U-]��hOXG��<v>��"!�c�
5�b*^�7��4��'�E�?��7����D�OXʓ�?��B��T�T�S�U/%rȨ(g'�?"N,�8��'�=+��E��
ɟ�T1��&��xk�@ˌ
��u�̼�I#yj|I�b�q��g�'���]�J��K0l�|lA�+X~~2���?I��?���<��i�"䃎%]��s�j��)g�� "O��(��W�lDQ��j>J�T���'�"=�'�?)/O�A�� �M�`�+˔mތ�;��Q1:�L�n�l������p�'Zf�v9�,]p��ٽ^qF�hJ'_-z�SP�A�DMD�)���5�l�SFdaX��#p�@*JQ���V�B$�xdЩE]fp�'�y���Y7g�˰<�l�؂/1s�^PA6#�a>���f؟��IT��h�@����8y�5X�JVQؼ�Dm*D��B%��^���q��L������<	Ѹif��z�Z�B�z����$ 8���W,:~l%�<�I��,���6E�4��
��#�6��ՋK�0�C�I
2a���N'ĝC@�ˤ��B�kJ�{`���U��ݸ�.H+D�vC�	�����a%`����1[t���dGNy���+�m{A%��F�H-������'?�l��4�����e��Zp�"s��3�

C��D3����L1��z�Ы5ؑ�uf>D����iH�b�����`ʡ7A�a�qF"D�� ���dm J��]H!%�A��"O��sdH�rx�$��3���x���ԐbpG�9j9��(�dAZ�2�s�Җ�Op���O��+����C%�T�J�i��T�?O�B�ɏZ���q�^�h`E��!����j\��r��O9J��)� �?�!�d5���sL1�'�λo�!�䋀@�B|�D/<5
��v�ҜN�"�;�S�O�
y:4�
�MiF(i�I
X����'\V#��'���|��)�8r��5�r�Z�I�n2���WY!�
�0���7V(H�s�D�G?!�d�6Jv���B�Bŋ�,K!�DY�J^,d	ìT;�J7�	,/!���$�J�r�� 2*t��SNM�,+� ��'�lI�'ՊpSL?}�G/�*b�.�:Q�ޫQ`4���O��V�A�4��4����UiJ�V-�Z�k�3T����	D���`���<$2�{`�@��.U;b��( ��=$����OJ��4�֣s8Q)*2�n� ���Oz�!�)�[v��D,S�=S��d����	�`q�	�V�xI{ЄN$9�QK�I>ddʓ�?a��?���4��ԛ��&:�x�R�=3dNld$O2��0�ia3cT��>�c#Q�0`��5�IǦ�$�����&98��,5��Ax&�[���	�~��[>���|�I�6m�q�IW�ta�	��xP���]��DT�&��=��O��Z��U� �z�ɀ�_�ao���@N^���k?���9OH�����./�������n�
�l��l�!4�e�@�OZ��O,T�k$�Z�ZP��@nl����4Gb��O�舡�S�Z�`�k�
͍(�ڀ�7�V6��	�b�.�'���'2�0�L���4`�^ѣ� ڇ|Cb����xh�<�'�qJ�(�����'ڌ�h�o���3�%���F�(��O�s���W�/?!@ S yD~-#��\�P��is�J��a+�<�Yv~B/	f�O��RGԯ[�$�D+� ���� {���&]���S��'O�1��'���Z#�E�D�4�P���g�A�7�v��$f���gU�W>� CkY�!�ċ'oU���ɛ�g�27 6{y���'�\��˫�$ʧ��i��0�B�~ Պ���}ID���4�?�H>��U?c��s�4�?g],+p��z�z�[R�x��)�S��� �ʃ�5����8��C��V	�`��Kǻh�
�;����(�LC�	�<{��Bh�pঽ�n�� �C�@a	�QG�TT��З�V�l$B�	8�V�+'���`���4P�B�	�_��x`��;<L�{d1ZFB�I�@I,�35 �jge��`. B�I?���R"קU�2���)X��B��>/'�8�FlM�k��[�O���B�ɳO ��t�5(��yr%-Aej"?q���?1���?I��$��+chT�����Q.N?	)�(�D�in�'�r�'���'���'��'�9r���qTՂ�BX��b����O��D�O���O���O2�d�O��Y�>S���F��@9���+�æ-�	ܟ��Iҟ���埼��֟��	՟D§̊;,:�r�ڮs t
��>�M+���?���?��?A���?��?��%�� `�$��FL��i֍@˛��'���'2��'"��'���'O@��}��Ec�`r� e��3wJ6��O(���O����O��D�OP��O��D����.��:}B`mTN��l�����<��П����T�����ɿ{7$ذ���}Ѩ���醐H��5a�4�?a��?���?i��?���?�(��!�H\��y�h��C�pir��i���'���'���'"��'2�'=��BC� f-���CS�^�}�2�r�^��Ox���O0�D�O.�$�O����O*qh�M�2Ԁ�ׂ[��0�b�e�̦��I�l�Iǟ �	��h����I��[H
I��#`�H5v��ء��M��?���?I��?����?���?�ڴ`�^ɢ�e�%���L	1(��7-+?������5�-G������>����*Q�5�<�[�O^˓�?9����lӖ牚h&~u� ��ڬrR��? Ѷ���O�Ij}���4ժ̛��O�K�!��V&�����X5��r�'���PQ�i>�͓P�lhyᯘ*�0��9XP���Vy��|��/�Sݟ\� 8��#Tsp�W���U��(A��X}}"�'32O��'j2j��u���!J��
wA�
���'F�c[��*<0�O�6�?q`�|��V�Wd��&���J�Jb��<�-OH��9�g?��Eۦ���n�2���`w"]����O�[\������vyA&(�|zDE���FI8 ���O��D�O���s˸7�1?ɚO�F�)y������8gƚ��S�̇IU��G�9ړ�?�-O�b>��d�<%N�1��S;����*�<9�S���'���	]�����%��Zy^�+���S���'���'���=ҧ���k@�1]N�X��"%�QA���M���'F�
۟�%�|�\��AE-ǄD�p�q6�M�����J�V���{�O��D7$�`�x�0A(X�t����Ѧ��?)�T���	馅���v>����>l\���CG�R�h=���^���͓�?yU�-"�r�����d����]�1x05ۦbA�V�\Y�"� F*��$�O����O���O��*�'\}�D�/1Z\aX�lCw�������������<���i81O����Q�D�.� Ó�_����-���O�7��� AA��j���zoN�h�S9�^"g�2Z�R���vC0��������OJ]��JI/����`�\b`�p��Hw}��'���'g��J$ř�%���&#a-_����E��I�8�Id�)���3.H�S��,~�b�1%d�V0�FC��M�E_�,���5��?�$ƀLR������gQ��q�� �>�r��$�ԟ�#�ƅ�|�x����8XT��OX���O�l�T�f���McU/� vµx�,�>cLP�v�óP���.b�t(���|Ӵ�u������FP�ΟD�z�X����7\��<�7�'H����I���������d���C3n�d�c�7I�Ic��J{���ޟL�	�H'?�ɩ�M��'=���`d��=i�� �B�I���ǳi>�6mZ�p�ӎv8�l�i?9j�!X����HC�N8���ß�"�=>���c��|y�O:���p5\b�"5��(�Eb��'~2�'��	��D�O�d�O
� ��ܦD\�P�%�yɦ?�	�����O�d?���3Mص���O�B9JDM_<�˓���g	�3�M��O�i�%�~�=OP�Pd���ϦY���<,X!Z��'R�'�b�'��>��*Exu!U��2T�A�X�Ά}�	����O@�S֦��?���>OL�Rd�Ħ2��SԨG?4�@��e��V�}�=nZ�:�lm�n~��ѩ0`nL��Z�M�0b��W�>�
�a��r�dbĐ|�Q�4��ğ���ʟ��Iϟ��Ʉ,�P�SDRi�B�QdyZv�I֟X�	Ɵ$?]Γ��PW+����A �<p�B���O<5lZ��M�'�x��ԉ�������Ѓ�`��	M�A�L ���������u��O�?'8�R�n�:P�p��
�7}[��K��?���?q���?a+O8��'��䕰y$��(��Ωw�*a�#h�@��$iӠ⟼ �O��D�O��	.ip��B�$ԛ�ML�h͔�Z��c�"�1i�5+��#�'�y7L�:Gh|uH�'ʋq�j(;u����?y���?����?a���?ь�I�?dul��TcW3M�$
>��ϟ�A�O��Mk�yB��u=.�s�m�%��x1m߉�䓅?��?Ԫ�3�M�'o�$�@��h�,A�]�� ��Bq� (@?!L>!,O���O���OTC.�6{�ZEc�%A�����O��d�<q_���˟���r�tgB?)8��D^�@kc�5���VSyr�'v���#��?1 $�BOh����R�Ԅ��=A0	�c��i ���?Apb�'�@�$�T V��9k�A �O�;R�s���4�Iß����h'?��'�(�F8r�Z���>
���q�ں�2Q�pX�4��'���?��+׬_��@J#���Zt�L!�OX)�?���=[���ܴ����V@23Ĥ?1�O�4�3��=v���d�ιr��l������OJ�D�O
�$�O���?*q�ë]�X�A'�;$I�m��Ɨ�����O����O|��������̓�ͭ�K�,���J:B&�A{��`�&�m1�ē��'/��Qݴ�~B!K>9�]���X�`"�QH�I��?��M%�������d�O���͎fpl��O�|���u�Ԟt����O���Ot� K�I�������yULM�VɖͰ��e{�L+��K�l��I���Id�It!�9�W�\&-��Ј��C��Ж'��dz��=ԛ����_��v�\�N]}�Xi$��m�i���ON�D�Ot���Ọ}J�'NRd���Z�ˏ0s�> �ņ�ٟ�2�O��$�O�l�j���Ru���)P咳Hx:	Z�BP��?��iK�6�ަQ��j�ܦq��?���`]�(��NR�4 �%� Z� 9k�hБCI ����<�$�<1���?a���?a��?��k�Vw
8����97 U �`�����n}r�'�r�'���~b�$9��ܩ��ڮ3�=�M�_��Iퟜ��E�i>]��ӟ�A`���SS�P3%gK�u-Qq���}$h\lW~R�A(����������8�@T�3J���4�"�dĞ���O����O����O.ʓ>�����L� Z0Ps�T,LN,�Ѥ@�����=OV7- �	����O���z��:�)JO��s��[�$�{G��|��6-1?��/%s�ȣ|Z�wl�)�*$G�:����Y E%p���?����?����?�����J-C����z4eQ��.'�&]R��'�R�'�듭��r�6b�PЪ�%
~Ѕ�'C �[�&��O����O�u�x�F�H���b�?7G@Y##�V�<�:�LD$+(��IY�	Ty�O���'mB�V5Vy��b��Zm����@�C6B�'��ɣ����Oz�$�OH�_��az�H۩��i	�⇲Ԟ(�'���u.���w� 9$��Ot"��M+d�H�T���!Eg� B'�E&w~r�O�J��n��'�Rh�aƦs�иxF�p�h�٧�',��'���'u�O��I��?���@<8N�eB�A�	��Q�([ڟȗ'�<6�3�I���$�ݦI��B=p��1`�jK��\L��+���M��i���)!�i ���p��ap��O݉O�>�c���8�Q �Y�L�`�����O����O��D�O��D8��h��>�0B%��N�RюE����O2��Oƒ����ɦ�͓(v�Q��\ ,�2P����06�����$�J<1J~���˩�M;�'����A9h�e*`O E�@��+��F��O�ZL>!.O��O �K�����ͨ�ոD�(��Gd�OZ��O��$�<iDW���I���I�X\L̐�ضgin�h�`�/b����?��\�L��Ο�`O<���Ǖ� x��D�=�BUS���V\�(]�HS�K��i>���'����Op��p��_� �ZE�'(׷/�0q��˟�������Z�O}��Z�6D
��Z�P>�a�̈́�S��>1���?1��id�O���:%,�!OY���Ǆ�_�
���O����O :��r��Ӻ��'Ź����F�R���ڀ�
Nk��SH�i��'j������I��	���	.&���A�ܫ����#N(I�깖'����?a���?9M~j�'��1�C�_s�����IC`aPZ���	�m
J>%?"E�:$�h]��gԾ7�z9SO�`t�BRK7?	rƍ�3����.�䓰��"C.�@��(b4H @�@L�!t��d�O���O����O�P�	ߟ0��a�#PnL�@�&!0D�eY�
t�$jݴ��'�@��?��Bb�Lv�Z)���&��A��b�T"����4���ދdv���'ѸO��.�888k@Y�va�A����%H>��'I��'�B�'p���,T������@���!��91%j�D�O���KO}b�'�b%Ӹb����]
J�H}�F�D�-���8�E�`��������?Iئ��)�'I1¤�ؤp2`��`�ӀW�DA�
�<IF�Q��>��'@�i>��I��$�ɞ+%4�L��G	��'��2;\-�	ܟ��'�\듹?Q��?QΟ>P �	*w1t����'&��`W��p(O���c�.�$��'Pc*	i'Î�mb� ��+�)PZP���
g%�����+?9���D�D̗�� JBG����{f|�k���?����?!���'��ԟP�DG��ȼ�u��TL"5RԈ�Or��Mˌ��>!�i��u���#,�d
� �P]���z�.�mZ ]JX\�Ig.`��0�0|�7���)��M2�ҺR�t�@�'������	��X������k��˹&}�I�E
 eˌ���(X���I� �	ן$?牗�M{�'� 1�" ^�*�vF�&���!���?�M>!M~�%A�!�M�'R�e �5Sa���$���*I��PL\3����$����D�'��ȓ��Y�U�l��/]�vx��f�'���'��T����OV���O��$�+��#e�\�}OXhcn��p�O�oZ)�Ms��x�,Q� |4� �)5���2cA0�@>�,��BI���$?I���'��)̓Z��i��h&R��q����<"~������	�����}�O��$�|?��	��.H��Q:D���>y)O��o�G���� �NʼqA)�'P6䈆�HL���Or��O�H�!�s�@�	9n�#Cš~���Q6R���+�����X@�e�IDyr�'`�'02�'�¥�I�d��IЯb��0xd�ƝTs�/����O����O0���� #\�
!X��<�i�H�}��'@��'Nɧ���'�ЗG�X��ԉ��h����u��k>|�2�i��	50�i�e�O8�O:ʓN�*F��ژ�ĝ/{�z�����?���?Y���?	+O�e�'2bFD�3m֡"F�,E���(P��|��⟐Y�O|�D�O払��]qAɔ-ھખ�ܓ\���%�|�4�rO�pqe#ʧ�yA�w��hp⍖}J���SmO��?q��?9���?	��?���i�r�� �m��:�B9�gZP�R�'��.�>i,O��mZ{̓c5�z��@7z��耗fI8Ĺ$���	⟔���\���o�P~b��B��q�Ā*�m�{�@4�P��P?�H>�(O���O��$�O�-Q���-m��H�#�\�Cl�l�D��OR���<�\���	П��IX����[����=o��9�o���Os}r�'E�|J?�y�I�OI�ɐ9�Eɜ/u�餬ݺ'ݛf��l��1v��9���d��������}pO)H����O��D�O���!��<q� ��Zr)��<�a�5�ǻ q��95�'�B0Ob6M.�	*��d�O�0�'��g��|��m�1�vͫ7O�O��R�<ڦ7�<?�f/',�b?U$x1�7A� sR��!��O�˓�?���?����?���I�y[�±l�K��uh4	�����?���?)L~��'���8OX�H�̐�U(Hc��D�k��u�RnZ������9ڴ�~�l�yd���+�4�V��$�5�?�G&�/e�l�$������4����׹U���`h�lİ�B{�[A�'���'_BY��;�O��d�O����yi�`tBŧ{�ܤ		S+:i��L-O@��s�̬%�T�ǅ܋z+�H��i�&i�veQł�<�#�ѧ"R����H~�O]����*��d�7i�\<���X�l\��GV��'���'B"���<�S��(�y�ȋoJp�AJ�h1�O��M����OR�І�D�~y�0ZB����=�q�'�L6-[ۦqqܴj�5q�4��$��j���C���u��Y�6rAN��"$�"ң��䓠�d�Ox�d�O ���O4��D�,,�!��mN�P�_�B�@T\��c�O�$�O4��8�	�O:uz�1mZAa��c��P�"	 d}��'�B�|���E�7�4��r#C?p�9�Ciǜ#�\��O-���Ҏ/d��_Xl�Onʓ��[�iܲZN�iU��C�Ґ���?!��?����?9+OD��'���F�N�F��L��~�0��W���u�����O
�d�O`�ɜi�4��.;Qx)S!�KK�Gb��� �-�#'�?�%?��;[�X�3c�7z�x�� d�	��������X��ԟ@�Is�O� ��F;<��P�&���I���?�����I˟��ɜ�M�y�	]� h�ۊ $���ۅ���?���?q�i֎�M+�O���Ӭ������_<�\R����"�p� ����&�l�'��'�'�֕ɧ���*Y�q�vn\��2�W�'!bQ��K�OD�$�O���8b#�ڌ7�6L�<6�� cay�>��i$�6mG[�)���Y&��%�daZBnm(��#n���a/Y*���'����L�Q�|�K��JI�VI�!i��Jb,�.
IR�'���'����T]��p�"U|�����8\���g��%>8m��z~�ip�Ov��'[�6MM�k�
�h���Q.
hځ�)"ήnZ��M#�F��M��O�������I|�&e�E�	��O��.�24I� �'��'���'���'���K=�a[��.G��4BCCR�$���'��'�����'��6mu�� d�������(�Uځ.�O��9�$4�I#6�6ͼ�02��t� f
�"s�*](��C$�b��:b��1�����4���D�q 2���v��T�UG-g����O����O�˓~���ǟX��ٟT#"��x�ΥQ�[,`�����U��w|�	��MK��i��Oh����M�zB��8��d�:�Qe�<���s��8�&�W~�O�Z����/��ٷhA���u��J��YZ��tR�'\B�'�"���<ic,�)F�2���9]���E���O��@`�f�d�]�
�pIx��Ǚ�3^	���O���O�o2HJTqo��<���b���������ݙk��c�Q2xUx �1��Ot˓�?���?���?��m)��l� g�z�իҁ= ��+O�e�'x��'�����'�4і�BH�޽��jƝRPTL���>��i�d6�J�)�HؖUj�B�86d�ZǊZ,Q!H�h�X�F&�Y�������ORO>�)OġBd����� Q�ޏ`�H�1U��O��d�Ov���Op�d�<��V�����FAdH @l�N�F�RVN�}����I��Mۊ⁠>����?���'��uٗ� u���7eI�>�Y1���M��O\����*����9�6���F٪�H�H�!���'���'���'-b�'�>�1b&3� Г@b�X��F�Ob�$�O<(�'�Ɇ�Mۈy%)S�q2JG�Qt .V��䓁?��?	�ŝ��M��O�Ay�&�;L�P�K��� 0!3����ˤ���')�'P�i>����,��"_��4�̛�4����a�)���������'����?���?͟||k1e��1�!X`���-o^�x�V�� �O^���O��O�	��;@�	�#�5�� �@*��L�V�m�A~��O�0����N�P$�7��@�\��^�.L^$����?���?���䧢���\r��)M�����2��2n�O��z�4lY�� �����ۅ$���8��"iP<�W��̟X�� h�mo��<���L(��a*)��'��ᩰ��g<=�ӄ=�d1���'9�	ӟ,�	��Iџ\��|�ԯG(4
�ܹ�F4G}8Ԃu��*��	My��'r�v)mZ�<QS����^سRo��x�H�B�����П��I쟰��I٦1���1�!��b�:�M�:�l��Rb ��G���$�蔧���'g  n�0p#rc�|[��8#�'�r�'	�P��#�O���O�����x�DE(u�ӵv@ޡ8�b^]�����O�@l�M;��x"�H���e����h�����C�5�"�'L��IB�B8�+�O<�IQ�?�W&w�Թ�	#"YF=�eЋ(9�H�ơ�O���O����O��}���� ��@�G&Mh���a��3��L;��']T듉?�u����䟼h��*B))��M��撮*��B�G�O"�n��M���i]�ꓴi��I$\�����O:TmRL�:r� 	�2	��_\�(p�!�K�Icy��'�R�'���'�j6g��{c.%��1�6�T7s剱��$�O��d�O��?��I�STI�c��;^��:tFƚ��DFݦ=�ݴA����O�|<��ߦ(v��ye�زsU���п=��y��W��Y��B����]�	Ayb'ůiϔx��ާ@oH���Ñ'�B�'S��'E��'��	���$�O�Q���#`P�B�I�KH��"
�O�nK�q�����M3��i�,��Vmr8�S��~���S��s(@�D�i�I�f�����O��'?��;�%��H�{"��uė�Q�	ҟL����������	F�OF�d�c�LQ�����.�X�>$���?Y�H��I���I��M��y��Ŝ{۶�a��Li8��"�쒎���?!��?!po�
�M��O��|�6б���LmKթ��7�N� .���$��'#��'$b�'}.yQ*�<�4���\4!�-!��'�[���O����Of��0Z�c�X򅈠X�i�ąTIy���>����?yL>����e+Z�\���@񉐌�@$��A�X�V ��i&.���B��x&����ĜsBй��̵��=�U��ӟ���̟t���$$?Q�')&��O�t�z4�ы]�Xq�E)�!��n���'�b'z�6���Ox�mګR�.]Z!�*i)ܡ��
]���#ݴJ)�fd  ./�&��DJ��xA��Ox��O�@�A����#}h�&ϗA�8�3�����O����O����O�9j���]eh�eA�E#v呤	���d�O`���OL��b�D�禁� M��ʵ' �JVT���P�.�d�
شJ��f�2�d�����Ġ��e�x�I-<�L�iR,G)9P�A��I�)j��	�&_r�s�'�Ԝ%��'f��'8�}��F!8ur��r���F�a�'+�'��_�,P�O�˓�?yQ��D�͚���[�H8�����'�B��?Y�4_��'��E�j�8�$�r�A�[���"���?�(ѐL��yk��l~r�O����	�Ye���$7�UIG�T4uv9e�]"�'9��'�B�S�<9���C�14�E�j�X��Uc�ş���O��
*�������q5���"�b} B�I�cʈ�!���O���O*�dׁ	��6�}���	����I#\?M���?嚹D�5"�8}q�!$�Ĳ<���?Y���?����?13(D��eQ�k�0[v�AæÍ��DU{}��'(b�'��O)��Th��ؿ@\��4���[��ś�u��$�b>5
���F�K���X����8���Q�%?9�FB?/r��_�䓯��uj�M ��I�� �C2_����O����Ot�D�O�˓?�IП��`n�+:
21�˗�탠��<��4��'w��O%��Cb�Vd��)~��x���0c��W&I&.�Х2�eӤ�&����Aj����>��;g�L}����K,P�h̋`�ru��ǟ�Iȟ���Ο$��|�O�N���l��(^�`�Ʋ0��K��?���w?��B~2�i�1O> Y��YV�ѶmX�75����#�x��m��?��(���Qϓ�?i�a��|�aUd���@�%A�"���ap,�O��H>A(O��O$�d�Oh��%A²!�ԉ�cBSS����O��D�<�FS�����X���D��N�$d R���x�fTǎ����	n}"�'@��|J?�H�A�/��٣��ݢx���D�<���=?p�	�?ub%�'t�'�`��nq4�J��Ȉ�v	1vL	�$�	��x�I۟�'?͕'�Z�1e\�q�DGnm�Y�d�|I��'K�f}��⟐1�O�$K,3sh� �>|����kȢ�`�D�O�p[��e�d�Ӻc���>����?����|4�e��3�V@�N�O���?���?���?i�������~ .(p��BNT��S*Hr���?����?�J~���r��&5Ob1S��2`���@<UK*�S�'`2�|���Ʉ�i*�F�O�AÒ	�kc�L�� �7"��h9��'��黖�OD?�L>a+O8���On�J�I{�d0񡗙kj�s�
�O<���O���<�Q���'��a��U2@�/%�� aD
�n��O^5�'��'��'2V��p(�2mUn��+�[�̡��<D��0lں��|��	�<!�a����1΄�g����aן��	ȟl���LD��0O��pd���8��Ϝ�a���j��'����?a��t\�f�D��L!*G�MU`���Q/� ��2��O$��O���>K6�/?�;*�>���O�BXy�)G+��q&��bg����|rR�����l��ܟ��IΟR��U'S1F1B�
i�|���CJyRƢ>����?������<���F�O�� B�R�{,Ʃ�����	ɟ\�	h�)�ӽ3,��c��ҏ!�z�1r!�4@h�ґ���i�)O�CC׎�~�|�[��8'��'Un����KG�O�|���M�l�Iڟ���韈�	ryb�>1�f���ƣ�=&�
�SgH��J��h�l1���dO}��'�2>O��4�I	5<`���mY7G�����bF�F����g��}���&�)z��HЎ-;f��P�ǙX�ĕ� �O��D�O����O��d�O�"|� �8袏]F�Qؔ)��h�@����'���'�r���dz�rc���B-
gЪ}!�I �K�8��6�D�O���O���t�k�"�\/�P��CN;.:0�X3�D�-Xi�� �-j:���Z��ty�O��'��@[(@&f��@J7pk�5Y�OI��r�'��6��Ĭ<�����v"�i¦LҖEx�AYVO����I�����O��$%��~���<b_ �R(�%Z�\�#�)��a����������'u��-�Y?�L>��)5��ؕ���fP��`�G��?����?����?�O~R,O���I�=G\A�*1xy�X�1�Z�����<!��i��O�X�'S�A�a��2��P���$>r�'*q��i$�	�A>�p���ΐgo���o�U9���J1O2�V���Iȟ���՟�����(�O>�y�+�|� ���[�4`ұ��T��'`b�ILۦ��r��!�2�9=ޤ�҅������	⟼'��$?�Bq!�¦M�_s��rֶ,G��jT�TD
|�	�+�`���OP�O���|�/��Dh'�^7Gw����ܛB�ڜ���?A���?-O���'�2�'�ˇ@�I�MM�@8�),z��O4��'��'3�'�P�k�5A.Z<�"S�:*P�Z��h��B-S�4n�\~�O/�T���y�jXn�⠄�y�cH�$�?���?���?1��ip��*����~�pR��'�=�%��O�)�'���'�|7�=���?�����8�B�I���t�ɟp��Ο��ɦh�N�n�T~Zwq��Tџ(E �`��N��2S(ŧ8�
l>�ĥ<���?����?!���?�ЯA����v"����;��d[}"_����q��z%b%!���.$X�sC�a���2�R��	�� '�b>��V��'�	k��t�!����NxlZu~�l�6��]���䓊�D��RN��d@ pb(��m���OH���O��$�O�J��	��jc`��jIV�(B*Y�zi�ц����޴��'����?����y�
��^+ԝ/rV�����?��2�
̦��'���)W,�E�O��NӠ�SCD �d����v+�M�"�'w��'�2�'�r�S�#�=2 ��Y\^]3@GA�,���d�O���a}b\���޴ǘ'�
�����|�"���&VU��yM>���?!�!4�9�4���T�1/��y1B0D���s��M�����BU��~�|�Z���՟ �	��0��v��<B����l�蹂�IW���Iqy��>����?������3��d8�nA&ՆUQ�iڠ	��	9����O���3��~2��V�li��Q��\B�l�Ssl����_æ�!)O���\��~Ғ|.O$S(]�7"&.�z���HW��'��'w���TQ�$I��R6��� ���I��K�T��IZy�mӾ�l�O@�$Ŝ}ض�Kڳ,��m�`	ɪjq���O<��F�r�0�Ӻ��������?娅	��=Zr݃��Z�;0�т�O<��?9���?	��?Y�������#+��ٵĊ/\*�ͪ6h@�Z�����Oғ�V������lc\�
�J�SPД��G��j���	ǟP3M<�N~BRJ��M+�'��0ӠC��`h�d\�uH5���:0����O�5SO>!)O���O����V���Pi?]��="2��O`���Oh��<��V��������	�O+̚4� �rB�,�2P ����?��P�L�	ٟ�J<�ue��U�D2�����y�cD6���:*�$����i> b�'#��Γ;X�bҰ]r�cHٴ�h!������ԟL�Ig�O��dɪ~�uZb�'R�`:"*�2s��>�*O�m�W����r)ݤQR8�膅ъsv�ڴN���?���?yw�i�mC�i��	�;8=JW�O���Fr� ��6E��?�X�S��G�k��'������ǟt�������=a��S2��+ |k��:W]ʡ�'����?Y���?M~R�w�0œ`EϒT�x���/
'b�N�2R_��Pݴ��f�4��� ��(RS��=ܤ����U*��dY1
��7D�U	�MJ���O�lHI>Y*OP8˦��?g����a�N�3N<�A��O���Ox��O,��<�PV�T��=XO&Q�t,F2I���l�A�l�͓�M{��E�>1��?�'ں����̂F��9�p�A��Ƞ�k��M+�Od�:!��6�(��权v.�ГgG� 5��{�	.X��O����O ���Ox�D.�'}6h��@��M8���o�i�z��ٟ���2���<yc�i�1O�� ,�,`��-Yb Є	��$��|b�'n��'^r�Q��iE�$�O�*�!ܿ�֨�0�E�8m���^ !�2���'.�'��i>��	蟀�ɏ<�Dp�"Bsm�
''�5Jg�!��Ο$�'��듟?i���?�Ο.h)�'�";b�pE&͗F�h�\����OH�D�O�O�1�,�S�>QH}�/E�j��G�
4q�4n�������@���'^�'%xI�F��n���;��1;�P��%�' ��'��'��OE�.�?)�_�bl����u`p�����8A�4��'EJ��?��NL�2_rS�*Op�`�aƁ��?���`V���4�yޟ�+�j�?�'f�,X��Un��j�`-=��'k�ϟ��I̟���蟐�	[�� .��f��9��s�)�~�2��>y��?�����?� �ik�$T11���`��dQ�.��B�'�'���'_B-�2i��V0Ob8`#�3vm��Č+�}����Od9�&о�~�|"X�|������7		�1�`y`FDѠ:�ѹ����������	Zym�>��?A��z���k� � ��_?��������'Q��V���y�x�$��K��ה7Ӓ�H���JNm �h�Uyr#U��ȍX����V]�O�Α�ɢVV��^�v><1����V`�@(̱[���'��'�2��<�R%<���zvF��%Y�|A��O㟰H�O2�M;�b�O'A
��c=D$ҧ�|G�l+S�'a��'�Q�8����̂�((����5rgn[�Y����tN�K���O�ʓ�?	���7��O���O��[`���MR��(QA�	`���!��<�V�X��ğ���~���<qD-�.�x	����^��y�kL�����O��,��i��&=<�S��f��c�4%dxA@o����X0����0%��'M,P�ł�	b�"����|�0h���'0��'��'rbV����O��$H�rUQ��
�?�0���@��	֦M�?�UU�`����$�?�
�C�c��ѣ#�6�&�0�ˀ���'r�Ԛ��n�O��n Hf�\���Y8�T���|`r�'9��';��'7b�'Hh<A��Âwc�xc*�~)��d�O4���c}��'���f��b��K��
�Fna0��l���8s�)���O�$�O���>�%�2hb;�����4w��Yh�ҝ&w��D	*�䓤�4�B�D�O�$�7M��e�c�}QD��(+@\��O˓r���ҟ4�	��4�O����'�m=��b7�#a9�]�-O���'��'Zɧ��S�N�y�����TrB�Ч�L��׏˅I��XZ�����"�^�	��t5�@aT�Haҙ0'_�G�j��Iן<�	Ο��IL��[ya�Oꬪ�h�r��3����}_�,s��'�2�'^�6�+�I����Oځ�H�[���ӷŇe]N�gH�O�����@|7m*?1���<���	8��N5(13���u"č���Y��S�����`��ߟ�	۟8�O�h�m�:�	�'�� ���T� ����4��W����(�ݴ�y"C�O,,�rs��܋'�S��?���䓢�t�D�۴�~2!Q�X���JR�H��CȞ��?��H�/? *����䓾�4���$f��֥�	^�pq�\��,���O���O�˓��I�����ƟdX�bZ�T��������T�@ ���i�I-�M+"�ifO*-0b��H�ᦁ$O�Rl�m�<�*��q�ZU[�%޷��~�PY{�E�eح8���";"��tmX�K>����Z2� �R�ԂW���%cE�$���C��,r]��o]�g^��I�Q��<bA��� ��`�n�z��V@ǅ$:lx� ��d7��A�)�}),���B��,���ҁC�ĵ`��W�̣#&B�q5�l�� 11���e�VJ$��`ɹt�h�����Jrd���$G�e���'.ix���5>����a��K1�0B!�$_[��b�ʎ�-~�� 	,
�H�Rt�!p��8�c��:AJ�9Y�8���.2Jb�q&�2y	�@��K�G�R�O�A	��sV�>��5C�&/�l��T��8m!�1y�*G%v}�Y�`ꏍlST��4fݵ|
��1d��,Đ�Zdȩ#J��h�#���g��Z�J��d���3um� �NQ�X:�QK�_�,������:�L%��"�c�e+��9a5q�@KZ�tRZ�
s�R�� ru
�h� M%��f��|p`��6��k��9J޴Mh��F���4[̒%��jU`��a#K�%��2�Be����f�F�n�1#$I��?I/O�D�O�$9�d�O�$�'\jk��ߪy'�`Ӏ(
�A���c51O Pa�=O��d�O ��?�i��?���iˤT�p�ٲm\5*ol�#�O���?�L>����?�Q�y���!V���CC��#�5���{�F���?����?IH~zU^?5�I+y�Jx��#�6iB-��Z����ן�&����ןغ���ӟ8�'�6p6h[�9��Hc�P:fD�-����?!���X̓�?.�l�$�O�$\�T����g�D4��i׋J���OF�D�O<Y�+�OғO�I�N�p�����m#ڬ2ᮂ$z��X�y2�'N,6��O\���O&��PE}���v��x���#WL��bΞ6�r�'�b�Ѫ<��O��'2�V��SN�6=Z���ØD�Cf鏍�?Q��?���?���?�*O����O�t�6ǐ;z٤�!��״+�8����OX�� 	*�)�U�<���R��u��������ܔ)P1kԺi��'�r�'E\듍���O���8b-�و�ĆDx��ah�1:v�Xg�� H�Dv����ǟp���[�P���<3x@�F�NI6$����<�	�����<q����w�T�iU�7qj��Z�Q���.O�t¥0O��0�;O:�D�O�D4����iB(( �D�A��BX��@��O���?�M>!���?��b�%Y��㐅ʊo�.��҉ڐ �*����q�VQ��?���?�H~JW�O�4� c�5z���Ғiɰ9�l������d�O��O��D�O������O��M�AѢl�7L�n�T6GI�>
^�I؟�	ٟ�'?��O��D�:L!X%�S�ȾhO���ćȕ~��'��'��')�����lȐ̚0DE@����LxR�'�ծ�y��' ��'�?q��?A`��z��t[�b��q ����޲���?��i�(䓏"2��e*�$ `� 8�-�w�jI�&�'��]��'���v�^�D�Ol�d�O,Ֆ�� h�Q�o��;��G�������'���͟��Z��M��kY�j��,�ի C�X�J�b?D����'���e�b���Op���O�$��(V<��
L�]�>���q����O��D�O<�O�	܀��D�O��@�+�i9~��,�w�25 �̦m�����I���I<�O��3$����%M3#.��c5F:5���'\�'��Õ���$�|Fک�`�F�Y�A��".��?����?,O��'��'����H�:=��@j"('Z9`� ��|��ۘ%ƞt��O����O�	i�TrSdT}��3tK�m�8L�$��OD��?����'�3O��M	�1~�a#��P	��c�'.j��H������O<�4�r���$��zolq�� �y;c%�	�?q���?	�"�'@�I�~�ʹ�ET(�V�[��݃^���"b.%���?����-Oʧ�yRhE�J�QR�U�I�z�1���(�?9���'F�	)B2�'r��RhJ�=ߐqz$�شb������?I��8]t�̓�?�eX?����|�;w��͸�АT>`q��t
�&�d�'���'n��y2���R!�TJQO�
6�F�@� �*�⍑k��Iϟ �	������'�����A	p���*��=/H훠�'��P�@�B�=��|�� ېD7��Q�@L4#
�ԈA	¼�r)O��d�O�d�O���<�O�<��(G#!��ؒ�I=d�v� R�����4��|2K��<�k�<a)��^�3�)�S��J���P�ieb�'wB�'�O���<q�@�F+��W�WC����ş��IM�Ο��C-g���	͟��ɄF���v'J�"DT�Rbִd��M�Iٟ�ɖ��S���|R�[�!dD+�cC1]�`��)��*&�'���Y*��D�O�����N扄nlR�L��$�����&1����<A��?�����yw�B�,�����J��%����2%�N"0���'���'�4��±х�E8:X��s��b�`;�T�������'�蔧�t�'#�Pb��S���$&� � �*03��Ԛ�y��'���'��O�'�?i2���Vκ��-�0yI�i����?i������4��� �w�(;�$��V��p�`�)L�`��ٟ����o�,�ɒ����Or�dq�##�
=/<|q�3��'�J`�-"��<���?�L~�+�P�e	V6%8 e���af��!i����?a%�iZ��'KB�'T��!���Rc
(�����_�!�$d���?��6	�'U�Ig��ʊ=(T.�b����F{R��#P/t��u�'3RLe�P���Ol�d�Oz��'/�|r�5"f�9x:�j�!F0_����:J~����'��)��ßd�d#E9[g(r�֧V����CG�M���?����?)Y��'�b;O|��G_�M�ԙb5��M����B[�0�'��Q�'�
x �O���'���Q��S��
,��h8�>N��'<2$�>1*O���<9�w�n)����p�D�� �
�A�A)O*���>O��k�+�O��D�O���<�� �.*��y����3{��[�!;�?a%\���'��[��������'���B�)|�(��7�Y����c�|9`eٟ<�Iӟ��I�?��O�b�I��"��T=|($X�FƓ1��]�$��]y��'���'�f���O劝�6e-83<����4��1�A�<I��?����?����X��S�P�H��l��������ILyb�'���'\R���'��ɧh�><+�C��<�n�9�k�����O"�$�%<C�d�O�1�OB"�'S�@\�sr~T@�CG4K=
�rw(_�ϟ������2,>?�)O8�M�j��'>�`��%�$#BB���$�O&An�ğ\�Iԟ��ɚ���C�4��lD��F@j%l_�w�F���P�	�/����4�'��S>!��<CE��(WH������Hp�V��,�	1�M[��?����?�_�p�'J((c[�;DX��E���c�'��ԫ�'��'3�Si������0AZ�S`��K�g�!E}�Suc��M����?1���?!�Q���'�r?OH�Q	��D�8�9�	8��)���'��Z�4�No��y�n>m�I����I�`�����*&���E������p�ɢ����<����y�-��Θ2�P�����aIņ�<��H牎SV&�Iҟ �I��O��i�5;ӄ�0�Ty��:��IEy��'f�	ş����T`���[����FI�z�(����0��%�j�	˟�������O)B���I����x H�ӵY0L� Q�P�	��($�T�I��Tс���*���n�d	)���
Jp�<q^����O����O��L��O�a� �$h牲 ��u�s$�!"�'h�' 2�'��Q��'D��tM6쉆w��(i��=M��$�O���U-9��D�O��O�2�'bbAV]v�� �O��I���X��+��'���'b)ڎ�ԟ�1%GM������2	F��c�'�*I��'�r�p�X���O���O�'�^I�7��4v[���R�����?i��HQF������IN(m����G^�rhW�+|�2��O��������������T8H<!�{�t �3�<_b�9b�-�~'j�Q�T�d������i�����Oh(x�m��P����`�*p�QdC¦���ן��I㟌S�}��'��� V"�J�
R(���CCh���r�'��'p�-;�'P�Tۚ'�r�'��I��>�(�����4X�i��ݠ���'JJ9��OV�$6���r��ر���5"��ЌL�U�˓8���L��|̓�?I��?1˟�0��䄕��� E(ѺJ6�0�'�HO��D�OF˓�?q���?�w�Sj\9�+D�<����,Z8A��~G����?���?H~�$�OWX=xW�	�NMi���9*��`+O���OJ�O��m�`j���O���G�˒')�q��˗UJ."��3+�D�O����O���hq�OZ��_&s��ȃê_�F=�M�B���?�'��'>�'��'�I���%�$�M=/6�훔茋Wb��d�OF�D6v���O:(�O32�'�RNV�A\�`ӂǑ�E��G4GV�'�'0����'z�'W�	�+[��P����-��ϢPR�Ѱ�y"�'��6M�OH���O��� _yb��?���!�42���w�?�?���	�5�&�IU�IY��*�8V���G�����Ccڈ?.�%���'���o�V���Op�d�O���>����W�l�g� "D�Uj���?q���?iL>q-��c�6O���a�d	a댌6�*q�@OE�Q��m�⟘�	埨��-���|Z�O*�!�4U)�|;T�h{�L��?Y/O˓�?i!�E�<����?���i��$�7�#g���Q(ӈ4<�����?q��m������ɧe�h9��۽u���-M6 F�O��$��_���O��$�O��It>-a���R�����$q5��Oʓ�?a��?�H>i���y���Q�t\6ϋ7Tz�����?Უ�B���?����?N~B��O�d��$%�#�Pa��!�L}���?Y��?Y����'��5:O(�{e� ��F�Y�
Ii|�cge��y��'�B�'��t[>��	ğ��	-c^6�IsIA� ��S���i�I���%�l�	@y"I�������S�	6
~�ʂ��k�����O(�$HSGz���O��'�?���?	�Ě����qѢP�3
Zp�ե���?Q(OġY��I}��y���0���8�-��N;r��	C�I,��4�?���?I��!��I�d3��#b%G�J/��K��9�V�%�X�c S�����@6�27�G�*�6�y�g޳E����r��7�?����?����?���?	.O�ʧ.[�Y�J2.��I�5�_� ��I.OFM ��i>!�5@�<��K���B��.�$�E�I ��l)D!	�18�J�2X��,�mNI��Cb/+���1a�O�B���=�2	�Yp�M`!v��xmڵ�?A��?��'��'�?	�w��Xia@S�q����QP�]�8�	O� �x�,]��$�y*�6P��4�����a�U� Δ�I�J���J�߈܁Q�Uh�Y�&��o�ض
� &	�% �N�zZ�aمc�X|�ҁXDM�Ęq#��{ 7�
:=�Xh���z���EH��^�������t��A�oE�b�(Iu*�+(m����R�.�GM��B��"����`�*D�槝�dƤ��N
j��e3d/LXI� �N4]�� �^3Uښ$!d���L���K vѸ���,KL�<q��M-��+F�c2d��Ҏ܉/E�4ز�:@�*�K�����������IayR�ir@J��%��7��;Eҩ��F��x�n%���t��/������}�#��[���аJޑ ��È�:q(\چ@՟\pcgģ��1rH|�>9��o�",҂kߘCq�%���ƽC��	?0���$�O��=��q�j��#.Ԟ-��zd�ܘ~$�C�I8:��L��ցu6�r�/P n�	��HO��My"�P;~K4EC�� m��[��E!_�eZ�ds�4���O���<����?9�O����o�7Ih��m�x��e�Ȍ�(�j����:�0>��J�������N`���S�S(kS<��D��ͅ��> ��7�<Y���g[�xh2��@�aW�z��]޶�?�,Ol�+��*�1sf�	fyLM�t�+2� �"O�i�ChV�v2��QI���A�>�TG��\�'V�5{��~���M3�ϋ%r�X�Ț,	�)����2#��I�d��֟�s����݃��Bf��X�Ӻ�ІV�^����M�d}`�&�m�'�<�1�ڰ1��	pnN��i�2g=@��wg�:u�%�1n��jv��$���O��d'��H;t~��Y���"k�@�G-M�oc�İ>��m��Ƀ�G�{TAk�SW����'5����'I��y��ж�>�ZR�<�wI��aZ���'�"��$�'қ�,�=_n�x��KА���̞���DQ�Pȱ)�p��D����t�3$�s��N�/��ka�,��D� ���T�D ��;k�>1��d�'*<-;���X�Rd#bI�>��i�����	��M���H����S���xP�0#� ƭV#�И>���װ=ACG�L�t�j�i��7F�E��4uў(�ܴ�?��tj-^�� * �M=JA<q���)3����Ox�dҙ+�l�� ��ß��D�Y�  `�gaξYJd,���R��BM�Rh��!,O�a ���;�z4rA�8l���e���v��um�4X2���'������%�x@ K�+��h���B��	�	`��������O�7-]0I5���F�3%^�Y�"S>?
�~�_��Q `�*��rn§K�~ᘕ½��Bٴ\�V�|�T>͗'̼8� 64!G
�5�� �J�L������C��M��?9�����O:��`>����'���a��\:��T�Q	UȐ����r�@��$(v�BqB��)r��Ȃ�@�j�a�&�MC')��\�R��P���sCֈk!�*t��|�'���a����K����	u�P� �@m�ȓ"�: Am�$0�q/(�4Q�O��'��I��9`�4�?I���M��̲Cd2�+�Y�Q�T�ŝJ��I�Aj����<��	���ŃTO���pv�ԇ!�XE~�H6�H�9;`�֙P$J�A��Z�<�mc��	 Q����-��xT���"n��ѺF�ө;3C�I"��'�O.K��ls�Q������\?ٕ�׮p=шP	M�@k����D�<�Tn��/�l�WE�3�$H�ˍD�<Qt	�U'��s���x����F\���f�H��?�0=�P
�X}�O`5I0��CX~��ML�_̚I�"O1tL�c�2܁,@�j����f"O�A�a-S9^8Ԙ���	e*�]I�"O.�k�HŶiv�X�ǋ��F+V"O6,)2L��	x�I'�>���"O�yP -	�V5�pb��CRry��"O�]aDkɟ&  pqkДwA$�
�"O��#rmDC����W�19���"O� �LC��"�k֭�3>:�E��"O<�Ê�C�i˛�'dm�"O� g��Vz��F�U2��2f"O�}�	�W��aw�S2Eȴi%"O����):��HaC	�)�TZ�"O�0��L\�A�6S5(��W���V"OT=�
�tհ	9CfE�:tQ��"O����--"5 ��Xm�9*'"O�U��F:lM�1c�\6^��	�"O8�w�7@xd����]�Q)�L�"OZ��#�Ȝ.:\���S D��j�"O�M�æH�B��Z�.=��"OF�`d�F�{�\q��%��u�U"O��s�P)���FIӀV�~�H6"O�Ȁ���.+AR�AFi?}�x�d"O��#���1Lf�)�U.
l�U"O�$�䤒�u��r�ŝ
�=��"O�qQa��$p��]��/(����G"O�zǋY�
D��m��I&0"O(!чĭmaX�0lC�(��"Ol�&�Ac��`��W��Cg"O�xp�Qt✑�lY1t��"Ozh�!(_�ᾕzC���Е���T�<�en��usF`#"�m g^�<�"����8�����ūj[�<��'۝<��iX�%���ň�o�<��&�[=z��3���LP<#�EIo�<�j]�)�0"�KZ�"�J�f�<i��:1h�%�&M� � q�cL`�<A4b�
H�^X��X�J���D�\�<��$�`��Q����!n`�  ̗^�<�T1Q	vУ�j��Qr��w�Ll�<�B�H�y�Ђׁ�I�B{be�o�<�7�V6A�$@��v!�����g�<�U�[(W�4$�j��nw��J"AY�<AJ�0BRA��^;�P�B�L�<�b�Ύsd�TpU�<I�d��u_g�<�4Z&�hH�"ՖJfޅ�H^�<9���7	%n� �mS�L%H�+�r�<Q`.�+���C���Fa�TȀl�<9o��*�!�*�XH�ٰ��o�<��`�%��Xf �mr�$�k�P�<� ��C"�T�n�$�x��y�>D�P"O��ғL70�D����|]� 8�"O��ŏ�P���8�GBO6�3�"O���D!�v����w#I#C�f$�C"O
L�P�[�/��b�`ʁw<�P"O2%K���gw���RO�P}e"O��`a�43�r���i��c`Q:"O�y)Q�*K���	��ߕ����%"O�i˕"�m1t�"�ρ=��;�"O�4#�iW�0��&�[�`%3t"O����
�V�DL	��S�@�"O���`�ݨN<UC��G)oPډQ�"O����I�BjP���!�"4"OZ Q� ����QcH�U1,=��"Oc��F3l|�(�H�4&.�A�"O2�"�
�#d�-
F"���"O���D]�
�ԑr�ES��tĻ�"O<M�h��VBtY��D, uh�H�"O���(Yb�h]�)W Ίb�"OBh U���	��hT,�d��D"Od	��.\�a"����br:킗"O��'#��A>�!���Se�	�`"O�!p��Α_�&��B� _N����HX�ń� AqO>��R�'f920IA ë2&T�X��:D��z���)n�:��D�A�pvR yf�'����rsXYF�'O\̰s��W��z�۵~utm낑x�b��j����=�O��}Ѱ�FW�X���
5Gn(�# o֢m��t( E΄ܪXc��{8�0H���0��9����8�m೧���8�y����F��@sK~o䩢C�ن>|��]�_l8قB���\�������1.SB�	�^i4)��G��G��bG� �@y�r/C�|�[4o@)sH�@P��Ԗ+�<(��ǎ�F���Б��+L�^0j���y.����~�h���Щ �~�S��>�'["��t:�Zb��	�%�y:�}p�O�!4���束Q���Oz2�?I���u� �����#r��@�!n L~�K٨B��mѲ�\@�T?U������:��C�\����2�è=)�8���.�*�O��.O.���'��Ͱ%B�]�ZR�0�S$�H�b�'��1�Gɋ�����A�G��E��.��$u���Q�w�h��%O)s���%�4V���	�=��p�>, N_�e`=3'bL�&3h�
� ���}� �V�q'Ȭ	��/18��4�Frg�0j��N��T��
+F1F�>)WfN"4��;�Ʉ;��d���t@�N�h$��[*�(yfHY��%��e-`R'&�,G��'@L⟔�U�]�$M��9���x'
��G�e�PZ��� HtD�bP/~U��av
8���C��MY!��w�l��s�\�3���P�"�E��s4R���JNJ��ߓ>�D[�B�+�r@ؑ(3o�R���s�tt�q(]1l�Xu���5+�t���G������UǼ���?Gg���ա�h{8�`a+V����e�k����@b�X�J����S���2�|fρ$�0�;gl�;��WPr�'�Q�q�O,&���Z�ȭ���}nZ���ą�C�f���k]���D]�q��G�Y����qbíFp���F�\�$�r��y����䋑:_��M���'H�M���L^��.�e�>�dN��|�h���X`��Wv�rt
bHHl)&ݒ�"O�\�Q�M�;��5�S�b�2���_��Aum@9��$c��oyZw�����d�$8�M�O�G��ec��
�e�����C2Pq�<��m�(��T�]�fд����@���:(O�U붮ΐ+d\p��dW�i9���&��H#zM��T�;Q�Љփ��<hm�'u��m��������9;��%�^�k����h��8�mٶh�m��a��q��`'��>9�,,q�'Вy��Zɧu� vi��K�1B�@չ7N� [l��ȓ]�Zmp�' ���Y���_�d���'�h26[.~�ɧ(�~��f�̪*�����-�2ar�"OF��m���y=X!���ăx?\)�
Ǔjs�Y���*f�G��L%��>=���v%E�F�y+�`ҋ`�`}��'l��GB7�8Ap��m��G�F�␮ �Y��*A�ȓq�����%,r!�)e��oڣWݚT��� n�)��!�+i�\�3j�4�
�0"fԩ�y
� ֩*2[�+��<�E�����rS�O�UdD��*�4L`ӓH�N�s�&��-J����Io}dM:4.�%b���x�L�<Q2�P�E�j
� h�GHh<ń��s�0 �w.�e�VtH�n	S�'��5!�ʈ#�y`��I�'w����mJ9��+��˪3O!�)q |�Ћ6(�ᢴ)U(<�,�*�@ƣ��I�r��<E��'�� a���"tRD�ל>/��s�'c�����Z -9p�K�ހ2JH�9�'X��R�V<3q� ��'<^ݡ'�1wh��׏+��iS�O��Ks(�����I.]vA�f F)8�R	�&��2W�x�x1��pH���fo54�dc"D�N`D��CY�
�b@	��1?���G2bɀr*��i�T�P	��Dʨ��db�f�r��B�QY�4�@'/��>a����_PDܰ��'|�ʍ��H�W4MR�A,�<t��o�{��I�Pe�<��I�?���yR%K'r��`�qJ&��PC`��(O��rf��p��t�!�������� �@���w��3�8��V�OPP@h�?�@�	ׁ��S�p�=�OSR����ܺ*�$��"��w(*�1ՋH�ĵ���J(X�Z���Oq�n�Sq�݈(�ZTrF(�6�8�* � L���M f�h�CCʓj�	@��~�/٨�\p���[�f!�����������ŧ:{��*�B��oX|9�ψO�9Qc�
?8쬨s�)�!���٤�ik�A�wg]v�<�E{"��en�L�C�H�f�$$��P�6w�*dk�$
�Գ���3(�mG2(�!e� �3O����f�Z���"�&����a)�	�<?�8�aeL�E�Ly{���!#O�A�O��uj�Z8xjhВSE��T��S�}ծfˌ�æ	]J�O	���(�;��]��D�J�������-�@����-G����J��h�j�	H�	Q3j�$f�<&)B)Mv�L��0��E�O��E��O�E�����@��	�y��}���Y^��hp�!�4&���/\�)i���	
o$(<���#ba*�Hݢ��6�DD��cפL#�HOe
��ݠ�Ș���Ô�^1g���.JԈ��ꛀ2a�`��q��"?A��=R��9#E�O�C�@<ONp���9M�&M���D�K��Ac6�Ղ���"�˖.q�T�'�\	 �
ȼ8ބDږ��,i0�>q���~�Z�<�'a;�j��:�@�b��6?~y
�c۠"�
�s�U/S	:C���g�O��B��,P�&�� -�$(Y�� �,�#�l$h��'��>���R��T���&"0 �����/w̪�2Un��"ub�C�y$8�2�l���">�!��:�v�`���CC� K�<�c)G'�أ>!��S��U���G:G&pqP/�Uw&�{1��Y�Vt� ���2!@UG"��B�6�?7͛�(Z�<k���
aH�Q�4n-���-�6ZV��9V��3ʜ ��~
���{NP�ũ�!����e��]?�S������r�az�KDd�aı�I[��ơEO*���VLH ��Κ�w{h����.ڵvd b�DB	Jլ�2 ��Z�zY��_��JP�CO�����L��pX ᐓ3��P�ԧ�ϟд�-C�5Hv�ѐ���N���>�,�ͻp�
���"J�;�\P���K'PL��ɟ�H��R�^�x���х��0vD�( ��A�@�qj؜X�\`�E ��I)ctve�������a�&J��Lp���r<�iD|���w~:��d��W�',�>�K�Iľ9�}P�㖓l� ̓u�J���@6`-�ϓ\�v�9f&�6e���J�x��a�'�-� �G�S���ו#�$ѣVK�0<���F'���R5H���;&���K�O��z0,Z>)~.���?M4*�Kw��}�p�U ٶxT�T��Iϸz�V�����-x�f���}�<���]&>���F�D\��WE��[��}ڣA��Mj�0I,O?�	5�֬��_ƀa2ghΚ(�fC�	/I\( ˕�	�s�r�H�!L13�d�	�H
���kF`az�4{�A�D��\����՜ذ>R�_�8��tj��xx�Z"#Y�]F�yJp�L�_!�W�� @�f�@( l&��:�!��*R,��W.j�6�a%�#�C�5r�z��`��>4,���OY+��C�	�1`��cgaXWr��9�C=E�C�I�	�i��I3`H�2&%:o�C�IB�]#g��1��Y�qLܽv�C䉁n�rt��'ѳV��1��H���C�I�X���1��
�ry��&�,`C䉭A�\9Յ�:s �(��Q97V^C�ɾ%���8 ��+x�	���K�q��C�I�3|b�����n��o���C�ɦ9\�C�3���umܦzC�)� h�B���Y�(A��G�h`�٘P"O�P;TlF3j�2L9� 	uS�HA�"Oй��F%*ba��O�x\B��"O�	��S6@*�Ag�-w�|��"O,���X�v%�"
9*<���s"OF��c_�q��bŁ]�pJ<D"O�}��b�F�9!�߈Q0hڤ"O{@��.<����*4(�)ʢ"O΁I����Q�$|����W��t�s"O|��qME+Z�Y�0'��Q�u"O�h#A�Za͢��!K0<�Haj�"OZ}��"�1�Yxd&� ;a�p��"O��b!�R�?����@'S�|h9""Oqj�BQ�`�$�m˹3��|�"O�ppT��77�VT�6l W�$y��"O~  �9}Ǩ�;�eͺx����d"O���,U_�8A��f���D*f"O<�G�]�	�"��:V�4	R�>i`�r�2UjT�� ��T�G�Ya��F%��Y�O�+8S�)�P♞iQ�]�ȓ	Ҧ�Q$jX"���/��ܝ���� u���_�Jq`���2-�F���b.@�!*��0¸�2��4�e�<��P�0y�E0b�Źv�rܙFǃC�<� M&c�����R���L~�<��I�T���C
ݦzX�$�b�Ax�<�g��'�f1���y�U���t�<q�ER-0\v���A�Y�<�c0�g�<��
�f���	+�+O%x��cn_H�<YE�c���h��o\4M��^�<���6F^���'�۶T�%��u�<	�G�3LP�����M�Qn��Y�kr�<�"=�� ���ur�)3��m�<q#�
h���Ф�< �� ��/t�<��d�'r�>h�T'8B���؂i@n�<)&�P�z<�c�I۞k��9t	`�<yT�߰�LR oǯ�d ��w�<��Ш'F����M�jlR�k�"Ir�<�όEB�;���~� �Zn�<�c�D�(oΩ(�eځiٔ,r�� n�<�H9}ځZ"�WD:X�s$�q�<�CS�>���!!,]���
Zs�<�	ґG�VXY��Ѳ{�^�a��Ap�<q��+Izݢ� ./��@9���h�<I��9%�TQ	tC�#&�,=�6��f�<95(>�	��5J��q1�ń`�<I�mΦbl�i�2�@�W[P��҂�\�<Q�ˎr�vq�c��ᄸBED�<�&�
,}Ό�%Bg���p�j�<a�� �\���U�$_IK%$	q�<1��PڰP�������Th�R�<Is,x��X��O ��kg��v�<����qג��&�A|1�-z�L�<!��ֵi"$a��d��94Ǘl�<y��H�N����Ь ���i����k�<��'T/VD�Ւ���@4�Dk��e�<��H�H��A�F��(-�^�<�L_CNX ӗ�X�F�n���	�c�<� #+:VT��[�_����g�c�<y0V�,<|��!��l|�hD �E�<b ^�4y$����G2t�tTP�#h�<�poոx��Ȫ�BK�ih
�At�M�<1b
2��%��M7()Q��n_G�<Y��J�Q��H�p�ZY�V@�L�<a$ҲA\�����pS�!�;�y
� �C�(A,��%��%~��q#"O�)�/7k9�P�F͎��fH#"O�	@U����W�Uτ-hc"O\Ͱ�!{@ D�S*>��=��'��Q��dTx�;AmX�" �I�'�1Rp
�Z�L*�'Z\��''�ă�t���0�Ď4��� �'����(K=1s�h���6(�K�'�U���Y,>'v<�ݹ��h��O^�8�Yy�S�O^�9ie�"A����2)%f-��'���e�W5_����'N2�@�yb'O0�`��I�c��]�����L=�5�d�O��C�I�g���땉��Ʃ��f�ޠ��-ٿZ���DTo$����f��@�C��g
ax���X�=y*\�o(A��2v��q���D�<�v���)HF�k�bH-tv8���Al�DĒ^���>�2��P�x��}��!S��J%ط&R_�<)���~�4<C`�*�$�+W&SQ�<!��!I��\��g] &��eK�P�<iD�S�I���BDF����R�f�b�<QQ�1H���HpD�k��"*b�<��͵of�H�T�^��y!,�X�<�3�ΖnL�A�zذ`°.�^�<�q Z�{&YȤ���&T���Z�<���+R���8���Vs,�i�#�Y�<�A��M*��ЅȋG{�`YG��S�'���"�S�C��|(�I�2tvh��A
�i5�B��?UB�ʀ�ǫy:$+aS(!��S�(D�L(�O1�a����>Y�)L֎�3ц��nj���t�<y�c���U�'J�~~( �� l��$�:����'���8�T>񻔠Q�I�$B3��1d�r�A��+<O$@7��$7r�C����`	0i����x�a�,uI6):5.��mS��٫gf�P�l��c�`4Q>q�=	$�U&��U��a\0��2 QU��ZC�a��m�j�@b��Ԁq0���$��n#�5���t�<�3b���2jJ�Z��`B�c�xcaz���4��!:����2�˖N55�8Jwg�C��|��'��UQ��$R�h��'?�T���ޓ�^mxq��D���*R�J��S�v�xhkS.�5,�
�*o
�4>��?�OZڕ�`[�-Jř�Ol�P9��1,��bg�ԑ�܀��F������:�q��o�΁�2 B����3�h\�;��#�	;(�\�9���j� u���Y�q��b���g�֛2� ���ǅ*Ik8�t�2}��+�=r��H7pL�xWn���'�Zp�֢�4�@��%ϳJ� ��¥�(�ZH��)8��=���ȫTH�'����3�ΠK
�t��I��
t�zf ����=y��2����oې���`��P(<ICɛ&��j��F�\�
�䆬������.~�yvKF�V�5dM�&"�P�٥�K-u��M��JR V�xrn�"o5��3i�	� YS���_��xQHLfw���B�Fo���=!u���	���a̛ ��1��/�t�	�E�f]K�޾R�`�t�ݜ5Ű�'%:��@��y�`��@ƌ+)��ً��ڭ
~�ؤO���dxҬ�)<ʬܨ䯙�z����h[��0=�E�ţl�Y؂ ��]jUc�B�6\=�Ů��m����	ۓG�bū����qK��C�"=h��
�'1�T�7�5;�:HqG�&VՒ�%
mX�t��Hz�L��!�[4p��2�k��	��iǶqHV�Zvb\�p<	"�Ɔ][� [�bɩ1���Å"��s̗!��hЄ����'�HtӤ-�Q`�Н1���P����bc֩_��|�`"�0"K:X�O \�&�T!Ėu����`kƉ��'Xʵ'��-f:��U���j� �L1���f�H8�D(0#�= �\X��N9\SL<��HU�B�����ݥ�악�	�yWe6�D�i���A<������Px2�#�ne�֩_W�>�6@��C���E|r�ō,W:���"�'9@�q� 6�ybk�ux0�T�ߪ�5"�d�n�������^3�C�ᆍ�jU�0����(���X{�qAa�OhYX5�ѭp�X�1o;W��U�4�I�_���X�o��0��q���'_<,c�K&6cX���ҼQc��J>�r��>*КC��q�B^(���9�J#�H<��ɤ9Gf`�R�
m
�ɠDL�rM�wl&l�l�Ң�x�	$h�|��	�L���*C�aޥ#��yFH��>w�N̐i"4�|� Ёb�G�=���zN߭}��p �&�$��ۭ���	'0����>	W~�����剡5Z�p)�g0��D�u�ځ#S4��dMg�E�q�ʡc�4X��Nb 4�$��n�}�`��6J+�q� ��t����&?�PXǓ_�v�0$S�,@Ly�r�-��&�x�v�&mA��f�K�2��̄w��O$ͣ���y���bCg �	`�̲PI"4�d0�D1|
�a�ٶz����^&3qH���P>V\�l��Ϲ��?���n��SF�ҧh�$h��	x��rE.0D�dj���47j�,XB!
e����>QLH� AjU �w|24�tm�{�'L��@�@�^\D(��m�h�P�n��I�2�V!tU)`fE�r�:���'��sp,�AF(BP�)s��X�4�B�����H�*rʠ ���_����S�+�	�j��W��.��5�&�*�ҧ2�,.j%�%��9Y�^��U~K-w��:ӓw��1_5k�[3≠�m�
<�`��N�:oA֍z&�1}J|:����s
���f	!u���bl�"9�fѱ�M�A�<C�F<VV;p���C~�;�mX9��C�RsJː2j���{�8t�?}"���h�PD���� T�(���ۓ[ J����W}L�$�ʣYNtQ�D�����5#[%r�=��H	���ZD'���*HQ�5�/�I(TV�B�''��(U؁(�c��>qF'�E����H���'��u�,!��J1
��1[�@3?���f.!��ɒn��lu)��wH����Q�l�?o!�!��⛶�K�r�D\�ʟ�x�kH�xm��sAB}�Z!')�.
q���A"O���޶z��P�%���m*��!f���l�S��h��P�ʻz��	�Ǯ~�yr�T� �TD�7�K�����$�$��<�3��A*��L�d�$�9g�[0>J�@ �)<əO�?8��t�(4�~��뀼iq���$}��!��Os0�MS6+b�'�1�ECk�����-.�0�2K��?�O�KS-X5Q���Ҭ�3Dp�
�'��� �܋@ (�ʁցY�*X;��/2L��
��|�������M�|:4#B%+G�[e�H�S�������ƝE?!�DI�OZlU� T<y��02�*C�s<L���^妁�#E<&F�d�p���	�٨�I<ғ�j�
�dE>9��	0G�7V���ɪ<�"(6h��W�})��@:vv�2�⊊����� �&r�Cbk�鮩�tC�/��{��E�JNк'�M���!Cԉ�ēZ����'J��S���kO�9:7ĸ�g�¬]��đ�29���A�İ��#ǂ�$}��XQ [��!�D@2\�`Ai��-h���
#M%�#�v�X����@*,0�Ib`@+���)����n�
�X��88s�u�ģ1D� �F>U&P�Y���D��D��D��Rg��e@HmV�,4<�	5��6M
I���'����R�!$���%ǒ[8��k	�I��-���ԏv/@���g.�t\��&�ID�uN��v���A�%�Ry�@,H�U��Q	�2^�	3���]� X���(?����=��n��?=đ���U�1���9��"�?��G)Y/�(�P�y��7��	a�p�����M����74lT�Ae
+���9��ќ|@�J,4�&a���ԭS� ��t�Tc>�5� � `IC� i����ҕ�"O���`�!OV��S��ZT��2�X	O�p�`��ul,�B��-A���F~��/�4x��H��+�r�!Ve����=Qp�K.*��P/1<�5�m�
:t���$K'4���R��I�0����<un�h�④-�ta@蛓F>�O|q�����#~��H�v��d�dHЊ}2��[O}�'�$KJ����2LO,e�Gl�Ek��̫<�"���B�-peC�{��GSFx�4-с5 |A�� �|"�������V�(<�Ɠm��mI���[��Лn��Fz�D�4h�%�6$�K���vp�p�ò?��ҳ��
�$����"��$'A�/f����*�nZt���u� F�S��M;�$ҵef��
�a՛=��àhj�<aO�@��i�`l�?s⽺ҋ�cy"m��YF���w�+<O���g�p�"ِ�B��ʕ��"OB��`3#6(:�Ă	�~	��"O�E��(9��*�$E
���1s"Oj�P��-�f�����q�1�2"Ov�"P"�R���Q��O�M��xH�"O�ms��B
���!�K��e��"O�D�FW��6��3��0W�h��"O�%�vK�^�� �M��SμAr$"O��B%������	0v��U�i�<����GlŃz�b�#�`�<� �<�#�M�~ڢ)�E��c����"O�p�P�R9e�Q[�%Q4,�x���"O�Q�K� @�01���H<�w"ON(��*P�A�ś�n`�"O$@RsKS�n�=9�N�^�(��A"O���g
M�w�ޑ[�m�4g�*��&"O51ThJ�RG���������"O�a��^�VN\��P�p{7�Z�"Op�s���%N^@���M(���"O4���F�.��I��G\(U;V"Oi�`�߆@s2[Ġ��V�h�"O�D�҉S.ph����ء"O��S��,�"H(��F2�0śc"O��3A�g��m�� 1b�<M@�"O�x��c��xf����&G�P��$b�"O�r&�l ��5�Ѐ\m�9��"O��	���3��z0�N0ub���"O�!ҥD�R�x��A� �h5�"Or���$��
My޴H�"O�y�c��7W"DPnX�|nH`�g"O���.Y T�(sR�
 h�<h�"O����ʻy��;� Qn�V��"O��`�o��rX�� G:<�: "O~D�wJE�Nº8�2���-� <a�"O @�LƞATj�cF�Q�/�R"Oz��1�V�_�� �/%���2U"O�� ��)T�(���Z�<���"O �	�-��&����cLƲxS�0c�"O`��k��y�:��B�A1.D�U(�"O�@�3�Q�D�0'-b1"O �¶�44���[pT2m@m*�"O��I�'�<3�lu4�i�8u�"O����BL�"nm"�@@���"O�Ip`�Q�Od�M���K�:����"Oh���	.�|}�al�w��j�"O�=�@C��(��dW�Y�"��%"Ol%	"dN,O�\`C �Si�C�"O�L�gJAm(՛�<,�1��"O�1��'��8����@�,(��z"ODM\�WxZ����ΤP�����"O�ax�J��vq7�ӡBy� �q"O(1��"�29����Ѧ^rP�1"O`9�ʝ�<X|�E��Q�4%�"OB�UhӉj�*�;�	 � �pK�"O�y���+J��� �� ����"O��ȣ���|M+'Ƒl�tȲW"O��@�
W�5��JĞ(�:�v"O��)G��L�̅xE�1e�xYq�"O����#@������u�1D������X�h!p��P�#!��m�C�	T?��t� <�V�j���:7�C��4~2lk���2T(�	�!rZB��
1�I���<}��S�RPB�ɪR�Xj��ia���i4nt�B�W�⥫�bȲ#%6\J�엂f��B�	_X��S6h-[�UK���JB��-áS,Y�[?�!��J��D�C�	�?%,yt�T��YT-T@�tC�I%��.��`�5��K�N�zC�	ER丘��Kl(ة��b��jC��t��/M��Q��M)",J�"O����A)^��8��K!88	sf"O����MֳG���U��Q2�"O�c�LQ+��sС�1 �&��B"O� jEBĒ�v%�F��S;�Ȣ"O0�s��0����1dE%e:��DY�<Q!`	 �A�AFre�P��M%T���q�����7K�&6��1RSH"D�x���J�z���ƞ�I_|�:1!D�t���$�D!t��)�"8$�=D���!�� ��tSR�A|Z����%D���,
�Y�XCF���p�r\1�8D���CI	yH+�L��~�ʧ�8D�L��G�?5fl9��Ŏ8Qj��FB;D�dp��N��h� ���4�F���:D��XP�^�{����&�**�>�i��.D�(R��?/v� S.@�N� )��%-D����Ob3����@���۱�=D�,���?��m$�6_���Xҫ.D������,/��4��F�-�"�,D�@��HJ�Qh�K�]G����O?D����L�D�)�G?L�@:�7D����G�31*%K ��@�����%9D�<�T�y����Ô݌���4D�� �I	,N�E:��@�}٦���3D�D��&L�e@��*R�B�qHq�-D������?�>�sR�P��b�3D,?D���q��'.�]R�@��@(�L9D�HW��b����6
4$��;G�6D���j��T�ԍ�g�U&Q3�U{�h"D�P�%�%i�څhR�b8<0��>D���t"��~\��;�'ԼR.���.D���#N-G|j@S�������,D���W#��5�=;�d��u�"���N D���
-u��Ǎ�
K B-c�	:D��z�΁E4X�
Q8lU��6D�p�6-lթ���#h�\e��>D��a��.�n�8��Z��b��q*0D�|�V���x�,Z�xuc�-D����I<%��{˖*,��� D��cw.���Ӡ+��A�< ��f*D���')"!0���B��B���.(D�H:�O�-r�����&8R���g:D��Z�i�|$��fI��Jmq�b8D�l�2�	$�ԭ�%��Zy�3h4D�İ��B�JZ؝q0j��L$��j�!>D���pK�?{�&9!����7�.D��� ��`�� G���$��qs+!D�0���Ӻy�<��e ��n��	-D�L��-�,��=
�Ǘ�n5b��� D��@&��"��T�KԿ0<!���?D�D�ϕ�Y��cVx!��=D� �2I\�z�U{H��<���<D��8i�����i�f<hlZQI:D�\#���=1�X˶��)�Z�t!7D��YЈˠk�L�i%�$#p#gh?D�X��@�!W��1�ǆz�H��/)D�cNV�1���h	} =�J;D���W�L�,jJȢ��"�Ơc#.D�z�f�&yH��)@�/dO��P��*D�|S�i@'( ��D*hLf���4D���w,�^:����aX��^�Ҷe1T�����B�?-h8`��D |�4I�b"O��r�7��HV���s�lEJW"Oz�[gdڒ2� �fF>��H�"O`��Gf>A�����`�*�"Ordc �@�W"Q*��ˉ.!�Ȉ�"O�#�D�W:��v��4`-���"O� ,4q k_*� `{��E ` ,{5"O��1��Lmj9Bf��1rۮP�"O`5	%��T� �k�Q̈<2"O�[�+�w��P��ɘɖ�"�"O�\PրVs��\9��P�C�0�"O��Ӥ!W�1�>���X�W����"O�b(Ψ~>��Cb�m�E�C"OdQ�Иu͂�1 F�,2��+u"OL�we2U
�٤�	^���k�"OL�sg��,��<9�Ì�0�dI��"O�܃s�U%2JȜ��a��&��H!"OB��p�X	OGZ����G$wd���"OF���C|��Q`$Kͧ|ul���"O(����ňr��`��*��Pc��R"OH����\��i�_7qJ�$ �"O��B#��"&�b���P7j-�R"O&����F���
��J%K5��5"O���H�GeX��_�@B� �"On�{��܅E��i�f	�i&b��"O�)�ˌ/!�`�q�ג#�}xB"O�8 �_w*
�� �_�	�x��"O�q��i�I�t�S�e'L�p�z@"O֑�`�U�2�|��c�y�N��@"O������h��ܰc�&��ȓ�"O�%�B�-�@ �L
N���"O��¥G��@����z@��f'!��N~
Z��v���I_NU��|F!�$\/@�D��;RVl�� 	�z&!�+c0*�`�%�%8Pjp)��4!�D��	 ���K���4a�o�%c�!���.:)21��͙4�t`F텾e�!�$D�-W|E�J	�tlp�*L��Gx!�D�����Tʁ�;�-�D^#*;!�֒@B���I"� ��5N��DiӌpT�ۍM��=�s��4t��"O�u(@�_�6�� N�
e��D"O��֊�{W�la�'@B����T"O���� �^�
�1�F�ߚ��"O�A��j�3&Vb������6��W"O�A��ΫQ�֩��gIl�X �"Ot���M�&9��}��a��u�!!"O��!%�æ(v��A�&AX�@"O"�v�R����{��^�Bdɣf"OΩQ������+Њ��D�\�!"O���&ŏ*B%B�)P46 >�S�"O��.�\�.U�iG�I
��"OZ�R�aִl�}���(P,��b"O0�r%Ȁ$ndR�As��D$6��"O21����Zy��D�L}�}��"O؝�$M+?ܞ���$^4Z6#�"O
<����7j��!TDZ��"O��[��M�
���i�a��)J�"O�����=?z��s�Hդh�� sf"O��s��}f� �N��F�&��"O����15\j�T�A��(��"OB��OX��������7n	*v"Oz��i��Lݺ<X`��0H���:G"O2|z��W�n�����	�"OR��r�Ϻd�Ĕ��!�
^�t��"O����eE�k��uK���0t�"O�ZwkJ`L�1B�8	�R=H6"Od���%� .�`H �f9|��0"�"O�����_�,�<U���=KȞ�W"O���B�K���3D�[���/�y
� �(Ӡ��9SN9���Z^����"O����锕L�X��O�6�&@i�"OV`������+��+rW����"O�M�g�$(.��ï�x8BQ�"O�q��E^+�AQC�Bذ"O
}K�ƃ �	���¾���"OX��t&��  �j\2IƒHӢ"Oh�+�fH�S\)R�.ŬK�8��@"O��)��Z�و�J�mB��z4��"O�hS'��o �`�e�Y2-��*e"O�й��I����� .5�8R�"Op�+Ջ{cr1��.J�i�"O�P��M+����3鋾 (q��"OV5��+צ4��u{V�+4-@���"O�
���ĥ���0uА�p"���y2�M�P\ph��Տ'ot� ��)�y�h�F�vkvg���� F�M��y��.5�@cA)�T�U�Q��yr/DpBQ!�P%:ěĦF��ybNL:.2��AD�;�4����(�y�C�}��x�-Ԡ+��y��*��y� ,�j��H͚y(DmAࢀ<�y��	}�d��.ԢB��t��$�yҮǨ �����D��4�&�#�o־�y�A�<���Un20z��6*��yb.ނB�j�؀M��$
�)�壍��y2�A1#6� a��2�m`E���y҅J�?����:T_�hpT��y�G�+�ީ���QD�t�S�V'�y�%��c��,8�A�Q�d�BC��yb��jc�D���F�إL�*^�L݇�3�p�� ����0��)z��ȓS(MR1&@&	��0�c<Q���ȓL��0r�_��Ѻtℴ�6��ȓ �9��k�'!Ҷ"4 7r����]JL�päJ6�D�HT�8���ȓ6���d�ז�� �7�����y^	@����<iJeY��I|~P���S޺U����=b=���� 2P��[�;��$�j�u��<�ȓ�~G�|�FM�B�ݿED0��ȓ\��0HX�*5�8!�Z:y�n�ȓ^C�D]�M6y ��m�2t��Њ��.U!,Ui��`͙l�b �ȓ(zP��E�0l�QZD�Qcs.Q�ȓ%��cc�Ԣ8���IgLB. 쀇ȓ81�Coׄw��d��f��-����w~�yrҮɠ^J��sA��{���ȓB{bX W�R�xD2���G����6d�9X��[1J�L��A(�͆ȓ41 1Ӳ�ʯfR�فPH��(��P�ȓO�l��W�s���[���k��e��*��嫥�݈t��ib@�N3lB��q9d��Ӣ�j�ԝR�6?�����O�r����9z�Uz�鞗|'\1�ȓv^�8Yuܖ ���q��>XE�a��3_�a`�w���1g"��G�
���2䌡PG�=1y� 0@�A����OxZ0:񠄺�����O9�ȓ� X�V��Zu�&���ȓ!f���B�/��m{���?,��ȓK6蜑�B�M� -{�$�l���\Er�&�BIX09�O��d��ȓ|���k�:
�
��� `�p��S�? lUQCdܐT�v���LW%`}�x�"O��R�%�&�Kܝt�ق�"O ���B>JhZ��d�^�S�����"O�����b�L�)T�����37"O.�ȑ�(��#��.j���ɕ"O6��`�v��pE@��[�N=�s"O(b2gC�y�^���˴��c�"OV�����fTb�� x�lٻ�"Oj��ªWx�r {aB��v@y�"O0��r��
Y&`�`�O�UXN�"O<!˖O�/���a  H�g�A{�"OB9P%b��`�鍤f�����"O���QKR	43Z�[���.��"O�(�����S� �V��,�ș"O<��,�:4t�s3fT?���"O��	��a焹�E&i-��@�"O>��΁
/�Z�{��	)�YSU�$>�Şk�%��! Q�&Ă�`%G����9�f�H��D�
��H��^<`|J�ȓJ�6I�#@�k� D�f$Z5M�~@��C����\0Q�2|R�ئo$,p�ȓ��)!�g
;�a��J�3Z���{4�zq���*S�a
񨔦_���:���25H�hږ�f�ڬ %�ȓ��xR��z0�7�&9H�]�ȓ^�zEUo�"�s`��$�\4��8���B�C>YcX�#����&��X�� e���\�Uj�hC�Z�ڵ��eu�*hU.CV`�K���	S�ņ� �$��OߟQ��C�*X��E��W�T ��C]�$�+�%B�� E�ȓp}h������6�X�YD�1��<��NklT��%G�8��Fڤ^<��ȓL��,����l�%R�/������ȓTe����)ҁ̞hq�ȓw�����SZH0)Ѳ��2��m��~%����h-P�Nޗ�r�ȓY�r	Qd������n�oo �ȓ5�f`�GXuL��RX�4�ȓ
4�թ�&��Q	���p��6�$; l 6.ʽ�!�I�ThjՇ�]�$�9ū�jh
� DC�z�F!��2s�9:*�
 �"�B2�R9��=����a�9^mN�x���/g�1�ȓp$�A�à>��6M�7Fn��ȓ�D��vF��>e(4����.��ȓr�vHR��L�t}2M�4()K�����ri����j׆gj�*5.�<	�ȓM��=��"�/3�5 ㄜ"+b����P�h��^yD����u[hP��a�Pp�	҈w����Z�Z���6�`���`-��f��	hD���o��]�a���]O�i��	2���T�N!@KǲK��x��OT<g��y��QX,ܚ�(ٷ<B�P�2�;����4�`�Y�bͫh̴u��9jK$��ȓyc<Lc��C&qE4��mܚ7�dy��F]~t��⑩_%l���S!�|��,�0�U���L-�E�4G%uz)��6���Յ�'3p�5 �OŶ���hіY��_.�i���]�J-�e�ȓ@�V�;�AP� ]��5�K;^ƠuG}���\��% S�G"��,!��۾�C��2nL<
��2k�xq�%Zo�$�S�O&� ��:�l�[,���V@ʫy�Ap"O2�HG.Y�}5�}�-��w��g"O�!B/�aZu:�V��qE"O�u��ʞ55���Dk��&��:"O:�f֞Q��P2�/ �4-�"Of�R�N<Z=ج�ƮU9W����"O�qH��ק3���91.�� R��C�"O�P*�E�r�����M�/B¨SR"O���3b�g�A>UA8� �"OrՊ��	l�tݢC�Si"tՀ�"Od-��'�G~\�{C�'�A80"O���A�_�O�f|�"�V#6b�Zt"O��N������;� ��"O<�B���+G-�1%�M�KNM��*O�1òc�:;��4�$��D���'�#5M�?B��\cg-� �p��'�&��FĐK�E�fa�~��'
�m(����ȻŃ��6�:��'!�����9�j�����)DH	�'�,������<�QY?1��x�'����$���"#`ߵ�~}`�'h<4�-�1v��ѻbφ%~�U�'j6���#R6�h����x�|�	�'�\a!�7d& #Cܬr�X��
�'|&�H���2[~�A��ׇS$�
�'�yH7� (8�n4�v �G�ƽ(	�'�	hRa�5xd|:��F0>�`�'S�H��SZ$DP�,_ 3���'�D���
�<X����
���I�'N��S��^��H��s&�A�:Y �'v�"���=�UqrKV+J]4}�'?.4k�i�)D�n��K�#J3r�A�'|�Yd �t�z�A&��?��9��'W��9�"&��}���)<�>1�
�'��P&��.2�i���a�8�C
�'�j�!��Z���"ӟYf�!�	�'&��3$�B#Q�T�1A]�#�.A��'Q ��j��S=�آ���&���'D�@*4h��(t2�#���%U.�OB�=E�4F�EPP
mz)���Ώ�yr�_+A+�MR��DA@ `��Mc���s�����BJ>'�ht���B�* ��C?O��=ͧ��'�<uQ6�q�P�f+�4D����'#�����bf���bͷ?ڄ���'�,��)ħ��e*ֈʻ/Y����'� �fڊ:��z���8+�5��'�j�(g���Xl��|�xhC�'�
��u�0PT0S'��w``��	�'�$1K��(��*��t�䄺�'#��S�&�M%�9k-r��8��' a&�q;��S �"����'����u��u��X����/+��@c�'��J�O{h�rb�U!s:���'a4}�r!ղgʠ�Al�?kR�K�'�	0G�4R�쬓�Ņ1ct�Ȋ�'k�Er��>~#t�c��cɦ���'>M���Ɏ��i�E�M�a:���''�,QB퇨\M�@�Ud#W�Y�
�'z�} p�N.���c�<u�2 h�'����OJ�{F|�q��0lh$%R�'� K�*(%��P���L� QA�'�Z��V͉6E��C���+E�4�(�'�NT�ī	 )Z�4/�9��y��'>0�A���9�Ĉ�4�jdR��� Hp�e��b����"Ԋba,$��"O����� 4�AO�f�SbH4D����F�L�����Ν#l[� &D���g.<�Ќ21��
�f )b- D�H��Ē�4|إr@�� �H`qB�0D�T��ϤO�4��#Ȗ2���f4D�X
��g��з22ʺU1�E=D�x
�䙈}��yĊ�"�Xta�9D�XZP��#G�HKa��}�X��S�!D�0�0EG���Ȓt� �D+ k
=D����ʹ��=��8N�9�vF:D���&-��'b^\i��ӱ8"p�q�9D��y	T&60�0��������,D����F�X}�G��e��E�D�6D�`���L�X]a&�A�!he�6D�� �E"QA�Rǂ��hU3�i?D� RwgɆ�����)��� �(D��	1�٪ �1Xb˅W�}(3�1D�����)UKJ=���M܀���0D���m܁D�L��\�A��QcA,D�����SM��Q�af�	s��K�/D���6�]t�4a�c��H<�b��+D�`�"�L�5T���a=?aeyш)D�l�'Mؗ:�ޡH����r���Z��%D�l����D�ε�P��	��,R��0D��YB��Gd�L��D�wH�8��j/D��r���4ݡ��	h$b�b D��6���.��L:@�]54;j��=D���g�`DH�%�xB^h���=D���h�?Q)8!�D�>tl.|)�/D�h3a��ᨃ��Sy���.D���ӤM&�\����K�����d,D�ܓ!��O&��@��)Y��q�r./D���FO ��c뛷Ԓۂ 8D�4���r��Z;0�b�'�#D���I��N|��썤/4hw���'�v��6�zС�!эFX�Q�'<�D*�o@꼲�	�' }�$��'o8Ң�A�+��%s�����'�,�� �×;✝Zt���n�|�S�'W�ZӦȡo��l��e��b��Ѫ�'�@PšB�?�V�肄D�a���'�4�@���2EcV��R�<8�ʓ ���T���x�Н+Ve�(M���ȓv�#W!��*����r*^�|d���ȓ/�2-j���c~��s�<R
��ȓ>P�x{ŧT<D{��� `U�P4��ȓAs4Q� �	���m��E�7��]��s=�Ѓb���S���GjG�̱��Fd�*W�W}h����cX�w^���V�Q�ţ,`}����
��G���ȓf��� !�)�,�R�&� r�b��ȓ|8������XԈ�)D�<9�xT��9��`�-S*Ф%��;~oF��ȓi��ʄ�?K(�@Zgo��v�6	��-uLd��D#'F��6�m@Ƞ�ȓ��h2��H(k���)'FE�P�R��2�x�)�5��4�3�D�r����ȓ,��;6��5��P�Ŀ$����ȓ��5@t����L�;��a�ȓh�T��$8+��}(�� ' "фȓl�S��H�:16�Ip�Ɇlj�Ȅȓ/%��7��9{����#�I2���ȓr��<�0���K�(Ӈ�=8�=��S�? �$��Η��ԙ��8e�^@+%"O�A��!#ܖ�D�@�x���cV"O~�������@��l�c�"O8�aH:����#J#c�EAA"O�-q���P���Ӥ"
	pm�"O(����#j 9"���{���c�*O�Aq)ĩ*yZ�*��p�|���'����d�$U�j��w#�eF���'�Z<0dU�t~���V�8���'�`�zB�e0~x�K�	N�B)�'ڀ�Z��	�h4|����7_�X
�'��3ҭ�.@sR�F/F�J	�'I��;g�S�o�T��A����
�'�����#ʴh��a����>���'�� �̞a�V���E�'CHT(�'�İ�#���PB��A�T�N���'�T$���2� ����#X.�,��';�lR�KZ0 ���1�TM��8��']���u��9K�I�F�C-��'��)��lLz�y��m�>1t�
�'
 ��a��qF~d���
J4d���'�"͓vǕnF3AK�n₝��'�0�q�ٸ~T>݁0��!0�Zũ�'W]C��4@��"�T#���P�'zx�`t�ٹ_5*�q2��7�5��'���Р��>X��Q�3a��'sX���ΤC�꽁�=9���'"n���G�]��� `�Z�ۼE��'= ]x�/�>�8�"���z\Ƽ�'ܑ�PA�N��|�i^�j.�S�'��8g˗��$C2e\��'},��0�Ġm�����h��Q��8��%�&��P�R9�ĸI#eВr��ȓP�Q�M?�Z����\��&�⸹�ϟ��~�Z�*١D����FiF��'��V30L����hs����KlbK�AHg@�D�V��/[R�P��G�1BveC�:.��%j�^����ȓ�ƌ�	:���)\�Xv���I���bC�>�L<`��H�P�Lp�ȓ4x��%iܖ6�h=����Q���x��1Sn�j;���� �n��I�ȓ>���!�6K]�� ��P�C��d���������d��ӥe�=�쐇�1�MR� ���䄔
����[�*�@5�ʘ-��H�DKK�`DP@��4��x��c�2�hgAN�J��i�ȓ�n����W�&3�ݸ� �"2����P.��3è /x �x�II� ��l�ȓWHB�k�nu��� � �Rk�T��q��-���W5y[<�j@Ë.<Ѕ�c�J��a��)T0���n��J
��ȓN�X����9lږt�G�YDM�ȓx��Ps�*�i&vDz�C�?M�r9��b9*���?�ĵ8Ap綈��j:j@Ia����,A E�Z5x�t���d��P'���D&��C�6p����ȓw6*݉���B$�س���a�"%��pv�Ցfeеa�(���-'���ȓ
�L�*����?�&�!�O̭{x�ȓ<�L����N.j�>�!��T�m���2/Ftز��:V�6p��	P!/�`�ȓ��
�<Z�#��*PGܖ�o�!�ā�$j�s���(��!e�!Wj!�� ��+C�F�j5���`dƂ<29�"Od�hW�>K��E3���	+&��"O��@4gB2����7lޅjƼ�"OҜلA�ki,��U"R1|��7"Or�t	�e6�%	G�ÔN��{d"O�05,�31�+Q�[1����"O4 K7�Z :UҮؖ�RS"O����EY(?�D��2���m "*`"O�@8�b��8,��[�@L�lg�4��"Ot��D���mS4b�>KJբ"O��QՇ��C��U��*O2^}�R"O���t�ͬ}�d�e!�?j�"O���_n ��mE#z���s�"Oʱ�s ��b�E�6m�!0��e`�"Ova��I.p<�2q.�0�T��3"O��{�IB�I�\PQ����)F"O&��ĆM�i�X	2�)7ʔ�@"O�b�l�3��i�@!\�i� ��a"O(؉+1lj1���c("�"Oe R��2&�T��O�*=�v�[�"O���φr`���	�%�Ne��"OnEp�$UPz���N�8��2"Ot�����#.�6�� �T����"OB��D�&z?*���!�)��m	%:Oh�7�)�'j8H�耩Oĺ}�`�<
t���j�m�g�Є�4P���w�4��(�؄�fm?|l����ПE����ȓ����a�Qw�!�1h�!;c4��ȓ<���/9�Ǭ9Db4t��<��{A!�/j�"��S��h�ȓbBpL��V;W�4���ڭ1�X���Vj�S��,����toO�d,��'iў"|�V�_�L��0�6ꐆf�*|���D�<y�F�=H�hwɉ9)�l���~�<iVI�(�@�g�.�����*�y�<�O] E6f��-�3�쀃]u�<9�O�0��Tʁ��Ȃ�x��Bn�<�JP+vDq��l�|����~�<����"7 ��Q�� n�����@~��)�*O�H%��=&�5�ҧ�b2>Or�=E�d폼jN�����BQD��n�<�yR�Dļ!BęN@Z��v��/�yb�ݡ(�t=��%�?5z��{c��&�y�DE�>?D�) ��3�H$�7 ׽�y��E X�T�&�Xָ��I܂�ybF��/�\=� M+ز� ����y��'��O1��˓TI !�)X��d�qa�aI6I�L>)(O1�1O�MYNW;x# ��;v�h�f"O�AB� G0��@KAl�5ln�"O�d��.A��D��+�U�M �"O!��fV9?sF�4�I*u'�0ч"OX�s5-[��2��F�Ӈ.)`-�"O�m N�&��d�%��[3�*��d6�S�'�9i����\H!��ǎtf*YEx��'����v��A-b4˂嚅T|�R
�'�<%i�àP��7��{YҴ��'����`��oW-���w�\]3�'SPa��H?F�x؁�_�B:JDk�O�ʓ�hO�S7r�h����%j�>y�M�]�B��>r`HB���Z}����6O��B�	�c���b_��,���H)��B�ɟ�L�r�i�+1@�#�)��B��1W$�H�RC�.	��@FH.$��B�*	O�!fD\3Z�{%���lZC�)� �x���H���p�!�5�.�pR"O���_�$$���ᙬ:%F��"O �@@C�A�L�'@ڬ!
�h�"Oh�:ab\5{�XȳS�6~�D93t�'�ў��`ŚTHz�9�� �@t*OF�������
�B�&�Ʌ"Ot�34኏Lr�P�mI"O`q�*/y؈��֠G
z`"ʃ0OĢ=E�d��Ia΍����&|	F|�qm��yҁ��ीǫ��v2b6nS���Ox��p��|��BMX�N��X�B����C��1_p�ɥ�H!R�T�6 ��)��l�ȓk 4����Z�� �7n7Ol2T�ȓ!_2I"����UY ��2�6P�L��X�V1�ch�]~h5B�@A�$�T��O�����톀J.b���C.1��ȓ�\��	�8��Y�E�2XF�pGx��)z�;� ��ޙU���(U,�|��X�?�$�+׺�!��� 9mt��&�}�<�&��		���r X7�TMH�b�|�<�s��F�SffBL���y�<���}~
�+p��mH��j�v�<q�l�E$r��d�#s{��ɷ/]�<�4���V�'H��a��y!�C+���8�?�|"�!_�&�p�$iP�M˴R(8D!�D�i���WM�3ۼ=�v�L�%!���,��a��K��Y�#�j!�䆆?=,��$y��˞X�!�-w�`x���5U&t`d��DX!���^�)	bM�&X�ck�S�!�J#xR���Lhz@��n�!��<����R��ZnX	ҡj��6�!��d���{03��"vY�:C�I"<=�ux��!�
xc�N�=u�C䉎1(h���тe��%��6N�C�I6��q�t���/#��$c^�u�#>����BLl5	3O��o����ך7���G�-��dP����'D��`��`��y�X)-��K@/
�e��5��4�y��8U�)aeʅ^���8�f�=�yb�)]>x��,��� Q����y򋟜A'q����0W.`)��$�yr�>VUB�P C7z������O���h�ܩ@%\+Z@V������?`Fy���'���d���>��V�L
'fD�KÂ�d�!�d��}���*��ћxR��h����m�!������t9��S�cD1H^	Y�',�`�\=8 D�tH�{RF��'ծ�c�k	%Nz���Qp�� �' \m!�'ؼ�v����_Ř�@�'�8$���tE8Q���j�h���"ON�� D�~�NP�B�\�I�7�,�S��y��T"*���rd��x�ę夌=�y&Q:T \c#
F!n>�����yb+� L�B���	%Z���+#����y����0Ft�ѷ̈�ZB|l+3�R�yD )0�J�1@�[�K�Y�w�.�yÊ�Z�a���{��1S��T��y"�M$t�ex!��s��3�C֬�yrm��0I0'^
_��t�G4��'c�{�.L0N5b	�!���V�"��tΎ�yAA�F���H!�<�Hۣ#	��y�ϙ���Q�5����C����y�
�-pL��w�%3$p�ASiB��y
� ��K��[�M4ƤS�DMqSd�1e�"�S�'";����6V%�͠ �CBT�Dx2�'�漺�&�%j��#�\�	�X	�';8y�Ůǻ=��p`2�	�*���'Ԕ}��ݖmCj��F6A���'�D��Dѫ*9 �1�H������'�:h23��K6r��lʀ t��'dlQ���D�-~�D��'X+jp�I�O��=E���̗$h "�ڨ"dP1�O��y��+/��32���w�K6����y�#ґ�v�b����!�A�&�]�yBh�,[�d��0�$?B�
��K
�y�&�G4ȴ����\ة@��P$�y�吱M?��8#J=P�x�v*M��y�J9�.�rB��JS*P��J�1�y�Z�s���@6#�z�h)��7�y�	��8(���yTn8�%�
��y��%/1(�h���5c᪱X�,Oc���=��VYΘ��!	ӂqa���C�<a��F�L���y$҂5�J8�$ME�<Iϟ3�x�C!�7�NyV�}�<��/B�	��1�bO�9X󮅊@jx�<Q���9A�n�B�X6`��q
U�w�<9���OJ�hW�Ʈ(J���׫�K�<!w(�99xH��b(���@��
�<Q*Op���J�C�UmN�Y-v�9���0�!�D_*��#��B�=�ʄHU�z!���A!�i�&�<c\b�"�o�8�az��ɯ}�`����Ip.I���ZP!�dP�O  X�B'��}\�t�4Ύ$E�!�$Ⱦj���3Fa�nN0��Bl��f2!�798�qI�����`�##�T�@#!�$�-Q؊�:P��s�8�%�Q�!�\����ӇC�UM�M�1ce�!򤘺~�*�� �uJ.D�� V}�:�O��p��G��{��N �P��"O������|@�Q��b��J�"O&;�)�!y pQg$����Mie"O�P@B�B���Y
�BS{�x��"O~�c"+��Fz�I�b�%rxA9�"O�)��R\}�E�P��"O�ɘ��߀p�x8��44F9�<Ov�D�Ox�"|r��O8fZ��$�&p	+ �I�<�f�C,;^l 3��kQ^���L�<1F�y���[3��O�fyQ	 D~"�)§T@��vB�>*j�p��j�Hs���#��r��S~\ȓ�Li���ȓE6��D/�!G�\����O�py�����?q��ޣL)\���:cK29�-Pf̓�hO1��d�5@��"Q��,� `"O$H�b)�>��,�QC!�x�"O��p�ܳK�A0j�?7j�FF8�S��y��2e��q��Q�^�b0!�Ő�y2	T�t�.�$��m����I�3�y��#Q��@;F���n�jqK����y��=ht� ��m�� �V
Q��y���`M
.�֔�'O��y�C2��|���	o$�����y޽:fԑ#�P<6o�3D� ��y�)�'7^��uFʮ_��i�� Q)Z����ln |�G�]f���ۛ6iX��ȓH�E*𩂗r��%S��s�F��ȓ `����S)/�
T�s"�tV��ȓhx�)���)N�F8z0j��(̆q��S�? �1p��3�d}���X=hU>���"O>0���1@��1g�h��1�"O�="qAW�
���C�F :�0l��"O��V��p���@( �~����"Ot	p��Hx�#�ɷ�$�"O��B�pc�'Ũy�~�z�"Oz��aE�}�~�2'ۚI�2�qT"O,HK���P�B���#'QĨZ%"O�� ���EٚQ�p%��(��'�Z<"�b�3_�ఒ&�x���'���+EDD�`���v �S�'�vP��C�.tP�ˊoe^���'�0p(��/-W�(��N�vx���'�����G�� ��%hƌ��'ł��e�%�f@�����H ��'�\��	1<�p�+a��7'�5(�'k�=�"�Q(T�p�#�'ŐF5��'�I���ݪ8�| wn&-��T�'%�:��`l�k�h�O5L��'O�5� Y�)^�L�P��0��
�'�X=K��Հgl���dP�%���8�',����j���#rAU�!��'�"�sv�x5��iB�$*�K�'tj��AQ�Q� �`Ro�� ���'&Z��1��*�.�Z�b0"�q
�'�
y��8Z�2�$鐪b�`�'�H�vl-rP:��'��
���	�'$�XqBR�~���GՁ2Q��'���k��Z��eʳ���Q;FԒ�'�T��Ȟ"'�8��n�L4H૏��(��`��W�.�,��tAɝ.��A�"O̤J��X�H�Ųg@�t��%"O&m�m��- "�9�)�*IY�"O�E�pf�;�6��/[�BHK"Oxq�˳m6�a�ǋPڸ�xS"O�t���Hv?
iqw��)��2�"O⼺�
MNyJ��t!ZSH�̪���K����J�e���O��Q�q7#�4O!�Ĉ'
7��a! �V�Z��$#f!��ޝ�P��� ڱ~��h�a�S-Q!�d�k�̙�RiQ�fji
e�V��!�$5>�4Ԣ&%^�K6�k�.^�B�!�$��X�(�K�j�?0�mf���/�!�DV�!�Eq��Ń
��D ҈�)���G���D�%�h�b�G^�+|��0�ڒ�y��Љm��T@Ģ�}7|=��d8�y"씭8 H�D�o㎜��O���y�`�/R���#M�kbX@��.Ӛ�yB��D�١C��c�h4#B����yb��d U�e���V	��HA�P%�y"�q�
 b��[i��Pऌ���'s�{��4Il��W� )*z�*���;�y��P�[j$@0�
Y���ĻbÕ/�y¦�``�KK���A�Y��y2���6�¸����yH�/	�y���wRU�Ҋ��ulЩ`@W�y"	0��\��f\s��店$��y�!G/I�DB��Ƚn>\XAWF
��ybj�"��KBMJu�V�*��ǽ�y��3 ��j�܁k���Hu���y2��CD��H�Ɲ�yd�iC�K��y�
R�s4�4B͟�r��V �/�yB/_)8�TQz�IF��%�V�B=�y��jb�3�.�qR�QH�)��y
� 9�FH7Mݰ��`O�3���s"OR���K�إqp�֠QH�"OV���F]�F�` p�J<'��}9�"O��&��A��u8�o�W��!�"O��
�&<QpލY�NH#VLq2"O�%jv*�3L�6N�>j�ݡd"O�))���N����M�\��r7"O�A���Pfp9��+ �|� ��2"O���K�B	R��k�bdFA*�"O"wƈ�H3Fl*qI��=RѸ�"O(|��Bs�0���X<&�-��"Oȩ�p�:��4����P�X-"p"O�ͱ"��N0�U�$t��t"O
]� ���03�X��j��!"O���,�9F���f\+[����"O��B��1\x�h%�D/oR�q`�"O�D��gA)�tj ꓰI���"O����Ғk�
�	��+,	�"O���A�l������+K����b"O��:�
�g�%
�J�k��h�"O��$,��q��U���ν~<��pt"O�h���^�K����4M>Llk�"O&�2G�6���CY~�����"ON5Q7NR�&�B���E�����"ON��t��}V�ى���:B��"O~)�D,�^���$J�7z�� A"O��* $��c&>�UD )N���"O���F-PޜYǣ�"H�1�"O��
�ΤM�
	���+``I��'��'�T��,ޮ�����
�$s��	�'��Q�P��>6<�%`5��$����'���c��:T�-��t�A�'jĳ��3^�8� dIO�s���'��5��˰_ѐe���Csy"��'/�]�"ؑ�	
8#�bd0%�?D�,(��X�yh����g�R���>D��8�ጛv���W˟��%�Ռt�!��)B�Z�h�$׋��@gQ51�!�Y�qP<�)�ꕽ8�0�`�����!�C(a��)�C��H2)#�T3`>!�$�);��i�.�)3��dѝ"!���0+�\a�.R� ���i0b�04!���Y�t��o̴#�|5�f��D"!�DT�3$>�H�	���	�P�F;,!��Ġ&�,��OA(���FY�^W!�dY7O�p BM���E#P�hF!�D��#�� �Ē4�������9�!�dS����y�E�4,�:q@�L�hl!�<`�<���J.�
�f@�/P!�O�Bj�X"�(�u!$�����!���$Ⴠ�ȽF���I3��?c}!򤑥y�pRׄ,�ȗ�U9�ٻ�'񆁱E�'[�@\���M)P�Py�'�|��C��4D�}yt+&G�fl��'0� K�(��Gv� u#@F���'�X��j�?��`�a�C�0�x��'N|գY�
!A!eK)y��|��'�&���E� >�=���MjB��
�'K��{��I*S�l ��,�j<��1
�'�@� �@��� @1`�dT��'=�5���7uw��3�gֽ]��H��'N��E���F�\��ER�Iu��K�'�p��fJ��X��	�9w/�E��'P$؃ �5?/$��sA��uQ�݁��� ��4�
,�I�� ������"O����41}�%i� j�n��7"O~�;և�zJ��o88���ת,D��XG�2�p�ˢ��Ae��E�6D��1�*�<9,� 3�N:
p%�`�5D��z�"�0*j �ew�t�#��&D�p�!�S� ��	�,V& ��d�:D�8�&� (_D�I����i���k�o7D�܃�i�7*V�J�nG�o�΄�'o(D��� &Thf �)Ө� i�\���c&D�l��'��R3,���d �P0(*b�"D�����#%D�T)Mʙ3��"D�4r�&�^ay�b͕s��yA�H?D���P���;l�s`�E�R#���3� D�(Rw�O<d�x))� �=ײ� �!D��8(�.Y��ĕ%}�b\y��>D�`���r��P[w�Ŧ=B��m<D�Xr��T	��x##�$okf����8D�����Ԉ\Ҩkd��jv�j�"!D��x�IYu�`��P�'m\��ю>D�l;��O3�z�"�#ʨQ9X�إb;D��hK�l� 1��HP^ٚ#�4D���c��={
T�dح8�Ah��?D�p;�a*N���Uo1a��Ag�=D��D�>�����0	��i���1T�x�e��=�F��UE�WB�Q�P"O�d4� )
uْ�݌Aᚠ"OJ�Q��G�B���Ҡ"���D"Ox��Kٲ]�Pi��L�35����"O,|1��D2,�"�� >-OT�X"O~LBBH��x��L����-5����"O�exP�N�)[�{E���+ ��A"O2�pR$��B�H���}���A!"O5Kt�X�,D<�!dɜA�qٓ"O��q� ˯E(pٓ3Iݞ85���"O�d�(�*MS<ш�*�nN��"O�	�h N�y����\ A��"Ov"A��;���዗�x]�Ms�"O�����2Z=��IU(\θ��"O�-j!!V1t52X05���qV9S"O.��� ى
��h�
8Pm"�"O"�(g]%@�X�A�;K�d�R"O��Q���toN����W�_a|�q�<1�7[H��2�t��t��}e�m�ȓYm2��ԠT�l��5����S����^���r�`L! �<:0���rY����0:�����b���7�y��K�ҝs ��gu��a��2(�f|�ȓ]h�SӁ�
W���A&B�-�0��ȓ(f6IQpʹ�p�̀C?��ȓr��ES,݂D���@Q�E4A�"8�ȓAƪL�$��'!'PH�e��n��d��\��ࠁH\�p�T�����T�lф�+%~H���.��8�i�?&`��;�|�K��
�����_�C�C�
�~�i�M%�EcBeh=�B�ɯEq��#v���$�mەR	ޞB�I�uܚd�s�i��%�%�Q:$��B�I#&8U���	��kiݓ'�RB�ɥ<H𼠀����P����30(B�I"b`pE���ޯi���ȕj�G�B�=Q.��R��H�'�l�� Г+N�C�(�>E�&�D�nl�=�ª���:C䉣t��	g#�"y��Kuɉ�5��C�)� P0��� 0;ZH��&@�2�"O����[&��g��4PT�P"O�)QpL�`@:�)�_�@���"OB$c�ł�+Z�!�Ă��A�X)�"Oj����@���b�₵
���"O�� ��zƒ����D�D��2"O��R��`��+QE:�d���"O��c��"�A��ʔ]�li��"O<�*j �X���C���"�V���"O��K@� cp�m�"W�ʡ�W"O��x��T�{�"+E�ܦ��"O>���	�f *�[j%�L��PF{����/^xH`��	^>w)�*V�F6	c!�$/Y z\!U��_�e���6a!�V�+`bST$�
IT!��e�!�vf'�̫ *��!�DƐ2����$1����ds!�D4f���!�#��&άBC��2a_����W�O͐Yy�ꁧH"�`��ҕU��y��'�|e��@=�h��=�Z}����8<O�=��I��H�^Eo	�m	|["OH iV-͍'�b�����+�P��2"O̙�0($�ܨ ��H93�F��5"O��fW�$�z�hC���Dͺ��q"O0���S�L(8@B�/�t͘��'�ў\��MA��Q���B�.xQ[�e�������ؙ:�r5H2j�m*�y���-F�!�H�G�n��(%��,��D(T!��[��aBgǄ��H��&�"I!�dì^�X,��o�"1Б� ��?o=!�ą� +z՚��M3 �8��G)�X5!��
*�̔9"��y���PT&�#�!���^��I�J�^p��a����1O��=N>��JY	Sj�1(��ܘi�-��l�8�?����җMZ�l 6c�}z�����
z�+΃8���V�ȌK��ȓG>�A���6��ҁJ݊	j�����H�1}��c4hF�V���aφ1+��.`���,�6-��0`���ԗZ�Y���^�V�N��ȓu��-���(d+Q3�z�ك��<!��T^�q��
Z�*_�d�D|�ȓcH"]âP}-8�`�g��l����)�V�r!��"L�i�b��ЅȓD��׎W�t\�/����D�ʓT�.ku��=@�P
�'d�*B䉉sJPidOX:��!g��cR����<1���m;��UAȺz�<8cU�HH�'��	y�O�\�t���b��]9��O�����'�����(L$R������.L�ő�'����@Bj��
tK��7��	�'|t�"iєlv�qsjS�(��U�	�'�0!*�>���P@�Tj�z�'Lb��4A�{�6�Y��5	8T�'Kўb>%�';����^��!i#�3���'�ڰ��
R3rz]T�����"
�']~)��
Ӫ7�����8���'o��U��B�!#e-yՈ��
�'\.���J�dl�	x���o����	�'ԍ� �FMZ���i�de�,i	ӓ��'�A:�� 9v��b/��W�hI(�Oܢ=E���]+F#�Q�Ε=&��TG	��xR�'�|-Bǩ�W�L5�Q(Y�F$<�'$�,SG%U��b�y��U�8TR�;��� ��(
%;*,�b�!-vX��G"O��S'�0J��@��Tl��A"O���m"jڝk%Hr���;g"O��ڲLĬb�'6�����"O�ؐ�F�fM��9�L��oT�P�܅�	!Q����f��S��5���MOh�C�	�_
�M:�F�$|	Q%፯��C�I K�|�ǧ!9Z=���`J�C�	�*J���D������Y�mF0B�	�U(�l0@���X��I�,r�&B�ɰU�<���� Y¢��#/l8B��<��+B��l܋��"J�$��?������/gD>U3��G�R�y$+�ip!���	N$	C��Q=q(����J1H!�Dh�p1�B
��2Pԑ�DV�1!�$E�GfE1�D37k��7dT#=O!�$�;y�$��HؕL\���!��9!��p����Ѫ�E'b4K�j 'j!�����Q̉��̛��W/= ��6�$�<�|�'%2��'H�0f2Q�P M�|����'���b�@��5��f��t\֬�
�'�����P�gĄ��'$lG��
�'t��W��^��FO�8�b {	�'�F<�-�;W]��Q�@�������'�V�;���A�0i����]M����')fT� �D NI8u+�'��S�)�<aWJ�4+�Ú�hS���D�|�<�䡎.DAČ��)�� �e�R�<��h�60�.�*E,�><��Q�"�O�<��&ګ4��p���7_J��᧝q�<��t�
���
�2��yT�RX�<Q��[�"~��Z� �.e���Q���_�<!�ˑ"_��B�ś��c�g��<!��Uju��C����I�bO�[��݇�k����S��n�D��4E�ȓS���q����DEQu%�<  Y�ȓd�ā���E��Z3�6A����.Pl���O�N���;�~�����d��U�	 G�n��Ћ��2�� ^�n��C� W/�ɢ��$R8E��@g?�C�	�
$0]��>(�[E�-s7�C���LqJaפ[��e�cЁGbB�ɲ�
�B���
	�<KP$�<�xB䉗E(���#>Zk�9W�~5NB�	�~��1��� z`s�̼ �B�IF�`3�
$�H0-Kj�,��'�IH�)b)O�a�B�M��K��Uc��x�"Ov����E� ~����40�Ɋ1"OnT��*�8@��g���h}z�"O��	g�ȿ^y*�҇L#V��-�d"O,aA�
�!;�A*3L9�2�Z�"O}��!��ЩB�q�<��"O�Z��ɾ x�<r��Q:rX���.�Ş!�Q��4:�DI9BƖ1<܄�ȓc��`��d��&�����\~��_Z� ��ʶM�1����1�ʱ��%4��ELިI&"ɘG���f��r}���w��SΚ}x�/�)�|��w#88��I.�$��H.��T�ȓOW�l	C�Ҹq�4ᢟ.6�֍�ȓM�F�A���d��� ��^�w�؆ȓQ��%�"n�!�]"�؆�$+�$ó�An�	�F�n'�P��A�P`�>Zj�BP�Z�G�!��S�? �ՊՊK4n��2e*�-x�2Y�Q"O.�1G���:����F={��L2�"O�Ѻ�Ă���ة�M����7"O���s��D~&B娝.`�久"O`t8"�CS.)brFɏ�<ɤ"O�y�Q�]�!��P1Fؠ'bH �"O�]��EY�Q��/U���:�"Ov<`�e��d�x	���ȕU��{�"O��YcC�w�<"����.���"O��iU�^7!v��je����"OZM G�
`�@��g�<-V�`�"O��x�	kȞ̀sώ�L>�l�"O4��W
�H4�,��蟘3�����"OmBͥ;M`(��7��a�"O�-J���+:D)bI֋���"O�p��ؓ(ȑ#6HȟT��7"O�Y�#��Ě��P��0�8��#"O:1���2v��I�Pk"O�����>S����Ɓ�1��%Y�"Ov���eƝE(\cF��H��2"O8�Ⅲ��Ј�K�#$Ԝ��"O&��fG !By���F� �Ai�}K"O�(��¢���g@.~WN@��"O��!���+瘵�� ��Q8D���B�O���(��<�|ΓRl8��f߃; pb�˯F�p��>:��چB\�7�D�;����,T��ȓ��T���V/r�\�p�)�*�ȓO�,�㋁ ��ȑe��HH�ȓn3�͒�
r��٘1� G�������P��CcP\0�$��	��`��Sӌt1k�+��M d�1�x��<a������O����j\��.I`�ȑ�d��L��'�$-*׀G����l�	Z���'=0�yG�?1���w�LKl&�{
�'@��a	WEtU9&`<��c
�'��А�� �ld ��-Ӛ
�'���b��
����A��@d�	�'\<��D�6i#h���+L��d�S	�'���hξE#�̓2E " ~J�[	�'Q�Hkn�-�>�K��_&E�1	�'��\ �+�����ac�����"	�'�"����J=Zx��ra�
$!O�I��'��Ջr��>g�X���ɗF!��'q`���h
�]�B�ڦk&@��'��͙v�^:+>��![��~$��'�� rc�T�� 	��<u�Ը��'m�e�W�_Nq�-x�AB&g�8���'�����F Hȧ!ѨZHti3�'��h��ڵ\By�r)ݷQ�^�3�'1��B1N�=�����	�P���'~NiP2 �E�B(�c&6�L�Q�'��"���;~�!"�+S"����'TE˖�B�r4��M�eTa��'�bp!Q��YT�H���.L&���'O��!���5e�6يA�B�*�!�'��Hc�ڀ!A�=��  � ��Л�')0�a��)�웇h�f
@�	�'��b��ɬ�CR��}]�p�'&����K�T�lBq��"+F��ʓIN��0��	W�~hؗ
�Y��ȓN���$+��n.dQ8�W)I�N4��,� @�6�J�<�Hb��"=$-�ȓ�t���j�#BH��e;D���7��y����vF^#\On�h�=D�� �	��@  �혠�ۿJ�I��"O�jq��6�5!TG�qcT�e"O։У��Fvl}��L��7H�<IP"O�q�B��L�Up�ᙇ)h�Ep"O�̢�M& ��@��}�~E)�"O� ���҃���sn� Y�E�T"O` )T��$D'�=�^
+����"O���d���g�<mɑbS�-<��
@"O�]��JW�]?TI���z�� �"O��!sg.t���0�^�x�t�)�"Oڅ��ۛ9�bQ$���|&(A��"O��9G��@�"H�w
ե0݁D"O���A��1iV�i��h,8aN�b"O-ӄ	�[wt�AW��MD�|�"OP�z0� 2TF8�&ߤ*V"�{0"O�H� �\�n��MӁ�̝��9�U"OҬC�E#�h;�ޥD�ٺ�"O�Y�&&
�<�$��q$[[�a�"O6h����l6ڬ1�c�8��<A5*O�<I�M�A9�칤�}@��
�'tTa����8"�С�%+�fe�*
�'4r��ьV��]��H%d�H	�'���L�xJ̐�\��`�/)�y�FG1'1ꜘ�>��@mF�y�.s����C�* ����n�7�y��ƲkP������)!��J'���yh�3�vГ�V�sǶ���B�$�yr�Ȗ>;�@R���[��g��y��O�>�V�8����F��|3n	�y2�Q�j��7&R���ds"����Py�jʬbj8��$�L�
�����{�<)��3`-�=�0� ��� $�Am�<���U�6C��e�p׋JD�<��P�1 N����u�(tH�~�<�Dmً!w�P�ǥ�`t΍ �ox�<��N�KT���Ȋn��	����s�<qF��)�vPta�pU� ��q�<���[)Ą�it�%��j�<Y��=hA{� �X09p,�g�<��ȑf�l2��7͚1���Kg�<����%Q/̴��N�5i���!�L�<�A$�!Gq�4YQ��7bfX�*QG�<w�rM��p���AΌ�� $�|�<	&˕�'���t�I?|�ҕ���[T�<q]�_�n��Rd'��¡O�Q�<2�bs����M��?J���	w�<0�I�e�R���p�q��W�<��A��17��s4���V9�����|�<	���AƑA0+ٱw,�$ۧ��w�<YC��t�T����-+�`�d#7D��2��+�������	t�ZcC4D�X����D �硚�9ef!{��=D�`+��˽Z�0��ț�)�*AX�-=D��ӣ]
�جKs��	�"��B7D��3�J�`��C��T�*0yu�4D��y��7�Lmh�.E��t�4D�̨a�ʳ B�3��<V���v�7D��E�dA|"�d	�@�
��)D���1��٪��������|�b�%D�lj�ڪ$���6,�3r.�
�N.D�@*���N����(wx�[t0D�p�Bߺ8�"�P�8i�n�AT�/D��yW&Ӄz���7�Z^q>`{��:D�|3`���|��\H'�ۂ	�dz��6D�� n4�f��XQ8SeL̽R�a��"O�dA�֢z�8�6�]# �Da��"O�l��#F7w�)ci�;V�� �"O�%p�����\GȖu����'�x���Ğ��4hL\�X�	�'XNuӳhۓ>xh�3��#^��3���*��!Ԝ��"ɞB
H���1D��B��2t�L��e�?%̊�A�*/D�bV�ʯ}�ZIR�֟[S�(yT�+D�(�6 ˺jpd�b`��v3���6D���"Ŏ�V�	F��u��4�g� D�  �F���Q!!�J��s��=D��A #	/6�AZ���( ��15
)D��R� .�h�CBI ʦ�R��$D�����Z5L�΅XVn;&Y�-kC�"D�\���
7�Vh{�ꉶ�PJ��>D�X����0n,�A����#�j�D<D��@�H�$���CCO%Ƅ�d5D�T8�΁�| �Y�g&!�hhP�4D�� f�Y<]��(���)1�]��	2D��jg�A�t�hy+�%	f��%p��<D����$�нb/;�%�9D��h��#9Z�P��&D��H��1D��ǁC�z��\��Tr����D/D���TAE#l1��s��ˍV����ӊ(D���m	ig�\����!t9�����*D��i#DA:&[��\�E�N��*D����H ���� l��L"s�,D�4q�f7)b�l�����u�֕R�+D����f1�Y!!hڋ<qޥ�v$+D��(aFV���EZ�%̈́�nhx��+D�����H ���Ġ*UNؖ?��B�I�'��yh1e�1)B�|dDם&5�B�ə �BH*Ai҇Tq�h�4�S�3hpB�76j��ˠ���2b$ۀi7bTB�	v�*��-Ȩa� m¤�O>(8lC�I<x���%�$\�B���)�B�,@k�db��6�� Aǲy��C��	^���C���M�ܑ��#�s=�B䉃t0!k����i{#��L[�B��z���.���e��DEm�B�	<v��M
�D �pda��rB�	�Uj�A�H�I[~u[�m� 8B�&+���!	�UaLو�f�_�B�ꤜctiB�Je,��6)�&<�C䉥.�`�F �%���DJUKC䉄|T���E�]$�H��4�B䉢O���5HK��<%h �"Y�B�	�2>l�26�N$�B�!^�i�C�ɣz@��X�S�*&K�7I�B��m�Tl��f֞	���j�
K�c �B䉽X�8��V/#��I�V�ʟ��B�I�G�����ND$vȽ��(�*�C�ɕ6�^YꇏbK��QS��>0;TC�i��=�z��w��Z�Ba�M��y��A}"E0��U�	� �P�y����4����:��y&���yr�,o���"ᔰ9��-i����y�
��@���v$̃3� {햽�y�l���)d4��e9g�O��y�n�JN����@vDQ(��D��y�h�#)���R�}E^|P�I*�y⣏�~��w��de�}���� �yb�K�6VX��fK0�J��#m���y
� !����;��,rCn�-��"O搐
�K�0�U�F�F�A�u"O���%�P-!~,T�rBA�2$&�a�"O�����pK�x��Q!K�H`��"O��)�m�8>u@�*��- ~�5�%"Or��#�ܾ�hh�%) y�D��"OVl�@��
�k�g�Cl�"O�]���J4<��}hUg�K[xE�A"O$�2� �M����X�^��s"OܑX�J�`잩���^e,��"OI	0��b|4�0��1=,�+"O��q)Q.k�P�UC��x\��"O��b��D;E\�tBݘkh�h��"O����s�}���4Q��݊�"O����/>�Дjr�X'4��)R�"Od�̋Q:���a���#�"O a��Ɣ*�X�D�zȴbw"O��A͔���4�bi��Q
>yzu"O���V+8�ʽ�R��-��xӧ"O��bt��(O�%�a��"O�Ea�́$�����F�:{�bܢq"O"�r�3/�8W�ۋ���"ON�G���hP�5�W9��JF"O��Y�k��>N�bd ��1z'"O@���/K��(s�#V1�2�c�"O���C
�Q�3U��;�"x��"O���7-ɢ=��DS%f��ht��2"O���!h�Ҩ�I���78���D"OVL`�c�{$E� ����顀"O����	H8w�&����:d�T"OB�C$�	5X�Y@/�
��pu"OZi��oS)X��00N�1Br��#p"O$������y����%�\�dX���v"OҐ��HR�BF�r���
l<��R�"O Lxr�T%�leSǪ�08�16"O�@�#'��~��G�< 3"O@�ʔ%Z%f}�B�+I
h�qf"Op��u�BZ_��b�҂J��²"O�9+��6G�2�h7�I<�Q��"Ox���S0��w�8�T���"O��P˞�b�1�M��"�""O�ȓC�i�^���LK�;����"OĜ���<I�8`�t�_�t�p�"OvqW����<e�C�@�5n��"O���G�N�ER̭@牃nb5�0"O����Y*�����`�L�"O�3�%G� f�E��(c"O,52�ʛ�B��;ZJ���)	�R�!��
Qh� �6ÇI(q�Ո�>]E!�	�g-eb��<M��A����q�!�Y�@Rr�A'�+6%�uoB(�!���w�Xi��CS�\}���A�ǎ!򤇴Lb��G.?�a�-�>�!��G#$�����u<����m�X�!�dݍb��m8e� �\L��bK�z�!��DY��.쥩Gl���!�D���<��`��T^�b��P<}O!�ą02h\��8\�ua %M�!�$�m´%�A�4Q���
�!�[�>`||�gN�#>d�
>�!��:9�E�MY�p'��U�˴`]az�.�a�A���GL"@ �KU zQ1�ȓ28�aB��P?F����
Dk�l��\�Lj�g�9o �[���"[��܇�S�? 2$c�FA���@".׉o�����FX�<q�,R΁����@�`k':D�̑&e����M!As�H��y��C�I3R����_�.qf�
kc���d;扆 ��X0��&TZ0m�@]&U�ȓos�)i��	p�ȸ#�P�o �ȓ�ȸ��aM�=����-<
��5��r����%��`ʃAR2*Ĥ��o�~��Hp
T[�o�sT���Iڦi9o��<�&�[�yf3Yy�fY2�!D�0�ԩ�k>��(e��GZ��� �Qi �E��]"�
��AFO�P���k�'N��y��[�s����ܐI��r��H(�y��J����pز�XU�X&(�g�����"Od!Ӂ�K�8��rf̝k�����x��)�B*�j� �+=�� �쒧OC�I9��,�2��6���h��d/1D��v��0����a�?�4��!;ғ�?)��i��'�ֵ�S(E *��Ч兡G�!�DC�P���P�m��i��m��D�7!�Ē�O�F��e�?Z���ë�!���$7���[��M<��h(����W�!�$�X	�Ԋv�T<rX�PIR�J�!�$J��N�a%�<v`4J����!��A?*mjM� +ʧ�Ԍ��P:�!���UXb`C�M˃\l�I�E��cd!�ĞYv|\Ѧ �8a$���v!�T�+�ɒ���� �΀�7��>�!�K�ct��E[�4bE���_�!�d)6&4ȥ� ~�,e����4;�!��G�]�p�I��s��	ta^�!�$	(rqj��� s��\��ϙ$]�Q� D�TO_�%��Y�h	��\�rW�<�y��Z�)AZ�"F�ӨfҡW����D!�S�Ol-I�+��Bd�@�O�f�		�'��LX�B��L�^�B�:N�*�`K>a� "������5�,�{�% �.%�h��v���+���	�PD�$�C"^����p�L�Ѣ�C �Z|`w��w��㉓�(O ٸW�ފ =��AV��5P�E�V"OLq��#��ܸ�T�
�W��$��"O�
$�8�j�z�O[�2��xg"OzeY1D�5V �(�mK')�
�9#"O4u���&Z�6��u��&��٠�"O��)C*a� �z�k^�D���""O�q"jE�^���F�a,t"O�H�B+�*����6�A�YU�x�"Ob��&-F�75�1�6�I=F�XT"ODЫ��O�7'rE��,d�
�s"O@�,?58I��^ ��	��"O�@ó���Z�be`Б7��2�"OF!��HZp��Ҏ��ԡP�"O�iIt ��VX�)��"m^�؀#"O�I��Ϩs��jN�Z����""OP��+����m�5*2��u���	N���I�'e��� b@>.�6�C��
s�!�DūbT����ݽe���ꃇi�7M>�S��yRL+:��Ӑ�Y�|$̝ۣ�
��x�	:9�Ta%)H�.��dE\t�
�'� $	���<d<��L�9��C���cӊ�5͈��%����O���a�U~xCa"O\���
�|x䇂hv�\��IN>-��-��V4F��!i��Ϙ��ҫ0D���e'N0\"W.ͼ�Z�3#D�� ���V���t���*I�}�E"O~�{pfK�\3�y�G<#C�� �"O����Ɇ��u3Dŀ�s9��"O��{qfB�I뜽锦6EPl��"O\��b�:[������<Zk �3"On�ɤ%�5/pݢ4	x6��1�"OPlj�C��o��xP��&%�i�"O"M� ���.�P!�=R�� �"O�M{���~`�Ug��pn-9U"O�h���Y�.����C�\𽙧"O��hqI��T�p�H!��I��P�"O�����؍U�TQ�� �a*���r"O �vd�(HφԀ�@׸]m6}+#"O��h��ymr�9&��	���"O���3`��$i�兂�h� �h"Ov�kR�W̆�K���N�VUi�"O���#�*`46�k''���0y"O��ӧ���;Sf�|�Q6"O����ѐ~󺙈��I�_�8(��"O��b%��,C�@�6C��@ے"O�J���eip�krE���
@�"O����N�9���T�]�C��-X�"O�	���\?^�ÍW

�j��S"Of���֛H��4���S�gn�P"O�[�G5N�V]Q��7QVZP�<�B��[��!�h-C�4�&Wa�<�3Ñ4�xv`ͧ
�Ĉ���]�<�`�,󮩐J�NU01��X�<��Ώ�8�.$��C�	HR�*eJ�<��Ձ�
]Z��P+�xh:F�I�< ��n��haG=Z#r�r��j�<11�Zw_ ��R���+[tm���SN�<��Ǜ���H�6n�!U0|Q굮�I�<)	f��@i�$3��kU#
B�<V�ڎA�^����
H�n�A�i]@�<A	J��xf愖7U�y9��D}�<�P��
��9Q�eM5�����ZS�<�E-ғ9o\p�R�����HpG�f�<	�ş�l��X`ffB�O"��!��e�<�PE[=d�L�����&Q����g��`�<a�!LH��p����J` C(T�<�&��?%0n���D֣#�qۀ#@f�<a��I&̌ȉ��q�4�H�J�b�<��� I5���q�¿*�<`�@Q^�<�@) ����	@ȝ6KMq�JV�<���Rj���QI3�89�RDFP�<ѓ+H�E�¨���<��I��SM�<Q�B�b+��bA��'ml�p�c@�K�<��L�-G-R��#*,T">����`�<9 ��%w�t���	�Z��f@_�<�ef\ned�Ф\&<����ba�<�
��ނa���E���"�B`�<��n��d[������\��֥`�<�ŬE�Qx��ĂG�����Ap�<Q��V���� Do��,\�{2�Vm�<�v�\
MDQ���>pw��
�P�<��CmP�(�d�Ƴ<-���d�<!u��tqVc2�ϊ3�@,p��LG�<14��5 ��	�7�\�`v^a��C�<� gJJ��=0KA%Btu�vN�I�<T�F/"��@���k�n����E�<��!���I�Ӆ�4��E���f�<y���D3�X��!��Yl֜a!a�~�<ɆN��=��3��M�F��-ٲN`�<� f���1S��%���j-4|��"O��q��� �X�/ؕ�n��'"O�ShP�H4��qD�7�֔q�"O`���B�F�@}cQ��svN|%"O�X�񫒰(�ȼCe�P6o���"O��'|:< ��OZ�>`:!�q"O:LZQ�J0z�hM��dݔ$S����"O��"�U�_�؁��Ã?%dp8�"O�a���)gS܁HV�_�<��t��"Ol�
�#��#5r@��`�7&����2"OP,�k�������j|��Q"OP����*P1"��d��r�j"OʤS��Yz�|��'�	14��	"Ov�N98�z���R9I0��jV"O�Q��%u2JD3��2`��"O
H� �KV �C��S�3nd��"O�Eڣ��,7߆���l�5���"O����'u���%C�^>���'��/?�Uq�L.��<h�ɛ�R�(C��~�xMy֭ŋd�b�7+ې9RC�I���H��n�^f�XW�;;5�6M#��2���zj��!
;�r���O)lO���Pr$�#�LS����/GTL0�)D����T4(�rb!ӖF>��ū!D�pzp(Tp��$0r��,�$#�`!D�L�c�ޮ&љV�W졣�+D��Ifԥ�����
ZJ�y���#D��8'3wC��qE���]і�!D��[���/�~P	��G7;h���"%lO���M>qc�KG��Jg����2X��c�$�A��Bd�� �JɡVg��?!���~ʒNLbϒ��BE�.�B��B�^|����VBHL����C�rDXD��!����""d���o��i���G&S�Js'�E{��dD�=�c�׮x�fe��J��M��'D:qS��oנ���ڕ6F�	1�'ֲ ���.� �F#�BO�8ߓИ'࠽�,K�s��u)w��@����'U�����p�\%j�/  )K�m�
˓�(O�,0�G�t�d��7��(G��@Q�"O i e�(zF���A��n��0�"O>x@�A�g�,]��`U+_��G"O��莾*��uM�
yC�ep"Oޥq"@��5�Jt얎�P��3"OvE���;c5r�*ٌPfFqu"OZ�'�O�(H�:3i�y���	'"O �֌�`Q�M��wܺ��1�|"�'�]���מ3*~��NQr��5��'��`�Q�J:7��b��n��U)�'&�)�	��V�X���e�рǓ�HO.,�$��<g�@�!����1>Q� E{*�p�1I�nVpM���o�t(��>a�����K&ȅA���89���Oڑt�)D{���'���s���P�\����tP�Y��'y�At�YdS���`�<8@��c�'��t�D�	�K��9���/7X��'�,<�F��`hqc֬A�t�ș��'�,@�BI��9��AzJڠ;��1�'���ŏ%�H��H#Am�	��'�V5sr	[�)�Q�s���4�j�A�'a�a�!ͺ6�*h�� �<�<)�}��'���*��+W�I��.8��	�'��a�e�Ig.�6�+h���'@�$/y�h��S��3>�BH m�<� Fܢ��Odp<�J��r/,H�"O��x���J �u����4��"OV,��!@�:_�Mbq�̅8U�"O�uZ��K9r4�P��<(혌p���3LO�D�2m�z9jX���_�y���f"O�ɣn��)�chO?�9+r"O&m��dX�a^�1��%Xkb��r�8�M�H�	_y���
��37)N`����`J�Dz!��ڗo��A��dBCᚭ8��͛@`!򤚱uMY�1(B�S�1@�-B��Ա��
��Q�cƄ�#d+�.\�R@FxR�'�`Ԉ��#G0�A����@?�T[�g[H<�%/V�fOXu+��S4g���U+�d؞�=Q�A�20�pĐ-A2��Ң�&��x��6
�0�����a���)ӤL��0=)�B�Ǉ4�h(���Ga�����2V�t�=E���fe��Q%V)�52�n��V�5��I�X����ƫ��&�(�ᄣ�$I�JEH�/��Ą��7J��\��%	� Ȭ,��@�OV�=�}��# $�.l��c�T ���V�W@x���'�<9�X'=1� `a�A�nÈy�N��@p�)��%PDq�`��'n`I�"U)?���'铐0|�fʕ.1�tH�j)8R���q(�m�'�ax��Z6|0~Z�G�F��N���y�)�FY�i^�9�H�	�AN
�y���-S`�6�@�,]{C,�y�Ƃ�N�0�F]?zŞU�E�0�y��S�um(Ya1��o�4m#Ei��y��R������]�kXlp��Ę�yr"F�	V���;F��3Ģ�y��Y�n�)�/%6��u1Q%���y�i�sU��.X/0��␆���Px"�i�<��.[�R�9�B(�'�`"��+,O��a��� ��h閆�?�<\�"O��	rMK*������V�����'�^���b��p}�@@��
xDB�	��phq��Ԫ.��p�nY; �B�I�N �1���6��(�����JC�	)�0��F�\7��2l��<�B䉾,g��k�F�!x�A{���5!��B�	&�F�Bk2�!��D�Z:�C�I`�l-� $܎4>���EC?�.B䉫/�H�1a��	W���br�^6;��C�	.9:m+W���Dg��+%���.��'�@x��=`-H`E�������p9�C�	-:�LD{f'�+M>0��G�E�xz0Oj���@��=P���jl����	�z�a�ORe kޗk �1�eN�V@�:q"Oh��$O��`.*\
2b[/ڀ�v"OZY�g�b��̨��2��98��'X�	6D͌���60����*18���`��I 1�TQ)�@��8@ ��b��>�B�I=v��5KЧ��X�rAC�k�Z6�?�S��M%%̺�h�B�윊a T��`DF�<f:3!lUڤA�TLN}�
�E�<�1��(�4��PB>pE)p��D�<�EG-*4%� @�V��HI� L{��$���3i����Tn����؁��a�<�'�j?�1(�AF .Ѹ�����\�'b��'{�gy��@GZ���8m��� Abǈ�?1�"��4���$|�؃Cd�
hI ��1��'�ў�O�X���g�SU��G�PW�}�	�'T������L��AM�T�<Ii�'��'��)���d6K%J'LTY�ٲu�.�C!�5D�� Ið�
#lt-"��*1�vT�V���G{���¥��,� �=9�՘䭉$#؉'�ўb?Q0W�Ņ	~<Mj#���y�'I&�D:�O��Q�LĿ����F�^�7��)���-O���l��X��.�H��ܫ!�	�3��5 ch�  �$�p,��o�!�D�#}����#%^�j���P�!�$*z��U7Q�'$�02�R8c�!��"ZKҡ���d�3���E{B�=E��'�QM�4eR�����y�8�
�'���h0(ի.͚�s3f�J��(�'$�M�G�ߑ ���,&nm���'��@�ϖK�����a�0�*�'�ў"~�����x�v�U�y**P�a�<�L�5nݙc~>TēuBa��ε�0>�!��n*��� �D��2s�<�'ߕv:�$��\# �u+TF�<�ץ��X��c�[9�����@�<���.s�@���a�/p� JEoD�<YRe��o�}CA��S��!҄~�<�bđ�L�4�2�<q�dQ��v�<y�k�\�� ��L��0I���k�<!��n�����	?8]�}‍�h�<9�㎆x�D\q&!8^�@�1A�I�<�R�C���
�I�YY��[�<��g48�D[V�����@�&FO�<)umņE=&8���-J��X���A�<���ѫYQN���@dY$I:4 �H�<a4�
�|�CD⑎R�<)R!�E�<���ĪNr��@�g��5�й,�@�<�$�� /�6�S��E�]��	�pZ@�<�EU=k��H��D�2�P��c
IW�<�@C�7�J2�W�5�Qٔ�ST�<)�C%���u@ z�d��dc�P�<��3v���-|�D�Xq�<`M�=⪝��KҠz0��1Á	d�<A�����X9����U�L�"�v�<�A�-00D�YV\�3��x�<�l�"��qJ�E2K;0H�"mt�<1��׷������6h�s��X�<ABI��uD�e��e-#�J�z�<ك�]��04��ۻ(��i`bs�<ɵ�� M��M��o���P�q�\z�<�p-˶q-�@�C�Тp�d��|�<�v.����D
t�`ES����QP�i��_#�J@�6E˄$�&p��.'HŊ�H�+.��!c��μ	a�ȇȓ&]�b˟&%��ͺ��ٍt`j���'Ș�G-�9{/�i"�H"����ȓq�u��E��7��y�"o֧_�v��ȓ���P�@8D��]�C�P*.�깇�L�HH��)˃4p�˧�"Tn��a<�ͳ�	�P<��T$X�iC����Z�����ͣ-C�D�\�*���O���h:OZn���K9>�L�D�d�� ���Я
ʁ��!�4��E��M��Z��h�lHsb!��O�u;$�2��~�|���͌!�CV�`�QBI:YӴ��p����!�JB�q�3,ѫ;i6���j�K�!�$� ��Ah[!M��S
�|t!�d��j���BG�O`8N�!�J�oz!�䊮_xb%����O0�p)�!�$.��8�@܄=�ep�(��[!��}���b��@�@�І�בJ!�� �! T�0��e��H��Xh�S"O� ��%j�ꄢҦrƺ1�"O*q�dG�V��Y�YU�|�Y�"Oڌ����)��;Q��;�8�"Oh�@��K<p�V�M�b����"Of�"�֯Vw���*�[�"Om � �\����	p�.X��"O� ;��P��� �!gx\Q*O�K�i�\�,���f4T��'��(P#��-T_v���c�'c�h��'~4ś≓41�q�1)��A�f��
�'� �˥$��7k��0f��0bڱ	�'5�4: �7>���6*�3����'��� ��X�|œ�e�9����'���a���#O� ��.яk��x�	�'~=)�7�hrR+ė`b�	�'��t9�J
1$id�a�$�=b8��R�'q:m�t� %��M�#n�Z~Tx`�'�8�*��|�z�b0�6Qk�a��'X�m����00"z�����5el�Q�'c����	>h�̀*������s�'0��Zg�16��S�ʀ$7�j}��I�Υˁ	֭G����DԤz���ȓ��A��[�����I�%\hH��Nh�raL�-Jd���m�/_L���ȓ��H�b�V�-wP���+ �.!�ȓQ���@���Y	�8�q�T�4y���2�\pcw��p��*�
J����J �� ��2|S�A9��%�ȓ/�����k��C���R'&իfo����Nz*�#!R�?b �b��ڤW.Du�ȓ��I�0� t�~�
�  ?���ȓY���@狮A hqG��:��ȓ��q��Ȝz���ۣ�2-0l��~\t|���Ml�sgB��U6J���$�L��`��VY�3L��PtRm��F'\����p�k⩛"7�����ȱ���faC�Ι�v0D��� !Q�,��PF�:�F��"���hsd�c��>e#�<1�D��m�̆ȓ�̙��ĕ
 6=��U�oA�܆�W�0����pi����%U�D-��Q'j}�	ܳ%6v����G� ���`���m(�� ����}�0`��=�H��'��2�$U
5I��K2ҍ�ȓ�� �%	{Ɋ����B+
�@�ȓe����L)�^m�J޺+ۜd��;�x�uǇv|���V�%�ȓ ��<9#4|���` M�2ؐ�ȓ�ى˓;�L�)SK�4���ȓ �&��Wk��;|��i��<@���a�,�@�.-(���)эVw�`�ȓ���ɴ$� Al�����_�t��ȓ)$B@�PM|�ڥ��l�3(��*�#'�S��E��I���F|�ȓ�~�*��k��,��?3dm�ȓO'.zU�m�̚�5b@�4��l�<y�(�m��1i�4RWf��&��b�<IȜ�@��M��a�/�3�/�Z�<�����d�z	���0=X^A���W�<i�(V�#u����0 �0���	W�<�$�D�x� A��2|wr`�1&�[�<Y�� �%�:�D3�Q~!�]w�9�=E��bQ�u������L�\8(1��Oߖ�y
� .cc�Au�*�B����ʼآ�|�����Ȳ�'V����%K�:T+�Å	~eCM<�v���'�����h\	kkrIQ�
Vw��h��O@ Eʀȋֆ�E�d�`��/�O��a������p��P��Q�a�j�I�Q��y�a���6q�ϒ*1��A��N����%�4�Y�{8-I�h�!�d%���� �p�ek5�^�[�R ��.:. �:�(дP��]�����r���む.��OuX�Q͕�V�k���2�\5���4O�Р7��)#�<��L� F���Ds�q�vd�e�	�� f�0tGkM�H
6�5|��8�4�D��앓n7�D�B���y���B/?��e U���K$}���������n>���,Ѵq��pA͞{����cI�3O�Y#'����]�ߓlS:JQ��
Xb��Q�}�p�f�3}�ʣe���h�-K�G%޴�K��Ƽ"�OیF�����_j�4.��� ��Zy��	+n���U����x���gH1���3_IV�8�Ɉ!�ZQ FT�(=* �U$ԉ����!��d��Xfl�6u�ɠ!@8N�Q�Q6�H�f΂D����S]vI��/dR��3�*[���]��!V�px�����?'��AʠH�~��7�ɲ
�8��d���*�~!�Ժ.���L�E�2-׳_�L��r]�P�G�J�?�nK�x�&���dϪDD��
�Ȁ%rD�Eƙ`L�Zd�.}�H��'�Le(F�͇h�0L
6aT�Z��H�괟@o$fZ5��%v�Dq Mh�8TB���Y��`�w޼ B����}_"�cEҖ��\
	�Wl ��&���/�*�ɂ��!v:�8q逈l�`$�p��d�c��;T����ķb7hyg�V��'ގ�X��OЬ��$�����HI�[i ��Dڴ5(���C���$ k�̠R�n�d����Z  ���$����w�V��M�[���CK$9V��}[��%�#(4�ʓT�Q!Sh!6����.!�IM+�Ja��fE^�81�"O���A��[�(��	+
�
�ڥP�Ԋi�:+HXexHWnyZw�b��BĔu��I�O���Iޖ-�^�+�X+
�������a�F�5@ҡ��鑆Mz(5�&�!ЊTK)O2��t��3
�T;��$�=y��!��	 �4���+E�~Q��c��ڜ@[T��'�<�G`Τì��p���k���p���Ck�d�PLz���8	O�"r>�ѧA�:�稪>���]�?��'���R��xɧu�=l[pT� �|��E �yb �PN<�	�T�~Ω�fƓ5���Q��-��:��}^��%)@�uإj���dB���2�F �p0Ш3�O�4#b��#�\5"�x"�Y�W��!�a�/\���M5�y����k28A燯
��|�����y"EZ\���Ԯ��S��	�+��y�
�1.�g��fk���	�y� �7��HJ�N�+���j)���M��fH���sM>E��4,+4\�ѯ�L���	D*7�͇�]�L���&�*��I��E�9�����7c^}0��b-���d�%A5xm��Fo�p��֡8]�a|�����"G#ҡ��Hh��ؖK�"�£Ƀ,u�E�O�Q���g�E� ��h1����I�a̸�r	X�4�ӡ<w�x�T��5T����CT�<��ʺd*bAM������\��ہ&C"��$�(O?�ɩ���Q�E
O�YP�I#��B䉃WidXIfY�=�B�ץ_���	Ff�e����~Z@���I�'j�eH�E |x�'.�4�C3&� �#�~���,P�Y(QD �Y(B0�c�N�D�&9��%�FS����'���كi��~�����`G�EI��OeQ'I�������;q$Mᑏ�<YR �?eׯ�E�dM�ԃӘ'3� �&'�Od�Q�	M�n��9���_�����U�n������r����Y_V��)O�mcP�7�s�����;p�����M6������"ʓ�*�8�'��r�����-���ħ^�H�G ^�`u��L�~��������coH�b����ǯwRqO��1(�~9 �dP��NL��.��/����j��bK
Yr+D������S�'vc�u����T�j�E�]?)��<�1ebZT햰Y!��Қ|B���D�w�Ƚ��ׄ*2�Ʉ�JM4�`���J�`m袃Y�O]��3�7Z��k�E�r���"��U)tg
dl�9xHּp �>Z�ў�K�
�;0 ���.�p�0h"Ԯ�[�P�{1��)���8W���C�џ�c%�D�g� ���'�T=y6J_|o�D��J�d4�9���C&2ad�2RU<���d�A�Y���k֒1Sr,�>�ਸ�ۈ7G�b�p�F�̒'�Ec��S&;�U��H.C��B��p͌�@�#Z'/ژ�R�)P���Y!��(ڧ�y��K�{��`W�ѯK�@x!�\����7�_�t7�&�>�S�? h�!���5Q��X�ɓ1�p[P'֟#Ix!qc��@��qC���r����  ����0~&.(���_�B�6-\�g=l�qf/��HO&,��*_�G︐��.CJ�X��1�_1�>�2�ڭc��I�$i� �#?y�AG�,�z=�e�O�@y��@26(�|8SeG+�ܙ��D[;Q[<I�B��caHl��F��T/��'} ����*(̪(	"H����>-*U�v��	o���}�� �/��u��gB	І5y�$ֱO��(��9r>��m�eNdG�d<O� *��]�b����'��	��Y9ī# ��58��|���鴢��
�*�/�.)R�O)�鱁kP�V����a�� A'&��?�QNa� �\��L�
@�� �����%�P�İ�PETZE���(�e6�!)׈�[�Ɓ�n�i���`��Ol�y��:�sӰ���P&Y���p��>p�F��ቈT�t)#)O�H���ɱ #|��'���c
�+��q K�1�&L�Q��p���[���߷�%�յX�бath��q�D8��ϛ��TE����E�	;�k�O�O�+��D�9��QJ���I.�=�&,6�>zd�ڼo9���CeP1�e�^�z� H�gՇ+����I�X�ł'jA&}X}��L��FoD��<q����KE�̇a{�U���*M+
<� �GiX�p�!��P���� �-PE��YňW	| ���8R�r�Z��X�S�l��'R��e+Q��<�s�0$PIFÞ�&��yYB��m�'|j�`F�+�l��}JqbBŞ��F�'&Y��I��<1�`-�"д��<��E�)[���Co[>'���9�%`}��ݜz��=�=�OLFa9��J?F>��� ��:j�t���_�BT� �҇TB@��J�8� u3ӢٷN�ڂ�ي[`�0{��+{�)�&�s�'T.&%#��ruh��p��Y��T`|-���T&p�n�!�&�&V}zyI%fW�~�By:GN�����s��kS��T�*x��F�}����N3D��� ��s�8�@��D{��+%����F&"���'�E1�'(�-�@kN�S�D���
�z�0�A�#h#b��IщG��xr �9����E"O��c�&E9���3l��)w��"O�006a98�(xy0�-/uD]�g"O~��s� RlX�Je
^�3a�lR�"O���AT{�����ǈxuZ�{"OT��M�#\v�A��W&%��q"O8A���ϰql]2t�C�2(t"O�(sdbb�zPC��
���Ub�"OVt�Ve���]�̜��X݋P"O*[v��&��؛׫Y0V�j5 U"OT�@���K/X��UO�"2����4"OhhpbO�K�HkC�0̴���"OLIw�؃\�:h���g��� "OL�"�]�x���&	�b��l)p"O�q���T@l��� v-, �P"O"dh�>F=fi�ǂʓc@�0"O��B��8H�H;��@�W��#"OJQ���:�8�I�p���
R"O,����A�20飑H�RQ���V"O0�U?G`�3��E&TLc"O⽂�I@s^��#�ʳ9:L�"O@4)1M�
.�>iQB��1,l�8� "O`�҅ A!V��@
�@ǿ,H2�a"O�$���ݗ�� Z�W;6�p�"O9C�&B-zV���1/�n.���"O�A��vdP;V@T���!4� D�Pr�,<����eM�
4�Z�8!�d� ��b\&:8�	��d�!��4D2ei f\�G�twd��0J!�ę#��i�@V�~�m�v$@�9!�dѾt��=C�
��*�(9��c�&(*!��,� �x0!�O��D��#��!���V�R����N�%v�$ڗ��Am!�DP.=ߔ��t@@�v�r\z��؜8�!�D�1%H@
 O��Y�ъ��!���
�Q��ļNDٰ�Ĝ/!��%��3�b #T"�i��G�v>!�� ��5�	(�2�h�8��Ƞ�"OL-{��ź-8������A��Y	 "O<��ă8u*X@��ɏN�V4Q"O�A�D�J!]�V9{	5Q� �c0"O�19�IW�}��� ��A�^�0f"O�	e��?�.���'L�Z�0�G"O��6�ɶmh(RK�3B�2u D"OV4�(�8Q���-in�9��"OFP3�K���*��rjG�l:x�y�"O��ʥ"�u�,��֧�Y�R���"O���$
0i�¥���b��4�c"O��AФ��8$h9�U��p"]�0"O�(��i�
F��t���B"Oht�ʔ�*�b��f�;p,eQB"Ol�kE*�	:��Ѧ_ ��؂"O��"�ײq�� q�Q��l�#"O�ݩ���n��H�'�T}�B"OƼ��EP�X���;7�Ϗ�*H	�"O��@�+�=4q��
�2=�"O �x�`+F��p�$ϋ�2�X<8D"Ox����lЂpas(�#|r�� "O~(A!!-�|@��G5�R!"Oq�R#��|J�A!�o�4��Y��"O�Y�Ŋ��j�R����/(��ݛ&"O� )�V��pX�f�gJ�D�F"O�P��o��y�)�R��a,��5"O
�a.o�r� 4.A�.����"O�Ձ�n_�q�E�'c�*m�2"O4�A-�5�\xC�	ې+F]s"O��ą��)�d�*Uȉ!Pf���"On)�sc���D8�G�L����"ON(�5�ӡۄ]��F�&|	[�"O���1�Ԍ+|k�DY�u rL"F"O����O
;��D�H+�LbR"Ohp�[�R�(����y��\y"O4�bףA���;2FI�j���!"OD4 ���2Ub�G&�4G�Q�"O��Y$�ҫz�|h��F¾0���"O��tӽg��9cD��c�8�"O��@W�T�X���ő+�A �"O|dS��\3�L��w�>�T�t"O�P �(I�`����X��`��"O�8��Ǘ�z�8,���;��1�"O6��7;.�x�B!�KXD8�P"O�0��8�l�"� ]���LR"O��R#�E�C.N�{ �Q<��s"O�9�����C�:���u�-�V"O"4�C�N<+{<@�%]p&i��"O�X��g̽`&h	�\R���"O��Iր�<�-��C&rT�-@3"OP,�f��*�*�!�B�vDPz4"O�ȃgPjW��se"G�`vY�"OtA���T��p"�+D`ˈ���"O�]��c��Kɰ��AӅhZ\H
P"O�(#Ed�.j�N�hd�Bh���Z�"O�!uH���p�ӵ. N����"OĤ�UH�#~d􉂖mG�(Zn9��"O>Eb���6��Dʑ>g��"O贱@�؁4��B$h�kQ��"O@@�$�� ���wa��P��K�"O4Hr�n�8[���#N�N((0��"Oȩ�Iޘ|�X�Hp�U�f��-!�"ON��%�͹nP�%i l�@�� �"O���a3 ��ѩ�ʼUF8���"O� ���a W�5�M�ׯ�	J�a0"O�a�%��?D��31�#@�ޙ1T"O|�;��θS�8	؆ �+3�+p��t�M�,WqO>�V1�Nͳ'��{3,A��:D�PCѪԠ^��$� Ǖ�q?P�i�:���s:Z�I¨:OD$�!�[6'5�� �b~M��x�A�%���=�O���bv��2�r��/D�0hȈPT�ɬU*��p�0X�F����H8���#�ADD������B������C���B�����gC9">hQ�X\�pm�\|6�]�
̺�h��yD��A`�.�C�	��qL�Ĩ��aA(5�e)tL-��Ѱ��L+L�S��A���Q�����C,5:|����h=A��+O�`��Ⴗ!��]��>9c�U`�|@�Rk�?A�81��.��0NJ�PI$/���C�
Ҡ�,�O<(q�?��kΐW`*�Qq��f̈�Y�Q~�B�>#��!è�x�T?s�H;$�d�y�/�!J2�;� �&�F�Y���f ��`�&uJQ�'�&�Bc�K�#T���Q'��	A��Rn��K#D��cr�]�[g4Q�ċ#T����$'����% ����"�74L��7�Aya2hϡI.`���H�Nbr�
�-G�F' d`0��$�ĦƩ�|[$��/�`�qA	L`� <���,~"FmRĚ�J��-�� Y�'�J��w��$0J����M?��+�N>H�A��K��j�ʽ��0�DC�%0P`���,d��Ի�� ���Rj��/GH@�0lܡ@EV�+�
͐�yb�D�	��:$�E�Q���'�.g�O�N�rC��B���7K�8���b����� {���C���)���	6Ξ[` 	�\ҭ�"��!)�J)i�'I����.��B�4˔ {@ ��Z����!�)�@��V|,D3��b��jE#��0����	�P 6���a��n�̳ťӦf�����k-�����A<Z^>ej���.�Jq��O o��s?!��:�!&��,�T�Q�0D�E�4h���8c֊B>� �P�H�VB�:X���Ӆ�8F�U��ǢI�~�І/Λ?_�� Y6�m�t���}I�'��y���LK XWy�mE#@>-9��A�p�D���d�e�\�y4�Z$>C�ɀo���$�2{�z���'�&,�ყ��,^��8()O�.�<~5t�����<Q�Ӽ8,�aB��ˉzQ�4ç	TW����TjK��r���Fj��"���|��!ǣ�!F��	�恂����џ�JV�X���!urE!%�!�l�aΈ��dZKV��d�ٕ(�xI������	�ZJ��M9	����j���]���C �1��T�'N�����\B��-4X�p�Em/������dh>x�W��"\Va��"O.@ZBȕA�aq���HѰ��[�\
�e�
N&A'��|rԪ�=�!cH{<��4f�|�<Q6�^ ���"�
\���y̓��T��+&OF-��J/q�L���p>�H�"OVH�g�,�̔s�ʉ�C5��"OȀk��E?A�B��(R<kd��@"O�]hB��v�	�H��ID�q�"O4�Pg�t�D�&]�p�"�i눴 ��4ɧ������;(��"��3�zcëT3�yi�^! aߘ ���Ҩ���~�J�A����._U��TQ�o��L B�H-��$�t�8�Oh��dƉ'x�����)B3w|ܥ	�i��>;*y�+�<S B�	L�p��F�=��Bc��P5�"<)@j� ���2�\���O���#r��x#Dp��Q�Y��а�'��bĉ�ME.m�V���P�R�*��.,J�����'lG�)��<Y��H+]@�dcc��o� ��Ya�<��M�1	��#�mx�yB
��<	����L?�]�&��6��<��L�2�ܨɔ���c?��P�L�ӱ̅1Fh��2��Y`^�Ua��D�<2&=�����-�Ɠ7RZ%ao�<R����v!�4{ ~�GxB�Dse��b*_{��8}rF�A	>��ɀg�K��)�v"O�9z�KJ� �������֜zW�#U���2�������S��ybgΩk�9�¡�2�Jp��j��y��Y#����0�89fKN��~"��zɊ���ሱ[p�]��!�)��-��5��H3���t�@�ЭL�����Z�*p����`h(Q��
_�L[�iQ�`����&Ґ���$��F��'7�x��bӏP�	��$��m,�	�'�!��eg���a�س����۴d��4�L�#��dM#�^���H~L��a�ًUa{�B�x5�;!Jڟ� 򑓆#%q�I�c�G��Qt"OL,8ҭX�,��Jã�-z��h�#��^�*��8R ��h�f���,��DA�+W�X��A2�"O���.�>���!��R�4�"���,�������+}R�9�g}r�H,xL����Z(m��3����y�%�w�����m�sn�dE��Mk�n���E�!�-|O=;��*\��Y#b/�B�C�'Fd8�A��*d�0��"A��Ӂȟ�"dykѨ��B��*Vg�|�G��~��5�ͱ;�b�Hc#,2�T�I��.BZ !c\�J0��,g��C��N�ę��R�\�;o�,v���
�{|�O��}�tZq���Z�&0��V,�/��U�ȓ;���%�*q�����m_q�hΓ(\����?�OE;�O҅m Qx� ��;B��a�i&�A���� �ɧ���VB�>/i�k����|�����ߟ�y�R<҈h�u�ɚh�B��񦍵�~R�.AK�P�Tb�O���G/�g����R�Y?s�Vx��l.�O��{�"��dt����&���I��MB����<W�C�I"5�cC�]�L��h k�6%�"<��`�N~�SFF����Oe 8HeJ�Q؄+�AL<R�� �	�'�6,���h�.�tnʧ"�� �D�=�`궨C��)��<�q�N�r�J9;���y�����~!�$��3pR<3��.i+��x�/�C)�d��P���F������d�u��2��;��[ҏ 8,a|�{��q%@;a_N��疍x,T�� gX�i��`�O�E���x戵HTA�
�f����I6"�ۄG�'���uB�2=`I�d�L'x����`�<�����-�!��%GV4�Ʃމz[��I��d�Tz,O?�I�W؞�	`f�~yq����c3dB�����6W_4���� dR���@�H�1V�az2JR7U�ȹ�CO��>�	�C���>4O�:,BA�jĂ\�,��p�^54v��X�n�!�d�&)��r#1W
�M�1�>p�!�d�� �h�Tʟ�(儨�5��#�!�D��z�<	�%�-�@D�"��[�!�D�z���Tl�6Dͬ A��H+B!�IR!�PB4�����h
R��'a�!�ΡnN�u�A#މF&�4hI�!�d��S�h��l��@(�"؊e�!�d�}�"�9���h�J�4��t�!�դ�4�J�J_�`M�
��ʚ9�!�d�1b�d��''�t�ӾZ�!�$ۭJ}vaP�-
δ@�c��!�$	�i��Ԓ/��n�`�U(b�!��;A�6�k�U51\���"[l�!�۩�����JQ�>9���t�Z'�!��
)e{v����F�v�P��ƉS�v!�d<p��f@9]�ޑ�
֮yR!�Q&��
%�&s��(�'��!��7��Ѡ+���Y���:n~!�#btjm��ڀ_T"�b@	�08!�$D�{��$@��Y�l9���m�y$!��Rɸq�牞�>ʉ��fY	5!�$�	ua*|�pP+
�('�!�䋍]���ʟ�Z%^A�kB6�!�D�`�H�B'��&+���jJ
P�!���V�<�持x��P�'H�1�!�D��xي��⯁.W:`��@��!�
]"�I��O={x��#F̓�!�DN*tҜ���$2r���S�àX�!�$�!ú]q��d��)�S%�3!�$J�CR$�Ұ OR��K���G����<�g�Ԭ$��yс�K'Vh]�?�u�J*AٺE`̓a���Z�Kr�<�#!�T���Y���R�*�g(�b�<� �t3V��ނu Q"<��5�"OD[&M�e�pJ��D:H~$��"O�Z���lx�p��R<�P�"O�`i1C�))K�K$DNQcD"O�H���Z\�~Q)b�@)b��b�'?�����nF&�s+U�+a�����Q���'v��?]لLPQfV�.S��i�-�4��)�L�CTk��*.|L�s�΃KWVј�MD<F��H�'pa�.ܑS�e�a��q����$D�a���hP��$#�p��S4X5�Q�!�h>�� �!<C��U��[}"M9��	���O�b x��&2�zYr���L�(�q\��A�K��V��u:A�r���Ӵ��X���+~��.Pw�bMۑ�N�7��a�2�
5�S�O���Ƀ�x&��F�
����!�`�3�4����B�k@�p�`�Z
>���Oh(8��g��Zy*��� R�P����H{��է�<<�� `E$���/��j(�S��\���y�/Q�	����B$�*�l�"|��\�@�؟���L˹x�j��oK�y@��i��O����/F���ԹG�Z��~����$�����(WD`���I�^������5��R�ʟ�U�Oh����
&'�b�`�K�F�Ё��Ɲ]ԦpRr�v� J$��̸OF�O��dc�H�>,R�W�&8YtP�d-O7�~Ҋ@�h$<����|b���\0_��@g��k��-	�fa���r��}��Nޓ2j�1_?�G�Di���$����޽n�N���C7�?���)��ˆi��x=��)�aip����;�6�HDOH�NC9ֆ��<O��� �x�����De�<3���s@�� @���NN��yBiēfg�a�B�.dJ��5,��y�A��L���j��U8z�p����y�	�Y먘����(�H"�@Ȇ�y�Ƌ0]�D�I3�	�V8�e�7�y����!1  
N	`�����yr2g�r���_=i"��b㍹�y�%M�\��G�bZ��2!L�yGC^Rf�ҡdK�Fv�)R��;�y��E����2�a�I�@�XA#N+�y2��5*�x���2*wR��g��yr��Ԡs��� CGʇ��yr�X'�f� �gƉ�� ���
�y�OX3F���t"�x!�](a�yҡ�/eB���C�*p�\0i�2�y�痵=�D3Q��`��9��i0�y�/Ll�sv�⊕�rQ-�y���V7�p�� v�
G&���yR+
J��ŉ�g\���HË���yҏ��4�t�R+S��%غ�y�I�u�)��Ǜ*p=�y��@��y�1x���{t�&Uc���ӆ�y��_R�\,���ֻL����Q`��yb�b���BeFQ�<��p�uC�y"�J��Y���6:B���[3�y"n^�$�̕`"��B��$��y�kP�����H�$�c�'k��'H�����4�<eYuLI23�5�
�'��[p�PG�X��1�H.κ��'܊����ؑ�k�*�Z��
�'La��^�1�Y���!7��8
�'4�0xe��C( ��(ە4@�	�'�N_I@SO�O�,isd��.~!�K�W��BL�u�`�$c\�!򤐁J7�U� �Y�Lјq0��؛9s!�;we	*bg̔Un�ؑ i!��s&a��n�zER�N� a"O 0�OI=v(��c	���e*�"O0��p U�P� �z����A����"OL!�,� mxF�Z�Q���5"Oh���Mn7�@j�Җ+�HpQ"Or�t(�Y��ܾK�&���"O~�20퇜/h@����\z��[�"O� 2�Ç���Xc A-[�<���8F"OVA�-P#>4I������
�"O6�Flކ1c~L�Ջ��Də�"O4�K�/�w1�<��I(�<|�"O��QwD�"��$*�� 8|���"Oġ�A�r�`Ѱd�ѐO,��D"Oj�w��q
x���a4f�Q"O�ɡU�I1�@A�A�T|$��"Ol0�^%=	@�8�jS�FX�x��"OD��aƃ������~n,5��"OTu�ե�=�4(KVC	.a����"Oĩ���B�YC�����,6;��"ObAy�QD8H%c�O�� 3"OJ�h�)�#��CU(j�\ͳ3"Ol�Y�v��L�ԡ�+[�DX�"O\��֩�>-�d�C��I+U޴$��"O
�Rb �V�ִ�!�A���B!�$���N�[��Ȧ@a��%O-Y�!�$5[1�z��lm2�B���!��*.TT�*2��
.o� �aA�_�!�D�`�^�bn�7]f�� ��?�!�� A��:�b��)�A�s�),!�X�w�p`+VO� ���B�|�!�$E�-�r)Sςn�,��l�.A!�$����<A#�˪�F|CA(A�A!�{$��$N��k���0g!�C�8tz=)�oZ���
V!�r�!�dKD�����4#��|�mƓ=!�D#��Y�K��Ji���^�!��ȹw�Z�q0��CU���̓$�!��i���#E^�R�� &�_T!�d_�.#���S�H�D�)R
�#["!��@Z�2m��i�5 z���i	83!򄍋^�Z��ɣCҮɀ��^�AQ!��x(X\�c +8_.	b����!�D�J�9��Uu�|�&D([�!�]R ͐UΚ�~p��[��P�i�!��`Q�T"�菡YATx�UXP!��A�X��rL�>��Q@�X8�!���I���p���0ӎ!��'��U�!��M����*V�s^(���ʧk�!�ȶS�Z'��,�(\˰&��5�!�XU��H�kp��C��3t�!�$,\[�Ď�'D�)�U�h�!�D�7y\����3O>b ᴀY�M�!�×Y�̨"�O��+x�07j�h�!�dR�L|��Û""&5�Ǩ�+b�!�DȘh�^T[��Ƞ:-�@�Ж �!�ĕ/M F�#q�]�t*��2D� (j<!�D�	��uI�L��s��1;!!�D�@y���"b��ءƢĖ%!��ܰ6&��bͳ�F��s��"�!�׭3�r)�mȮ6�tE!��8l�!��T�x����l�2�
A.D�Zk!�$�m�`�ZC�R�]� ��Պ�/S-!�$�2Y7�(')����3�JƇ],!�Dԧ%��V�X�S��m[eI��\)!��3QPHYx��x�@T�鋦2!�$��H�E�"cX/v�k�&��!�dع��]A#.R�`u\-��;`U!�$G�S��B�H��Ab�--4�!���*~FdCӏ����Xs�L6(�!�Dȳ7��Y�[J�h!b��}�!�+�B���?:��\���H�{�!�� Hy�t����f�hT� ����A"O��SȂ)'�\�'.Q�6�0"O��PU�N�g���.C8y�J݉e"O���g"S�x�A��Z���U�t"O��@��5���Z%�2Z���W"OtPj�_�^(���J�w<��"O�z��9�����&ρ.	B��"O\���OAqIƸP�H+bKNx�"O�h#�/\<z(u�@� L�]#�"Olf�/�.I�1�1L��	w"O����"	'Z64% �Y�L.l%k3"On�  ��W,�RF�w��Z�"O�@��K�>o	��(+6�	y�"O�FAS1e�]CĉNf����a"O*�����d�z���/d��"O$x�F�H�{]���C�Ҹx�@8!"O��r�ǅ!U����BC�/m�Đ�"O`,�jנ���g��	�rP�"O"����P WnL�P�Ղ1j����"O�d#�jϷTb����ST����"OD12"�E�~��	���(ZM��y�"Opy�GF��$2E�W�l�����"O��2��t+�����@5���T"O�ԃA$��h�t�{��)'��U�"O��1��:/�|82�@�J�pY��"O�Xs5H#
�8)`�՚���"On���J#:�h�e�H�d��p�G"Ox�*��N�f�u#/�֭�7"O���4ƙ:.<�w�-_���"O��c��K!p���+ժ5j��B�"O�X0&E�(�.P �
�\Z�Hf"Oj���,�I�lJUi�MQX!�"O,���K��&�\(�梅6_1���R"O̰��)�O�|1�k�#^����"O�����*�ly"��i���"O�"狕�襀T��cK��y党-�4 
�)�M$-0ã���y�%֜z���5`�?1�E��cU��y�Mٽ&Z��V�ؘ@Zl��2�$�yb-^�Pux�2QG��<���CC���yr���H���Ř-� H��ג�y�)7�rXi1)�.` q�qFR��y�(l۶��� ��&�`����y�͌9!�E#B+�V	��L�y�n��KTt�R��3�4rԨ2�y2Ş�1k ��wSNB4�����y�����`�&���@��LW��yRE؈nپ rǆy�Ll�Iԙ�y�fMU-��{�0Z�4�����yb�,Vp*6'��J�����׎�y��&Y�R��<�����љ�y��&�p�@��' c�;�̑��y�.��M77A@�&ն1�G�U��yR�.k����T%5�͡�P#�y�-��K�a� ���j���y�+ˣYx s4�W��ƱqB��'�y�%���~ͪ����Z�	�����y�F�. .Υ�b��NZ̘	B���y�ɕK�4�0��9T@\�a�'@�y2�ɀ����Ǒ@떔�7���y�"��-��lr����-�,�
�!μ�y"#?i�
.�;B�`��y�ҭ,l��[��<�B��4ϙ+�yb���hU*cT  i|͡t�^�y
� $=�D�14|����(P�*X��"O �p�,t��d�Q�-p�|�"O�16̏[Ry!BmWlc�]�b"O:�Ic�Y	l� ���_�I(�C�"O����+	�/@3�I|���%��y�ɂ�?�>�J3�^��n� �M3�y�Oz��K�]��n�*�`��y2Cդ-]�0ca �x��[O(�y�-]�X�@�i��j��\�/�.�y�$�<T'(]H��
�G$�y�}Xx���(<Z��=j��͇�y�O# {֌��kS-RD�R3,���yR�κ̢(C$�Dxz'��m�\��70� 0Ƒ�`� -b�$�T�$\��E��D!�G[-����h�y	.�ȓ/Ģ��E�L0*����iǊw�:P��{�D:���+m���e��?�ڸ��EJ�ٱp�G@�@��K[��i��>V��V��V�8)�Á�N��Y�ʓj@ܲ&�.n�8��g�ӞM�C�7(�lyJ"kX�1�&�R	���B�-V�(�;��[�H��h�J�Q��C�I�OZ�	�@;V������K��C�I�B�n���Cʟb�������BT�B�	�I��IP���"�Z�I��
T6C�!fG�iA���m���g�5^*C��=���$�T/q|�c1dS0k�b���	�/"�@��i��>EK2��Ge1B�h�HL�(#��8�Iڟ `p$�0*+��?IH|juaΘ1�`���-Z�,PuA�m�"y��#��	82��&Ǻɫ�fX�����('˜�Z�cF�NH�P����'������?16�i2���.�6@I����U�\�P�뇃��A�ʓ���O>˓w
@+U�7]Hлr��`���<�ݴ:����'�@�W�J9�dءÓd�v(��oߵ~��m/aӚ�ķ<�+�����O4��l��}8�LB�dN���M�:BI2 �ɐ^���$���|���3�Pu�4�ƶ�������G�Z� �	^�	%�H��ɿ!Ā�F�ݖ�r��DI�-T�������?��Oޅ�'��O�L"(� ��F���q��C-2����/� ,Ox��И`)V%1fo�;��M���$���	L�'�?!ش�\�S��9	�R�d� / 	�=��`�i�i7��'��|�O���C�TA�`9�J/s������2<��Hf"D��0?yէ5S��L�ed�Kް9��� c�u*��I�=���4MLͭ���%s���9` ��0G[�y����q��fv�Г����8�M����O���M����(c��)�U~�l��A��R�<�ҥ�xLƱx᭏5e���±Ǔ*���'6�6mr��nן��O!ر��uӶ6��4?�ЋK+.Ā�Q��M8�����&����P
�@�Ɏh���s4jC�}� ٖ�=>f~���Q�[��e�7.��%��#9cB�Y�G��/L������m؞$b�E�Ol�d|�ndQ@8f@t�����P:�ܢV�>���?ٍ�O���8V?`��Q1+}zѩ6/�/>�C�4y�z}Z��� Y*�O��
 Ik��i�Q�p�����M+���Ov|����G�C�fY���Y�~ʬ\P�'?"�'ޔp�5�|2�'߉Oh�\�&@J!=��Px��s�����}��P�&9R���2D��DUD���B��I��A_w�uа!��ҟxN|��Ou( 	s��8D�Z�a�G�%n�&��@�Q��?E�,OJ��І�| �ݛd
�������'P7�Ȧ��'��iӤ�
Ե��mOd2D˒CM,�nZ������i�OX���O�7mJ21	(�K$f]�Fr�q�耎uF�&����Tfq��'Z �C�u�ddРm )1�~��v	�^�4R�h�^y��7�g}2�T c�ܔɳ�	�>���P�`���O8��'gD*�����;��3L'�)��M�Kܤ��t*��#����J�'ˀ�Y�ꕿ;��]�!��ko^��{"*b��l�p�'��ߴ,��xـ�ԗ}T�h�!�.�RD�O�����!6 (  �