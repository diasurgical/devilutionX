MPQ    �    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h�F����|I�,N���
��8J߬�Q��᧕� ?R�vl�+�ꗍKJ8J������8m������K��f�Q��y#^�]�&�ġս4%�~������&�1y�����3_��	v>�(��i�$E�8��R��y��������������9��|u��5H
�W�����L�=���hU�>Z�<� Cݥ~<1�q���M�{K�>Ƨ@�v�K��m��z͎y��*��ݟL�lb�jI���Dn�Es���䓓���Dᠨ��xa�>zJ�-��E�����4tV`��ǼJ�#]:q��N��i��7.䮐/fER��٣ڵ)B&D'��B�@�Zv���I��V��kE ����x���P~�RR{(4��э���P�.��&/����'�ѿ�W.݃&���d^�����/>�:�q�����(�H�K2���t�U[g��C�����VxPt�(���*�ð��D�y�^��������`�~l�Ng�/Ft����<�k3��>��ɼIO+eU���ȫ����
D:oL.�?P�uj߫J(f�) Й��뵱y0Q�6`v<���vGv��p8E������f���ۥB�l)����!��=�(�̥P��rⶉ�$Ml9��;���B��� `tv�Z�YF�|B)+�|8W;��Q�Ns��`?�`| ߍ+�����Db���d=�����r��Ϩ�xlL�1U�"��i���DL%��aV��A|Ų1��eO��Y��@`ǎ�=&�����[����{6�;���E/��q���Q�ѻ���Re|w��z {풴4�� w7�`��x�^�S��k�����U�=* Fَ(��0C�f�T��xK^�Rf�3�9����^nv�����C	v$m�������Tl��R�� j?�u��s����j{4Q�ʊ�Ј}=j`�F�b���u���9C�)|�>����X���7s�g5�c6���ti�g�<��N�'��"�Ε-,iX�*(�Bҏv��5�wL��S�E���`�r�8(�:�����>���*�������3p.P��^�?}^��6�L����&2YpBJu���n/����m;�\�T)O��(+��>z;8�H�����(��Za`�p3PS�:G�=�aH�������JE�6��$���|�Nm�ِ1g�Mj���z���o�T�[!4�h�'��h�qR_�v�W��魙��I���@9��WHD0�f/�^�u� *�œU�V�$Z#���s�ZDrT_)��	f*i%D������	eʺ�@�	��vL�s�!*��F�8��V�L���Xu�0Gq$ ]�����6�����^�k>XǄ$W�� �&�,�AA��'��l"�%���� ����9�mV���ϰ�?ԟ�W�s��N����	��I�M���y�
�}kNvֆ�J���E�!C��0��ADnG����<lI0.�#�m�{����dѯ�b�UNz(bS��R9��8�CG�{��˛pH�Or,�%����Ц aN��^%���J�/yw\J�F��D�� b�Ɍ�^��k�����<���:_\fR�Al�+n��c7v��EFpڮ�H���J0	� 85�]_Ө�S$&fz8�� ����?�O��@%�@\biݴR��6c��i�:B����3<|/n�*��ul5�_���;3�a�SH,�R Z��"Xy�C��q�x@��4���Q����X+�v�})#'T|��T48�_����Aآ�]� ��oI�#��5Dc:k7���7��b�؊ ��o��
���٭n��Ia��XQ�v���nuff0�ଣj�����"�u��d|&>�¡|��5g�ĴP�����cɻ�����W�B�J:gf�����Ћ�ҿr����R!�j�0���y�zFT���{_��kz��������<+�~:�=�O9��A����F�]�ֽ�省�V�(��(�QШ0:��+.]ܴ���s��쉆�5Q;L��XuS\s��@~@K%��^Xƕ��B���|K�2��tV��r���1պ�'���I�r�b�����ƀ�݂G��5���"Q��C~�^Y��)���"(�+a5%���Vۡ�߈��v��nyk�ã��T?�L�2�J�4xb$%��juW��+s��w�+?U�=ІX�1�Z�{j��ț긤#6�}� �Z��&n��_K<.~l�lݧ��/�jF�NDy4��~� $"� �:q�|�@�o�a�K»/��<X��0O42�i�弰j�v뷐c�Ypp�ոh�$Mۂ��7�ږ)CWD�Sɜ�).�mQi��m�Dn������!"Q�T!�G�My#�*�r���0I���,
O<�r�Y,��h~���a�~&��@��̳��6���۽��$It����_%)�\�E�i��>q���"�,]�,����F�1�J8��ۊm��?Y����z�,1���@�?žx��V5���Z��a��r���t����L�m�΍��/%c,v�����B�?-����� �u�,"����t���x&�&;om�+	��xz��D.L>����c�-`�:]�Y���$��$c�ڦ��ٝ���u\�����^�ZY\�g0a�JF\��2����G��Ð��t���EXN�}<�� �n� �k��ȅj�;&�
lf$�D�Jfm�C�T~}]_� ���\�}>Z-ڗr}yʹ�T������nLҌ9���0hwHmj��oe�S�
ȑ@AFd��ޑ$���b�c��o�k{>���|x��,�V��q��n}�!d"4�S2]�[J�%�k�L�\�[q��c/}hrǬ@d�B����U�E�1s�*��*����x�3+맮fG¦3҇�T�-Ȭ=.���a'�}�-����
�i]"��Dd�\]W�3�ɕ�B4@,a?Y�e6������i�Kx�Q���6U��j6P�u}��2���R�,�T��L��z�9��:U���^���m����<�pj/^��A6Z)k��{5�US��i��s��A^rPt'�Η��f6N(���I����-hƟ�R2�9\I�޼�@�-_C���ϺeP�Xb�-Y���}㴡%2��$�Z ��m�}����(%�ަcH>}у ߬ws�QBϑ�������"$4 ������ހJٿ���î�l���.h�Ү�����0��
`ȉ��gw��U�#����� �dq~7�'̌W���K��,v�۩���n1m��������Z�hl}�mjČ���~�Ā	C��By�����u��c¬x|hz�#�-\���sk؞��V<(�"j�:�&#x���
gN�f-�3�c�I�f@��4*a��}DBB$�AZQ빜6q��0fk@r#��vxE��P�S-R}rQ�T�P�gZt.�R�Ɓ�t')��#W�~&�'d�|��ji^>|B�q�"�vm����12��t�-gj�UC���#�iP/Y$(���*=����,Gy"�#�8��Ҟ��]`����i�]/������<Zڔ��_�2�I���e,�㶧��>(
xjL�'3?�'mpH	j:_(!� �e9���b�Q@�0`�0��u�vW�|8 ����L�
���o�}Wl��s�bm!q��=�]����s`��$���t`��BY�r 4X�����4�W�)f�]8���ұ�N�ETR�V�{���:���CtD�7�_h��?}�\H���\K��@����]���7˿:�������\�Ĳ�+�e*�W�D�m���Ԣ&M�7諞�[}ӷ8B:��gĀ��>ꍞ�����5���|��z{�!��u��;ӵǝCE�s���1e�&����q���%=��ɏ��ˑ\f�vx�Ӭ���p3�]d�p6�^I��b����vZ����^�Ǩ*T��dRǇj��!�>{/	��7I�8��`�@pbt
��a����i>�/�b�Ԙw@�RX�g��6�D�t�������N�u���/l��N�,�(�*��B�ҝ���w�^�S�^�$Fu`R��8C��:d�m�ң��MA���su�����p�s���?��#�ρLBtE�0V.&��rY�РuS����C}zH\O���+�sPzk�C8t-L�5\���Ita���p�an�5GĆ���Hc&��H���G�$�Ԍ|��a�z�1�!�M%}bܕ*���(��4I3'Qrq�ߖR��W������[�����9�RH�m��a�^?�T ��i�p�|�dB���:�T�����qN	���%�5 �����ʕ��	s�u��n:�*����^��q���c��u�!�O}� �/@����6��n0k5'��0㖿Y.�K=�,k@%���F��3����X���W�RܢH����F��=��R9p�A�	I���d�s�vM΃)� Q�@Zv��+�"�� #�C���g/dn"%Ϭ	u=�o&�n��$����d�D�b��z���,�p��dX�>\���ĘK4�pc)r���%�P�"	]�A6�N���cF����eך�w�=F�<ń�y��d ^�e{��%���Y<�^:�u�RƊ��J����� c2��E��p��aH�$�J�m���+����0�r�/&a���*���<{����OO�a 8w\����6^zni����cNS��h�*���lpu3_e,w;.�S��j�H�m� u�s"Ӿ]���q	6��4���u����X���˘�'��z��4sJ��~�6
�A3�A]��o�!Q���d(D��7N��2ʟb;~ A���	�b�;6�I��I�PX�l���n���0��	����VG���:QF�djE�Xlby�5��R����a�7�>l�hh?�J�=7�:�'����MЦ�A�:z�|ʒ!*=�05�/�t��F��Rgk{zZ����O��r.�6o�<����yR��}� *�DS�IsE�!6.��n�7q�Q�Q.�����K��z�]�����f��Gx���
�����RSw�z�~5�~�q�$]9a[��=s���g��[tqȰr9�S�#��W0<�8D��m�v���9�~�����¡45���]eQ��c^TP�������T+|&Ƈ�V�E���|�Ln	SF�����L�
J1��b�s¤����A��s�h�Ѐ��jX���Z��E���U�?��6���{���O�{ _�'.Y�l�9��D�F݉SymΙ�9��$3�"1A�:���|��[oR�K��ۚ-9Xz��0j�{2j�l嗫���A퐨�zTAT�z�h� i۝:b7v���D�����3��#Qįnmk�;��A��8!l��*TY��GkA�#�r��u0��/�H
����m�YgOyhE��ߓ~�i�@kE����.�"޶dZ,�0tT���\�)#��E�@m�^��H����,�;���/�,qJ����=���I��15T�U�1%��@����s}�V��*U���Vf��U(�q�AV�L%x�Έ(S�B��,�����`�E��;-/%����p��"R���/dF��CM��iom��1	�]����].��J�F�c�A���u�4��_Z
$����|�	��#�0Ə��m��㩚5� ܢ����������]x�ѫ����!'E3M������n�u�ƅ��@��;A;7���f�����K���~x}1�o56͂�\��YZ�rX�I� E���z�Y�����{�Zh���j���oj�����,��F_����t�B��~�o]�\>қ�|��3��Q�V|6*��F���48�2�FJ�{�����_�f[ld0���!h-��@�B!y��0�Ƒl���Ņ�ꃶ�;xL�%�§�G=���3�T�Ts��K.�n�auH�}>z���R
�5"�L*d4��W�~t3�v���YO@�8�t���I�ͻ�3iRÛxf6��ή��R�P^����%����,'�������t9z�U���y���O�����v<���/�E<(9Z�8C��3�p���H��N�7A@�$PM�Β�Tf�F"(x��d\R���z�m2\��X޷���;z-Ҹ�&����E�3�1h��R��92s/@�r���uQ��+�}鱡6�(�a��^E�>�J� �Qs��1�iZ�m��ܺ��4����� ��9%��v���9��� �~�Y�D߲�a�+Ȓ
j���DOu���Y��mU�(��3]� y�~2G '�c��NK&�a�vh����L��%���~��Ol��.j?x����4Ļ�I��V���%�h�ǠJx�;�z@ZI-7�I�95v�9�!V8��}�)����#��`�jNk��n�M��>f;�z��Ч���D]B�� Z,GR�q����k;�o�?x λP��oR����ь�G2���.���4�/�.���W$�&v�yd�i=��$>wj>qF���1.�*��N�2�h�t/&g��Cϸޒ~ۚP��(�-�*��Xݤ4@y]�=�Ӏ��Fz�C|�`q�&ӄ��/<���K"<Bh��.�����I<�e��:���{�v́
���L�@*?�hGk�+j�2�(�0� �T�c�gk�Q{��`�s��є�v��H8�Jӫ	�\/>֣#��C�l_��Lv!��=m����b���,�l'$����l�G B�1� �>�:�:�O��2)��R8�����1�N)�����߃ݮ��d�5��D�tY�Z���'>���	��n� ���X��=����˺P��p��7�w���'Ƿe���x3v���ѵ&����f�[+ �(J��GtĻ�ق����	�q��� |�|�z����j���vO��8GǣnQ��	�v��4ш�*2�.�=����b�f �fݸS�..�ȟ$3ȡ����8^$�=�I��!׸vgM�PS�ł�T���R��zj�c�\����b={*���@��`	[�b�g��n��Bj�_��>���ֽ���2�m]bg+.�6_�/t�3��r	N��ԁ7]F�D'	,�*��B�55�J�Uw���S�p��h`8^�:���J��
��`d~�ԮTw�p�k�ˡ?sQ���L}H��˱&���Y&�u���qT�Ql#�0\@��O3dz+��z��d8/2����״\ŠX�a֏�pi��0����H�ػ΂���K�� �$#�Z|,h��u51Q�M��Nܰ��e�c��4>I�'�y2��xR5yY�)�H��������J9,��Hz��\�^^�`l �r������?����P�T�Ĳ���	k�%��>��1���p2OD,����i�i��*ll�芥'���V��m�u�2I��f �� ���6I���)�kP0��z]���Ԇt,_a����"e���,݌��g�͐�#w�Q4��u�̳M�\����0��H���M�����m���4�v�vN �Wл��CVn��<0n���D�B�ֆk*�1�LՅ��d��b��(z���g���F/P�9;M�1�٘��p~��rS�%����]wI��k]N���Na�U��%twR�Fh�Մ
����7^���HY_�w�A<4][:U�PR�󠔅9��0c-T9���HpP��H�J&�/��?��]b�!�&\�ـ�/u��7�O�T����\�}洈��6Y�|ig��qKi��%�m*lAXl��_ y�;)�8�J5H�8h ���"N$X���1qQ�_�F�;�� C�T��X�F�˳#'J�f�Uo#4���d�A��]s������?�lD٦x7�b-�b�y� �W��$�/�}���$�dI�!�X�e<��Rn+]�0S�
���5�������\�"�d�̈́�/��/s5}J��ꢾ�ܫ���P��Z��8�7:	�]آ��=8ҵ���W��!e/0�$��ojoF
���{��'�a?�c4��ql9<ST��t�E�����C?�7���0.���.�L�|�Ҁ��L�������Q��f䫪��]�ĺ��y
!�>�۱��F���ГS�����8~��.�_{��@��8�2�0�E;t��r� 3���̒Y}�Ӕ��hR��B�v�9\Հ=��=��5��ј�Y�y�q^O06�ߓ6����+�7���M�V�	�U�&�+>nM}�y�����qL�
�J��b�⻤�鱗�.�s�-A���K���RX���Z��4 ��>&ո��^6�}��֐�jW��M_A%�.4�glSH��e��F��yȈЕ���$Nl�"��-:�0|6�o��oK��c����X5�0�d�2�=�r�Ɓ췖�C�RO24����hD<	۸�7�߮pDY6�&[Q�k�Q�m&r����@��b��iT�GU}#�r7?�0��XJc�
Exӽ͉Y���h������~��Z@&4��O��m�ޑ+�gIt�����yC)~��E`�u�/������ a,���'��'Y�J��Q��t�⬢Y�0c1`J�@-��n0�V뗆AӋ�k�h�L��|�L��΃�������������4���
h���O��k@"�V����f��.|��{m���	&{��苖
��.E"���c'�K�0"��q�̚>�$�k}�w���S�
��O^�1V���A�!�����π���f��sF����;��+P-El���1�688n���!� ����;\�3� A�f�i2��P	�y�m~s����tl�=1�\�aZ#ESr3C��[U8��	�d�B��6b�h�0j�����ɣ���%�FZ�p�G/���û�L	o�*>�fO|����b?�Vw�މIώ���_4SW@2S��J^������2[gЇ��fh�T�@�K�B�ju�������`I�!�v�wx�����TG�����HT$��Sz�.�p	aЉ}����
�Xz"���do�qWC�3�C݂��j@�0M��-,[͖��i�  x;���F���yP[F�*���϶�j�u,b��L� 9_<�Uc���`���?��Q]<7�/� }7VZ�%d�������ðn�)�A{:KP���΍�f�^�(3�E�����
��Uet���\M�޲'�~�-Հs�A�Ⱥ�f�4|�a|��㪟�2Ν��-?Ȑ�Y�c�}��Xq�j([襦Y��>3� U�s��χH��Hb+��V!4V����%����O?`��1M�b}�Y[�H�4�M+��&��
��a��)$������UgMg�nH �0~-�����~}KA6���!�vC[ɴKo~g������;��о�l���j��U��T@���ķ�],��7���5{�ٙkx�.z���-ѣ�t���V	T���.����(#�t�-�NF�Č������f6�D�ꖮ�Z�xDx�pB�Zú��ό�'��k6�l�ʅ�x��PϛRs�������4K��͖.�,��7$z��V8�"=W�&Q��dw�����>r�sq�	���`�E�h�2j�tj>7g��C��m��MP��(��P*3���\�y���n�$����`,�ӟ'./�>��c<}���ɿQ�dI`Ee����-X��{�
�SL0z�?!�9fjj�%�(��? !�k�a�B�WQ�?A`G?N��ӟv��8v4�$��s��~���l�JX�V�!'=('v�� �i_��G�r$�A��9�	aB�i �(�U�d��uz�8�)�\\8(Ͷ���N�dȠ�����;J���v�p�D3�3�U+���c�S٤����]���ts�Ӹ[�:ܧ˵��6f�ؒ�f��D|���~e��#
���[�̶b&���!��[F��./f������t;ɞ�Uj������|�
#zq�EW
Ա����j��i��d�G��vшף:���=�#��?����f�����(��l�3��f��^������U���Dv�X��@�=8;T�H�R�j��u��K��t�
{%�Zʛ�����`$�pbj����n�}29���D>�_����������g���6:��t��DN�q��������,�(*��dBc�<��pMw��S��آ��`ȝ�8y�6:Zk���(���;��t����Jp_�4��?���}a1L�<�f-	&���Y�M�u� O�B9F��f-\{�SO�J�+�Ǉz!�e8�V�֍�R��{�a��p��+13�N��H�eû�)>����ڷ$^�<|�$�pi�1x��M��^��.��m�^4yi�'�����Rp��I��:�=�Qp�v+H9g�DHs��W�y^�� [pޓ����<��ص���T0����	w;�%u���� ��̚�K�.m�G&B�d~*�g%�E\����Yo�uycR��� .�9��H�6��}��ӭkkY=���ߖu���ˁ,������"�}�W�V�E���ߊH(e���D䌖O�q�H��&�x�8����i��M����*��NI:v�[Q��v(�C8@��]j�nؾ��E|O?�ޢ�����@�?d"�$b_Hz�����|ۯ� �4yڌ�N��e�p�w�r��%������w��N�Q�w��(��w��FC�v�E��ܚn�^�����2d�<O�:�R||C���,����c(��`jp,@H�J�����s"�h���N&WX���Ԁ����{OED��մ\8ٴ#�:6T�i�W��,s6������*G��l�ߔ_��;$���rI�H]#) ��"ɩ����q������S���U���MX\�~��P+'ō��0O4�����W �1A�BF].���1��w�0D��7�84(l�b��� ���?�������I\X"~���n��0ů��o}�L�"γ�X��dMQ��& �58��|4�W�M��=JWXuI8�3�8:x
1������0���2�!�A=0k~ʮj��Fe>]ȶ~{��*���t�>�䬉 <�L�o�H�N9:J�x�RXn�?ò�/_�־�m�n�G�;�Ђɨ�i'�pE�]m�+�5���\݆֟L����)9S�c3�t��~ѓ[���W�F��3�+ɍty�c)�t�^ir/���5�͢R�n|�c��ꝫS���R�.�悸�05�4������^JX�:¢�S�t+�h����Vl�]��F��Gr�n�f��O�m3L'�J'��b�q��T͗w�Ls���<lǀn�>X��LZoc�X��y�h�ua6�-�1@�%��?�_�Z.�l���� 4fF�_�y#cG���*$iIm"'"�:���|q�0o��K�-Ț��X�4�0�,2`l��M�'N���#JC�0Sh�w-�Ӏ�7l�����D����#��G�QzFcm�8���]�.Ą��WT���G��S#翻r��0z#�e�Y
�$���
YݝZhOb���W�~7��@��=����$e��lP��t�ٗ���)ّxE���J���>1�꽲�,5���"aJI�C?�1�Y�'0�>F1�"@�~��i�VF�"˾�������Ͷ'�o����L[��~D�@�]�4�Ǽ��V�ЅJ����h��f�k"���k�:���&�mv�	at�I	9���.]���RcB�}���*��Yk��B`$4���r�{ٮ�������L7��v�%�������ޫ�0���Oz�G�M���F���E�h�.+u�љ�n�||�FȶI�;w���{��f�S���uu��^~n��%����{\��Z�*3r�Ҵ����TAm��ҝx���7|hȏ=j�4id�d����bȖFU��ޢ�c��$Z��soS~�>�Q8|).���L�Vr�����W�R�D4n��2γ�J9�T�_�f[b\��t�Kh��S@��B|t��ّ�'��,�	x���sx��g���7G3\.c��T_F���@.~��a+�}�so�B
 +"lZ�d�S�W��	3�0;�SR�@]H���]���q�iȝxx�_q���&�1AP����E����E�,�������e9��U��E��E�����<@ʊ//�2��Z:3-F]�c@�>�ƥlA���PE��Έ��fG��(�++���e�
)�0S]�d�\�Z�ޭc}Q��-�OҼ\J��A����v������N2),���\rȫS���t|}���p�(���TI>��� ��s�eH�HL�#Q��0!�4񠌶�j���ͼ
�M����f��4�l��y�览�!Ȕ
 �Ⱥ$�����xRUB�v��? ��$~(�E��;�91K\s&��vKQ��Zʎ�P���y�݋�Il��hj5�����1���Q����4�Ʈ��5x�Arz6'4-��ɯH�o0V���3ꈰk�#�r�
��N!٘��=�-f1�J�E}u�ID�t�B��bZ�^���؏���k1��%�qxv'.P�o-R�U�?͡�Vl�87�.���ƒ`���F�=��W��&,�OdJ�˼;�z>mEq�p����b`1���2E��t�v�g;T�C����4�P`�(8�*��0�Z�"y�Rn�	��"^���\`�aqӺ�r/2¾�>|<�䇔dվ�-I��MeA��4�<�lJY
��Lk��?�IDa��jK9>(R� <2�v%����Q�W`�*1��2�vh� 81>��?tR���Y�l.�l��N���!��=�)�AF����"E�$9��EE~�>Bj:� L3�p��Epo��2)�y8�-��Ñ�N�#�Ku�����y�c�|��쫔YD΃��P��P����M����d�庝��T���9˰�l�{��M�&��4�^1e�*2E�n�V(��׼&^*���!Q[afJ��U���>�14���A��'���>�+|㸅z�ƒ ����i�n�s�d���ٰWؕ��<����l=�o��z��=�fӜ��,�>Y83����� ^ڑ#��x�W�Hv�ߩ�����Tط�R|^j����(֟Lp{ �p��t�i��`?��b�y�i�����zF>�x��s�Ș��`��Fg!�6��tU�Z̨��N|����8u,�X*�B>[���n�w�O�S�i=�5��`�AO8��q:��$�c-����s����w�
ޑpKG�O�?iĳXZL�PƤ��&�Y�;%u����3$�Z4�
�\��OiQ,+���z|�F8����iz�SA�V�@aL�Rp�V��&�$����H�5�����4����$�3|b��k�I1�ZMV-������[�#�{.�4���'"���0qR�I|�.��Ub���X�Q{�9�<H�%��R�p^P˻ ᮓ�`��X���V�FݺT��P���	�+�%0������o�&^������2�_�*"�Z� �4��L�Ԑ�uT� by ɪ����i6������k����pP�P�7��B�,<��{/���'��F������K��1���׫:ڳC��$�:`"�7����:M_b�eh���}v��g���1��CSJL�ط�n��H������_�q׹盚��;�d=�qb��3z�A���|$ȋ/�����#�|.&p�W&r��j%rB��ӳ~�7:N�
�t����Y�(��wHDzF֧��E,�5O�^��R�����B�<j��:K��RW%���{ԇU9c#�P�V�KpƕUH9�BJ[����I�A�Cnb&R�9�;���m�:�0oO�SL�Ի\N�����6OiL����%�X�~*"u{l!�c_6r�;�֊�h�H. �J"DOQկ@Pq�yO�|�#���$�
�XR���'@~~�O34$�&�O�<��MAD��]�����i���P?��cDO�V7�#�bL�X r���Z���sn���E9IM$YX��b�:Cn���0�����}���[�Ύ�;*d����=�s� 5�� u������ϸ]�~�X3�.}�:�+*��Q����]ҫP��o�!�sX0�K�e�TF��#��{�g��W�Y�o����<����jZ����՜mx����ܿ��5� ��B$eb���=O��k��F]HT��p �WT�ѭ`����D�BS��k���~������2lr�.�9��lB�-�t��Qr�����(���	��^z\���Ш�Yt�I�9�3��5����b�௬7^E���ϸ�*+͹Y���VG�o�������*n����/�Ƚ@�Lc�J�rvb� �V�ܗ�Ms��C�)�.X�CZ�yֲ©�0�P�6���Ό	�ତ�Q_7��.��l�h�ě��F���y~]��j0�$�F�"���:�p�|�-�o#�K���> X��0�G2�W��(\�bF�y��Et見V1h�����Se7�����DϘ��\��C�Q���m�}����ES�T�T
�:G<�a#↔r�k
05����N
;񚽃!�Yu�h� �����~�}b@��+�X|�|��G���t%���R)4�iE�w��e{�ҹ��dL,p�R]|���J������L(���h��Y1��@c~�d�V���\\�0���^�R�ԓ����L�W��y��ZL�ά�����D�«8������>��a2�"c�y�`4�!e���mQ`�	��'�I�� 2Q.�˱�w�dc]�׿&�ǎ�b��g�$Ϣ �m���	�8�a�G�g8%���U��hN�S-�϶����)yK�JD�����~E�	�ie��l?n�4��"m�q)�;�`ŗ��hf�]`�6����{�~i�P��S9ͳ�Z\�ŜZ0�r�ߴ��J��z�����"E��-sh�<j
��?/Z�?:����cFP�^���k�s�\�\�o��>c\�|d�FԘzSVmy<�����ӭ4�=M2I�~J=��W��0�[]����h^b~@��B�����hj�����0h���,)0x}���ScG���>�DT��m��7Y.y��a�l	}o .&7�
��G"G{d��VWy�3�=����@�k��"!K�LN�i;x7�����O�c�P����`�l�j�� ��,�5���JU�Fx9!VU�f��J#��O���<{}�/�5�-kZ�`�����S��w
��w.A��P�}l΃�f��|(���������gd�a�.,\�K�ިg��e�-K>ռwb��-�ą!��#6��2��D��i����YI9}z}7�O(�UͦO�>�vr ��:sp�}gg��_9�k�4��
�����Jҍ�>?�, �X��V����߃D ���
{��u?�Ӈ�.{U�����k J��~#�r86����Kw�r�}�v�Z)��e��w�������F ]l��j����b���l�������9��yvb�O�:x�t�z���-�|��8�
_�V�����(�&#�#����}N����C���f,Ռ�������D�}�B�Z���"��]��k,z&����x1��Pd�Ri�.{�ա�������.�[���`X�X�-W�i�&��d���{	>h��qW�ۍb&R{�{x�2 ?bt��#gֳrC�Q�����P�+(*��*)>O�5y����� �@��T�`��,��G�/�e�$Q<�R���
$�I��e����O#)��8�
���L�L�?W�f\X;j�l�(�� W��^��E�Q,("`}6L�±\v�C-8�gO�Zn�\6�4��i�Pl0���ɹ!��=�p��,���_����&$t/`�&;��%�B��` s؋-Q��������)R��8^z��q�N:C>������(�W�*��DDi;�KT�����H��Ѧ�ߞ
�xԘ�I-�p�˫R�j�zJ��Բ�Y�e����k�G���&���藍;[|I��$��)��l��e��M�т_���7|��zg����G�'���	��_vW�K+�Z��#�xc=q�}ٵl0�7#f�>�?r��e�3.z�\�^��~��j���#�vN�a"ųG\T�F�R�Мj�Iq�&���m{)#�QUm�$��`Zib`@�TU���"7�0� >�{���QE�c7i�,eg��6��#t�*�C�Nw��H��uq�,��*�r�B�����wS5�S����gC`>:8��:P���>���9&@�1�)�g�e�ypՙ+�j�s?��3s�L.�Y����&���Y7J|u?���Dx/�
�Ζ\�P�Ox	+��/z�8` �foH���1Eea�p:��!���Y HO%���4���}��$�i=|��$�fi>1.��M����E�־��V�w4�	�'�P���R&^�4��p��G���,�29�s�HK�Z�M�C^��� �q�ܴ&�s����g��S�Tf��u	-<%�䳴����P�$��O��}W;�Zj�*}�/�9�����O��u/%u;� d���66Z`��Z<k�����+	��7��,�z&�v�o�3�4��Ì3e�>��������(�F$�>а�����5�R %�_�>M:���3���zv��^ s��LCnt��S%�n��&����P�8�
$ȹB��ն��dXنb���zo	��㖯OH�*UI�BY�7p�W�rw�$%M�����Э̜N���'�����C�)wÒQF��h����Oo^��ґY���A�<�A:��R26`0��oc�6����p�/HTiMJ�?t�g;љ����D�&M� ��ol�(t���O;�l�\���Y�66J��ix`V�����0���*�>%l\�F_��;��(�xH�X ��<"�PՊ�'q��ӫ��ᯖeo�X�.��'��<��n�4_����<D��EA�M�]�$,�����m��ГD��s7����b�ZL -[a�u���$���{I�U�XX����n<��0�R���BM2�i�`=w
d����t���5����;���M�ڪ�N�Ř����)N:.m�������&أ����!�g0��E�`q�F��>��{�V���Vʦ�9��"$�<$j�e�#�Hw�kW���)�5)񲍩P�����o��=�J�w������v�f��]#����s����ۊ� ��:�S㣌�jC~����FͱS�)�C�C����P�t�tBr%��x���C����F��Y>��S�j:�do����5fS�I���J��^@}Q��~����+�*�
�wV"R�e�}_%n��J��b���bL:��JR�bk�H��������s}<���Ծ��#XU�Z��e�,���˸��-6��l���D���^��_�%�.���l)<�6��Fɵ�y�w��%��$�c�"��:f@T|��Uo��K�%��W�Xf��0�[2Vc8�����K�7�@ż��ƏhuO�	G!7bKAp�OD
zќ�;�_Q0]�mW&���$�$�Mi%ETE~cG�O�#�m�rH2�0�&��^�
��p�^�aYSl�h����˛h~�n�@W���&����"@�Wt�L����)��ZE��Ԁp�4��s6�,��������vJ��5�H�g����r���137@���_	�V��A�Kk���������-#�L����t�e����ͬ�\U�L��(�� 4O�\�,"�O����<�9��c�m,��	��=�ۖ���.�i�2Mcx�Y���������K��$jn��h���d�o��b��Y��l5Қ�<S܎|4�Q���$����������0���E���᤿����n�	X2���,)�;�WZ�qp�fk��q ��J�~d=������nq�\�XZ�U�r�a�F"��@��D9�S�F�gC�h�	�j��K���z��ȘmFK̟�X�Ӡ.F��oI�>>�Z|�5�3�Vhz�Z�i����4���2ĠeJ�T��P˷([X�6�*h�hM@�*B����髑X@ �1T��A����x8<��.��G)u�#{T�1i�$��.t6|a��}*��A��
���""� d ��W�3�jk�	˽@�� �+V�S��'�i>��x�J�������PJ���{��%����,�O���	G9pC�U�Ԝ��o�;4�\y�<�P�/ep�(��Z����c4�4�:���`A,uwP{#K�~>9f�g�(d��Ј�� �����Y[\\�ޣ�}	-M|���꺃t�ҟ^|Tށ�����2ߨ��^p%�����=B}U_"O6(,<�Jm>Dp �$fs-������َ�ܦD4'$��T���^��4�GǷ��[:��/����?��H
�S��0z	��s�|PU�{%�� ��4~�[��دn$K�M���"hvԊQ���8
َ��s�L���Q�lzCj+f<�=�ħ���}���3��F��
��x�<z,tO-��%zjإǞV�g���h���#��  �1N�Q�Z!��P��f'���C���Dɦ�B�+�Z��Ԝ]u��)qk'����$x� 1P x�R�'tV-Ρ3���nj�.�cF�H9M�n�s�WL�&��ed�^��q�0>cJ�q����e���C�2�tG�gq3�C�ă��d�P֭�(E��*��9��EyI9�?k��~����<`]�L���/(),��V�<.�ꔚ`��'Iq�e����j��bGa
f��L���?�W,�j�x(�k r>�l�c��ίQg̠`b�޽Pv��8����u��H��31�@�lˮC��33!8�n=YE=�G����ͳ���g$���{(p��ZlB �� ���ئ��;����u�)�L�8�����q�N��� �)��ol��2��!�D�F��U�,�1�Zo��S������D�˦�GH��zҰ�,\�u[eq ��Qz⑩��ye&O�R�[�L·��]_Hħ��E%מ�y5�ݶ���|u�z�û�֙n�b��Ǥ� �Zm
�u!=���j�(���_=Lg���s����f� Z��s�����34�C��[�^��ɜ5}��}�v�b��D��n��T�7Rrc�ja+�HCf�E�{�qʬ������`u�b�/��.K�˹r>ݞS�)���ٱKg�6��t�@M�޳/Nr۟��Rp�0�q,�*
�B� �6��w�:|Sڻ���?7`��8�a :�F��)$�to���f��뉮��p���#
?_�E��Li٠�7`�&�<Y�x�u���v��,��\,��O��>+��z2s�8�a'���r���ya�x�pՙ���|�_�FH
5��:������X(-$�[|��a�1�N�M�Bh��U�Q���1�L4*�a'X�gzZR��EZ�����9ĝ{ 9�&H����H��^�� �"|��|��?|��(����T{���8	�l%� �1>,��=��	.0�h� \�UF�*���v ���hL��3Su
��v�\ ��Ԟ|��6����i�k����fO�E��r��,rîq��js���׌Nٸ���]���M�=}���-ȳ9�7�K��M�m_)����M������Gv���lgЧ��C��ʟβni5�0na�Ɇ�t�����q�dsdby�ozJ�S�r�����%�ڝ`��Dp�wr� �%(H�Ip��H��N�vq�*�ڨAa�^��w>5F�1�����kp^�)o��f)�c`M<�u�:A�6R�K�qd@���!c�X��Op<��HoJ�JD#�B�`���q�y;�&HVc��x��B��:��O��ZG2�\�&j��X�6E#�iӔ'�]Rզ -�*�(�l��=_l��;|劃zH��D �n":���eJ/q=���
�������X�����<'6������4�2����#�{A�]_���:k��'\�~D��7UzO�b;� �FQ��}��i۽��QNIæX����1�n��d0?�w��E��^��D?mxӞd���ˠ)I�5i�o�V�F��]�څp�,wF�1�$�c:�μ�IK��-$ҡ��|�!Q8k0<K��[^*Fv����:{fc�MIǦ�{��]��<�&ݾ`���_�E{���惚�f��h��8��>�T�8
�ZRгH'�ҸJ��~]�c`��d��Ɇ�)�]����S�s���;~b���K4lh-�$�Iɞ�T唔�t�/;r��*�S���~>K�?��T"��u��%ף�Y�)q�5A�xф�����^;,(�Kh��b�+�$��_�V�X�A$�xn�t������LU;�J�Q�bF���RؗH��sx���M�:���X4��Zy�8��+�*���F)�6����B��V�<֡_-��.�)0l?	��ъ�FĐ�y4�,���$���"�c�:A0|"�foYqK������X!�0�DW2ю���q����Ő��d;6��AWnh0��$Z�7���KeDE{���=���ZQ��mM��&�k���tDDT��@Gr�&#�t�r�.0��z�G
1꒽99�Y��ch ����mb~H��@5��A�����ISt[����-Q)��KEL�ԛ١ү�f�N(x,�������9�JZd�=�U��\C☘(���1Lk@��оZ<vVW!x����f ��T0���C��hf�L,���o�Q���/����+*�a��Tvc��I��W��"8a����W��2&m|�	 �+і�9�.n�����uc�R�ȅ�{�#̆($Zd�cFiٿg�׶A���]�癚�|0(�����mz��N���+��xSݐ4�NEz'>��9��~&n���+���Hy;�nw��j\fF�Τ��2���~_�q�6���)T\*��Z��r�V��G�-�%�����iҮ׈�"y-h�j �o�N5��P��3p�FF"�޳ě����#oİ�>ғ|�����5�Vc�������J4��z2?�XJ����ͦf�U[S����ӻh��@D�B�pz�w�����E�̗��<Ƕ�5�x��Ie�G�1��n�T�8��t�.o�Za<φ}��W\8
w��"�޶d[jW��n3��=�d��@�O����k�r�iy�Zxm�����u�mP��Öo������?�,N�?��	w���9˅�UObl� ��� �7q<�C�/ �}#N.ZK�P0
�����V���AgsnP�!�y��fX :(���?�{D+���x� \��ޞ�'b��-�{Ǽ�����=��zW����YM?� 2:��*���Ƅ�OR�}0�V]n"(�BU�EG�>��� AiusH���s➴���?�4o����� ;0;�.�b��N��)�4�߹ݷ���
1�����H�	̝����U� ��Z^` �2Q~.�Ja�jTK��c�sc�v��ɴ7܎Ӽ������iKݼ��l�j������.9�"4�����/7J���x;�z�J�-~���`�Y�@PzV�N�D�H���#-u{�N�k5���l��8f"�řV�J�F�D��B�0Zs�}��쵏��Hk"�P�6�Mx���P;��R_�%1Զ�n}��	4}.�`�ƣՓ��5����cW�N�&�(	d�뷼��>^bqgy��k���/n��2��tV��g��C�W�EWSP��G(`�*O���;�y�ܭ��uN�ܦ�
ϼ`\���/���ϩK<i�J�5���H+I�eierB����u�
A� L��?���R }j\3(�JV ��Y�1��w-Q���`��*޸
vy`�8b̫��$�ŭ��K�FlfeB��!���=:��b�)�U����$��OJ����B{�X }R����]ڶ��yP)�1K8�s�����N�!��ك������X��\D�
��A
*�a[@��B�GK���_��.�����N簾 ˡ��{��~����d̲���eL���W�}_^����&o�m�Ŝ[�o
��O�8�%��f�]a����8���o�;|4��z]�����Eԝ�r�?9��U�������{�C�-�n|`='E�+���m	�f�����x�o�3O�u�R�'^k6�p�5�(�%v�^���)׍T)�-R�pj<-����̟��1{�[�$���PN`��RbV$
�|�i��f	�>���քv����F�V�g�X<6�s�t���yn�Nm�8��+��B�,&�3*�y2B���q)�w�`PSՔS�F8�`��8��S:F%I���B��ؔ�g��=��)pK��㠉�?�����L�M���[`&��Y��ju�Ǻ+��%X�j�@\g/�O:%�+��Gz��*8�)B��>2C��~a�Fppk���↺�mH�d��UY*�p�3�t$Jt�|3W��\��1�NM���7���IN��Q4e*'��u��R��� ������=�͝�*^9S�H��T�CY~^aۃ G�x�el�*𾆃�����T�����[	㼧%a|��LK�|�6ʷNk������PB-*3���1��'��E��u�fX�f\ �EΞw� 6�o����k�=��j�᠒ԭhp,ط�l�,��;��B�Ќimъ4ƈ�j���x_��|W�4jU����k�h��޵�U[�M��+�М���v�� �.{�b�ZC�(��I`BnDrs�kfk��� �ݹ�2p�,�md�c	b�z%�鼎ɢ�Mы �����㘭H�p�Lrmd]%����~���WJN���X9���y�uw��$F����11����^�}'�:��j<���:���R�߮����&�jc���g�qp��.H�K;J�h�����	ȨR�&C@�L�������U��O1B"�q\�`-���6@�i.���2�}���1*�2�l�4I_�D;�֊ކ�HI� 1�"��Q�@�fqx
>�Mb���W���XH���:E}'����4Ս�� ����AU��]��,�(�c�����D f
7�.,0�b];� �R��� ����c�k�I��X� ����~n���0�_��'h.�8����)�O�d���B����5$���q ��C�
�`|�6�)�C5���:�OV����HR#�G��3�!��b0�$��VkOF�/w���{����[P���@�>�<Zk�[�o��46�Ɯ� ��+�ϲC��s���ٮ��3�Is\d�n�y���\'8]��!�L(Ɇs�� �u̷Sd��`
J~=_p�������K����O�Wt<rG�.�d̹q��g�O&?�	���ű���$���95XNѿ~��_^6�:���Ը?��+mv� 4;Vؼ��|���"n���@���q�"Lp�_Jq�b!�=ė�� ss�4¨���ZXOCVZ�X�g�x�e����Z6�-=Ν=��>+H�_�p�.{��lz	v�l�qF��y�����$���"dc:@
|]��o��K���OB(X�7�0�;2L�&�,ׁ糐J�6�Y���h���?��7XX�&l
D���-�O���Q���m͓��A����'�T���G��#ӛ�r�`0f���P�
����Yɺh����_�~���@͑N�\�������|�T�t�?i�~�
)EC=E��Զ�[�*{\�):&,!+g.�!��KJ���P��&�����wq�1��9@4=W�U��V����(����ψ��������L�W��j����lI��3}��Bϵ�<���e�V��R��"t@����Ƹr�຃ om�9(	M�&��ޖ��A.���jtc��ֿ���V=l���}$�ej�^�0�z���䄸�e�b��WD��{�χ䳫��'�:���3��Oh����EU����=`�n�$���Ȣ�v;��g��f!;���J���~Z�챑�]���\E��Z� lrzk&���m��_��zV�	�
����h4Ej{6_���t�Β�FA����à�� �.o?�>�<=|�n�i�yV^�+�q|�>�4چ2�XJ�������[N���^!h���@!�B*�RK?����g�����=��x��d�GQ��WTK�ܬZC�.jZ�a��}���w�
��&"��<d�\UWJ��3�$�����@I�7*o����3fi��#x2���s�tNP�ȴñ�"CwD,��c�S~�9&�U
��g�1	����<,W�/�EZZ���ia����*_�p`A���P����tP�f��X(�z������ƜJ��Iu\T�Xޙ3����-|ʶ��"u�y'��UpB�&
�$�J�2��
�����C�ʆ8}i���(bi�@AT>�� ��hsc�W��A��LW���4]'V�����[���,�}u������CT�ocV�T���H�
�RȦO��$�p�r�U���( �%~�bI��%Z(Kȧ���v�J��rGen�H��(��O.�wR�l:��j!��������Qⓑ�#�G~����x9�'z"A�-Yn�ɛ\����mV��ɰW�e#5���4N��Ɍ��䆭�f
���V�PTD�X�B�$�ZN��ӃR�.xkp��WxbZ�PV �RڶC����z���.�}����ڈ�}���8KWq�&���d6�ټ�G>Y��qhN���>����R2�5�t��g���C�
?��iPLI<({��*�s���y����u���Zw�e�`�D��&�/J��q<�]��k$��+I'�re-������Xę
�LWx?(�_M4Hj��3(>I6 ��9b�쵉@[Q�t�`N�޳�:v��8����Q�>�����5�~l<���g:!�m\=�N��}1����� �$%����B��$�B��� 8���ܒ0�1���T�$)7�8/ Ŷ���NKa�o6�8i�eׁ��̡�eD:"B�< ����y�Ǥb���PpA�	ԩ�� ^�A)�˜tO�#�9���$�	6e'��1~VM����&�k�Ȑ[ͲZ��/��+��9�{���1�ѓmO�*C4|O��z؆a�����������m�P�$�+.��C�P�^ដ��=�`�f�s�8�f���P���*L3j���J^F�0����Ð
v�T֩r�u���,TD��Rh�jOc���F�{��{���b��U��`��ob�8��[8���:�y>�D���8;�� qg��6���tA��I�Nh��YF����,AY�* -4B�&􄬧�w$�SЍ���P�`o8 x�:�#�Ϥ��a����S�v+�pF���?U*��}rL��K�mw&��YH5up@F8%��UE�M\�΂Oի�+�I�z腌8��]����Qsa8��p]O��ĆF�H����pMB�����$�)�|γ��W��1?5MB���R�m�G�����4���'�G�p\3R7�����G긚�����9�ubH0��>��^� � �ٓ-m���5P�a�;�2vET7�.��{	>-�%�ʹgr��<<ʒ5���>�N��K^�*�0p�����.8��V�u�7��R 5���r��6kS���l�k���\��Q��_�,���g7�D-�������!R����EZ�a����/�a�Ճ�&?���}ʚ�ݓMˠ��Q�o�U�Pv�F�"v���C����-n�ᬦ~�!�����S�7��r#d��vbo��z !����&��ً��S{9�h��p r���%��)���Z�~M�N���� ����(w4> F��lj8ܡ�^����j-O���+<���:7�2R���|��r�c�P�¸Sp�|TH�lJ�e��V�5Y򨯈"&>J������Yx�p�NO���9\:��*|�6;��i�]ʅ�1u��0*�\�l�h_��P;�d�9&�H� 2�"0%U���q�z���ٔ��¹�vn,X�3�U�',�?�w�4	0���k��UA���]զT�G����~)a��D;�7�|�1�b�[( ^~��ƣ��_��FݣI9�X)����unMAe0���B�>����� ����dTÛ�ٍ�5���Č��¾v��;�q[�|Ґ�E�:?�����W�c��җ.[�y
�!�|N0r�Q��F,�=o-w{7�1�C�e��_����<�ϋ�Vz��C񳴜�:0��A���#���t~��.pc�~��)��J��� ]���\���A���%27��0�QS4t_��E~�ͼ���BȖBJ�T�g�
|Pt.Er�wo�	Ę���*�u^�JJ�d����c������5�0���rQ��d^1�����u�+9>�{(V�@ٔ���N�%n��U����,�XL��ZJ��6b�G�BG��~8snk@��2��Xj�lZo�BZթ��w�|�U6�}��������dF��_#Fg.V5l�)a���F��Qy�[�V��$�z"���:�o]|��o�v�K�k�����X��<0'�2�E��^�N��Ͼ1x"��׫h����Z��7�9�?D��ǜ����s5QA�m����\Tr���F�WRT�G�j�#��PrYER0!�$�y�
'c�����Y�hV[5�qj~��@�ͳw�C��޳t�ɶ8t���y�@)��.E����ѷ�ҥ]��l�,\��ɬ3�	i�J����n�}�Ә�RN�1�;�@ϼ��P�V��r����w�J`�n3E��LuLbBY�e:��7� �N=���-�D�r����?�M�1"�hI�L. ��Q@��.�m�	�2�P����.$YR�c)c�^ѿ[�1�d��7�$;���Yd4�u���M*L��|�����2xB�?*�"{E�����^Q����j��v1E0�'�U���a�n�HDC��]�w;��I�⿀f��}�"��n�~U���T͟��\`}Z��rU��V�[7��E��d͐�D�hO1;j���P�+�e�i�F<.��iOL�_�O;�!o��X>��V|Pm��q!VY=ɉk�ť�A{4���25tcJ�T�C����[I��;
'hJ��@< B~��-,��	խ�M�
���¢xi�t���G�
�f�T��T��1,.e,a�}[��9
m%�"�,�d�n�W�Q�3��V��@��1�G��͸'i�� x����v�ϥ�P{�̃Z� ��9�,����Hyy9�jsU����6���1V���V<g��/6��
bZV����-T��S�KC�A�ϸPLԷ�o	<f��(�^c�!:��q�"�w�[
�`\�M�ޔ����-79J��hv��0��0��{���@㌙T2��������2	K�E�%}�L��w(��=�;[}>Uc �R@s~��i%�jۖ�W��4�ش�����#���.��|�D��{}�������ϻ��
�j�a�3�?���C�U�ʔ��>% �!�~��ߺ���K�u�iDveڪ��ҏ	�Ď�n��]Tq�2�lUr�j�hp��շ�X;,�X��������w2�; xT��z�WS-4T������v�yV�;��r�~�#PI�q�VNhm��e�!�Xf��ݙ����D�EB�ЋZ)J@�;Ïɥ�k����@x7�Pqt�RU���X���_�?'A.Ϻ��Yn!�L���ė�W��&s,�dqf�B�6>T�q�U��N1y�c�d��2�r&t�ongBrC��6����P�t(�H*��ݡ��y��'�����#��i�`�M�Ac/�3����<�Kf�k!j��'I�V�e�I~���,��2H
��L�q?ì�Hh/jz(�g� ��A݄�d)9QyU`��ޮ�v/��8�NY��2X��U֠��U�l�2H��1�!Iw�=��	̘��K\��i?�$`�L�����B1 Q ����I�ڬ4n�/�	)>\;8�싶�1�N��3*�%�S�������a���E�D�Ym�7@��P�4v��}E��ˠ�����5<���˽˗jnX� ��<ð45e����e�l�r�Z���\E&%L+�|[���������X�2/�������x����|j��zS���g��5��u�x�K��d����yX�d�=��L١I�裆kf�f��7a���3���H�H^!DL��s^�^Jgv�Aʩ͉�ş��T_ñR��sj�)��Z՟�U{Iʽr��v�`Ƒ4bLv@�H$�߃���>����:��O.5*�g�I�6\�ut|��̯C�Nce�����a��,\)3*{ "B�i���E�w��S˦����`*T83:<B��0�%:��x`�7��юZp�&�ֵ�?Гk��L�����&׿�Y��Yu+[�aə�\ +\ݍOpR�+���zC?�8L�x�T4aŝ@XaswWp�n+��"�p*�H;$����� i!��3$��/|i0j�R�)1�<M�Ҷ�m;v��T���F�4���')/�k7:R�-fv����S��3{E����9�`�H����9�)^�� ����H�R�wa��<��mlJT�S���y�	��:%ד�����r�M�m{>ᔇ��9O�F�-*�����I��;�u�(�'_x �Li�m�6�9��F�k���������#w`,C���b	Z�>p��5o���:�*U#� T���Lײ
��*��H �����<g�K��M����
W��dv��S}���8�C�\��?�n�������̆�/乮7?բPd�m�b���z�hx�0���9����ڮ8�#�_p;��rcKF%������s�c�N�qn�;	w�r���s�w�(Fe����m�<�`^����@R��|�<��:���R�Q��"1��\^�c
M'���pm�>H��IJ����J�p��J��&9tT�U��A��JO'��خ�\u5���=�66�ri�񛅎Q&� ���*i�mlH�_=�;\����>H�C� M�"�j���fq�
7��q���M5��XX���p�V'�.�R.�4K��V����A�V]�g*�bb\�YZr<��Dv�q7&�x
R�b� �9��f����ӭ!�&ItZ�Xı��蕈n���0p��]�w�.Sc����)��d�d敐^:�5�V�ħ2��93���2�"�D���:��)�z���~:Z�6�TW!O.08ݮL�F��*�{RSe׾��`���Q<�TǾQ�+�p�r��Ɯ����!�^��u��g��n��)S9)�H���#(w�R��]��e���^�O����n�����OSO� �VQ,~󄛼�Ε9���Dɯ&����tI!Vr����]�/�x�Im�E��_��V����4��mG5�)
�5�F�v�^,��\x/7+T/��</V�����!�鹀n�����)sL�o�J	�b�jѤ}qx��[si��^&��НX��Z��TB�����_�6��}�S�u��2�a�j_�;�.1��l�i�Ģ�F��AyE!S�m�$a"	�:ҿ |�e�o*)�K�q0��#XR�"0B}�2B���oU��s쐀�_,I�R�
ha~��uSb7N�ܗD�>B�cw���Q�
DmC���w�1���ըaT1oGC^�#�IVr��0ܭ�O
�������Y?��h��淣x~Yt�@C�/����4ގ�9�t,�"�t��)�[ E}�"���g� `��߽�,�%�d���1�JkZ�nS����	!S�-K�1��@j\��K��Vh�-Q[����ř�I����L�L��`�:b�b�|��i��8v����!���J��H��"*�}�������y]%m��	��_�lB��.̊�^c�����m�o�7�D$���T#t�Ж���w��O�X���̇�z��Ͻ1/�����'����q��`��,EĄ�h�s��n�����.�h};t��]�f�nm�]�����}~P���G�k�Z��\{p�Z�+�r0���F���.���0dҿVϐS�Chj~�jq����ֹf��8F7�=���4�	GV5�o5�>�r�|�sxԟ>�VT�b�Ƒ����x4�{2��zJ[��~�#7�l[DD�����h4�@WRB���-��D�"��!���x$����uG'+�uT����@�.`�aM��}`E�k�
�-"��d��W��3�^��u<.@�vL���]7͓�i*-�x>����A�*�P6nw��=:�y�g�,�^H����tU�9�U��s�QD��'z���n<�ݪ/њ�FZ\#��:<�H��� 4�&F�A.P��v�j��fi�(Pba�<�b����R��E��\��ޏ[�s֏-�ǁ��Ο�oZ#��@�b*���I2K"O�J��MZ���O_}�P��(���6�>��� r��s��O���D�E��ܒ~!4������z�Ȥl�4�������5�V�(��m�ߊ3@��=
B����ߠZ��h�\Ud����U Q��~
�Y���؛�<K�������v@���}����Ԥ��y��ӚlpZ�jT���0�ē�ӷ�,'����@�f��{�xoT3z�-Z�������V���U�da#kc��NC�F���4=fx]�g��w	D5�Bw��Z�Y�I�dd�kúG�
x�3�P�)R�����9��PW.��ƴjh�m����W��&N�Sd�SY��"�>O*�q}V�	DΪ�9�2gϏthg�qEC���V�)P�d�(�VX*����|�Ly5�∫U�����}`Iv��\H/w�`b<Z"����� I��e����ֺA�N�
�D�L͊�?^�}C�2jmMo(��� ��qX^&�?2�QS��`�PީQv���8�ƫ�3^4��{B{�=ml7IO���!���=E�̳������D��$�^�n���n�B�T� ���!n�'鬒
��)y��8e�궥��N@ �끃nq��[���7���Dp�P�2���r���k����/�F񷺿s��p�x�w�`˒�i��~د�۰O͍��"�e݋��*N�M��=�&�L��>��[����}��vē�v�ǐ��i#�I�e�P|�m z�ɷ�B]��N���代F�/�����F��sY�ߑ=������>�Yf�H"�������3�B|�ù�^��W�!���#<v�N:�(6Y�ZwTz�?R^��j����4�w��L{!��J-��8``᫡b��P�U@�,B�7�l>�j�֕u�
|�E�g�67;Rt�M#�J^�N^�,�H��m,w�*���B`̴�"�wZ��S��F�W�`巍86:���텠��`��8i*�;�,cp|?��{�?K{z��LUjǤ��&ҎJY�qqu�Ԗ|zV�u����\mbO�+�]z��8�|�2R�0�xO-a�a�pA��T���.�H�����;���K��O�$��|ͷ�M+1�KcM���܈�&�=
�򝫁4�0'�6f2�R퇈11#�����{��s��9l�HR���4KI^r� x%ȓcݡ��ԾTO����Tm1n��
�	�mD%�Oɴ�Jز�Ik�H��d�����A��*Dǻ�b[��d!�¶��uv9�b�� k �h��6!@���k(���RA1�rt>�^��,�Ӧ�]����o/�s���鋊�̒���&�)�w�M�E�%A��n����Ә����B�M�����WR��Y�v�6W�dxГ��C�&���(�n�HO��WL>�񂁹	��]N[d�"�be*xz�з�?�+�s����	�ނ1pV8�r��%���5iд�N�Z�V�-����w*�;F@i���<7��2Y^�9�� t��O�<��:-��Ry���]����i�c�9�xUXp(��H��J�����^���Wè�U&4��]�9��U���O�P��m�\��/�`d61�ai?�m�I�A�0���*Dhl���_�]1;<T����Hzc h7�"&�_���.q)��)���l�,cFXyt�ˋ�'"���-��4�_-��ݓAf*]KHd�}Z���U�j�D�X�7�w�ybn�� �5:��I��U5����9I�+nX_��㡷n8�0+�&�xr�����ΰ�d��d�jd�gk�b�5U�P���P´���_4�	:�OP�iQ:��c�5�_Йޑҍ]G�/!=A0�q/�GR�F����<�{m� �9S4�;ã�I֥<+���L�s���g���}�����ԉ��$pA�}D�$V��#П?	�>�k���V]j�ғ��׆��C30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸�x�rhK9�1�#l����_�)��ToڬrN�'|W�Ds��&�M3�i��P�E�d�F��FB*�@�J�O~6�I覑�	ߓc?F�KE�ַ1�v#p*�8s,Z�9lTA�'8�qEx��ϦIq4hF�w��Ձ��Ýo�,�b��<YAΓ0u��YH�T~�M�&a�l�"����|ج��)(_�f�O�jE�x�`�07M�8-��I� dh�
`�irr�����A'璩
�q��ƲLZX���h[j"�@����� f����X�'ߢ9{�h�2(k�J
>�
]�t"�*m�}j���B�I�"��+�E;�%	�B�	�LR6����4k�4T�$i��oj�C�I�n�F���F- �ѱ��:^��C�Ɉ���R��!+1Xc�6Q/�C�I�Vs��k��'M*���f��a��C䉃D~L��R�4}^�Q�D]�r��B�	��p�Q��ǘV����)zC�E�V$=y=L��dȫ^BC�	%X0�p�E�
2b����	u{�����!Ih����bEy�B���kT6pՆ]h6@��?y��&%A�X,G*�\�r�i�u�`)p!� JfJ�)Y#�M3�̘Ix(с��<!��Q�S`<4$����_�xO^3�LƷ2��A��
}�I����:u�|��|2�Ac�` �y���obv��M�U�� �Ԡ"��� "O�h2�  �.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   y  /  D  U  '   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=��J�E�TM�P������PŌP_`��7ju�r�d�O���<�'�?!�Ov�%ʢ���)�-#�E��-�����L9B8��	�}xy�@�]��4���N�.ς]�
Z�>=��	�=9A�N^X$4��Z.��(��O���O��Ĩ<I���'�xQ���وnB���J�AoH-�	�'�<@D.L�s���#&��C6L�{��o�4�D�<��*Q�?���HQl4�p�c�h��m3���ԟ '�h��?a����'��3NԺ�ȷ���a�r)j˓T��z�)!��<��P�d%X���&k���ay"�J0�?y����L�t�U9l��H�#�T;���O��;�)��
�`¢ȃ$r*��&ɀz
\C�ɰ0r��m]�����ɣy����/���?��w�Ͽs�����@s!L��,N)�2d9iB�'�a}�	I @	��Bp��{�|�q�%-�y�n�	V�x�at��rq~]����yBB�
RYX�Y5M�~�T`��Ά�yr|J�!Y�k���T��-�p<�c剌��(Ѥ�^�@�����������H�O���' �	�z (PЩH��ɢ(�Zc���a&,O�$
�-ڼ1V�pU猤IV�u����B�ayR�BNj$����n ����ϻ%���OZ���_x��Y����Ml�L�VZ�{c�0�#��V:�P�ēEq^�*a��O�����KO���O�<Fz�O�r]�pc�A�,�̨B��;W��)�1��jm4���?y���?)N>��T���GN��fg�h]$S�E�'*!���><`D��E|B|�f]�p�&��OnTh@�Ƀ ���S��;��L�Q����bi,�Oڤ��E?:���Aץ>k\�s�"O�����E�"��ƀ5h��×����'���e���M����M�@$S���ī�턙ZPyç	hBY�|�Iܟ �'����bĜ�$!DѦ@{u�@��G�Z��1DG�=�2��,�=��E|ҍ��NƤI��ןa�N��A��>(Ҹ���1(n�Q'�X� �	�i2��O�����'�@7�O�6��<��3�! �kUPub$�R�?k  ���,��䟨��\�b��&Z���T+h#�8���;n��B��@���P�h\�>ϐ	��$��>�RE�OD�G=���i'>��'Q��C�I�*�P��N�9��te�'����}����;��)��G#�e�R��-��`�)���HOJ��3g]�DF�YS��)
xѮ�3�ޏ;M�Y�'O^��'v�P����?����?ɉ��DT�p>�M��m���4	߂��'A��'�������(fZ�`�ʊ�u����ǓY\Q��rQ�:������/:j4�����	˟(�ɶW�t��ޟh��ϟ,ק� X����z5�|� , E(5۱矖n"��XSZ���d���g� ��)bH�/MªL��ЫFⴳO��2�X|R�
F�,��*##*�S�v��	$D�Bm���(w����t�@����&�'� Y[������dp�Ȕ��X�������aQ�LH<I�+�E��,����O�p����K?	�K웖fg���|��'�B�O��A�)��mIR��1�T��Ek�0�&p�ڴ�?!��?A*O�)�O��$�U\��
�F�t�q�1�W�Q\��5#װPm����'��Q�p�L�N�<M�&�J0��uv��'	��(Q׍�-~b����ҫR�4�3퉼"��h��X���Gwȕ��H�O����ɦ���xy��'�O�1`�5xq��h��Ձ����"OB��1�P�	cl����M ^V�<B+TI�	��MS����?�p������TG%R���
4.��B�$��?�M>I�S��򤙻G�4Z�'�� �ؔD�8!��ik�=�P��R�qЉ'e�!�d��U$pS'b۱'�If�w�!�X�x�-˗�V�_V$S�GE�Rѡ�D9<	ra��8=��,*�g� 5�H}`���Ȯi��>m���H� ^�4��c�0#6�d	���6�?	�°>����Z?VУ�MrcM���y"N��@5%�! �8�<��IR�yr$�@匰hGN2�~X���Q��yr� }_0:P�H�.�.0X��p<�7�	��R���q1� �F�*pd6�IK��#<ͧ�?�����kP���!�4Ӳ%s$��15!�d� ��أ9�:���`A!�D]�A��e"�-�+���C��G5d`!�	-q]��G�(�#� ��l)!��N�k�^IK#���$Y�f��(�����?U2�	�2�Н�3`e!���$}b��]�B�'Rɧ�'U�0a���@�r�I %c�Qv����d�E`Y���@��$�@L���.���H�*v�=�B�O1���M2V]�2�Uej�a�fIX��5��s���u��bt���1�]�i�=��ɽ%2���'W��eP��W�a�Z�pI�f6���IB��"|�'C�\t씙�eٖH���'�����ٚ���.�?�
�'.�TK���9���J�(L/��LY	�'p���̩A��nB�<��z�'G*�b��)��e���D�	B���q�~�'��Tc��i�#@�H��$�#��5Sd��9D�<���x��I-� s0�Ǘ(xX�2c�#�C䉗'�Nu�1��>�(����I#i�C�	���a�s@`�@�	�y�2B䉏=l��S�H,M�X5��� Q����ĐB�'J&qHt�X���b
*�ƨ��'O^9���4��d�O���h�[�D?PL$Xz2.¸2��Bڀň��K��幒�����ȓA�XSX7`d�1&�Q9p�@цȓ�8��g��*�� �Ƽ	A��ȓ,:TE�����ּ��LBR��p�OXPFz��D��$�Dq�E�A')1�@�È��	<1����ɟ�&���Z(qCD�gg͹ F0+�"Ox�[�&��Xb�uc��'5��0"O��Ѯ�4�t�hO�Np�0"O����G�N&��&*@!Y�T�"O�l!�OTe���N�i�d)w�DK�'�4���o#���v�D#)�D�86�� m��6�'�'l��Y��Ɂ�U8v� ���pf���Ш:D�p@'��(,S��s�#�z����4D�x�B�ң9M�mI'��=w_l� �1D�(xrN�T򔄁1`�*g����a1�� F�/�F�����k\r$�M4=�Q��F�;ڧ�(��"!�
m�z}������)��'r�֧� ���D�һ`JN8a'BA@"z�h0"O1
b���.3��K7@2C0|��"Ob}S���#V;�xQuOþz(�ŉ�"O84�M�!�Ti�##
V�1��'x�<�d��r\2e�1���n�Cw�O|?e�Tp���$�'�rX��:��*��˟,7��Z'�;D�di�lN�9���݉|�T!�
<D����
�Bgn.�Nb4D'D�h�ю�q9�܀0�x���g&D�,����W2�<�" Z��`"�*7}"�?�S��-$�H�Q�ݟ@��x�� �13����O*$
���OL��&�����H�F��'A�R0Y����y���1a�8���O�ay@�yReS�6��1�D.�E� �胅ܽ�y�J�%��pv��=>�R���@W:�y�^�Rĩ�b��/�r|s4�W���'�@"?"@�ß�1�)o>D�`FgK\��4�W�?qN>��S����U�3(H�ID��-p��eƚ7�!�_�yfh���6t'���d�k�!��^�2�� bSd@�x����i��	�!�ЀIЀ��!"�����$�!����h��`h�`�# $:�`TnH �d����9y��>a��㇧Y���BK#
6��u���?�����>�!��E��ى�V�2��� K�<����J�`�b�� �_�<���Ɔ!U}�X�$X&.�MG��r���YB<m��S�u:�p�㉧�(O�h�w��/�<��T�=k@-�"�O���Q�i>9�Il�'Gx���SU���#a�4R��j�'+lx��MA4.�RԐ�@H����'x.ЊvΈ��t��G�K8���'�R��I�
E�H`��Õ?C%��
�'����#�� -M8|�3�!SU�5�N�������3��� ���v�����( )���X���?aN>%?�!�C�}�� �h�3}�*��c�,D�aP��+r ���LǪh$�@�I,D��І�]�_4� B�)�v��|F�)D��0�B�z��/�aX�A�-*D�p��۴�<�Ui\�O`H���'�<��OV\6�' Ƚ��`����4#�)��a��O��O���<�`ac`Tyag��P������h�<��+�B9� �:@ht(�d�<Aң��� 〮L�v�֫D_�<1��H�t�Ќ���ސ:�<����Z(<���߂IA�|z���,u�*��K�'{��>a�X�O�I���a��a��� ~�L��@�O(��?�OH)4H�31�E
ìL�Y�m2"Or`����0^O�Q��Z�G����"O�]tcA	+ :=q�B�z4aG"O���,�h��E����.�>X�`�'�\�<��H�pO �hD�%?��Չ�A?��G�\���T�'_�X��0�׽p���j�DD9TZ92�+D�8�1�� ��A d��1�N��0G/D�@a׬A�@�eQ@|��Dg8D�lp��^_��`�u_�sT�H�k6D����٧s:(�%�O�ya���d�4}��-�S�'dX��h�^vRT" ӑD���OYS��O ��"�����1[�B����z�jL�1N��y�*PW�ƁV�"x�l��j� �y����#��q6k>:j��ֳ�y��;xI��`�#A��&�Z���'�y�+H"	�-p4�˳s�8�����'��"?���П p��^e��P��'//D)ȑ��?iM>��S���D�8�ƙ�1�!����W!�� ��)�Da㨼i�)�:���%"O�@��M&\��a�H,c�Bm;"OR�P	�<!Ш-��F�
!�p
O:�4	Q˞L��� H��mL���O�+G�Ӄ$YH��F��I���t|�=@���?��xt�	��'r <
����Q�������U9�n�qTeF�BXm�ȓ�Ρ	H�~;� ��[�PtdE�ȓu��E�F�	8 q$��s4z���	��(O��8�+�/.rP��E��y�h(�O��jt�i>��	ߟ(�'�ݰ��Z����Sc��'|\xpQ�'����׏�?.���U��3lk�i�
�'��=��O�/2&iCa�+jRT��'v�d�Iڸ
���6��f�" 	�'��а2*�T@.��L�32��PHH�����	H<��X[.ƣI* R��v��8l��K��?IK>%?��2���b�@"�Zq�����!�Q?V�*��Di5�=���5<R!���8�q���Al!�h�+�
.8!���G�@�SÐ�#X4�7�!�Dݐ9=�Yw
ܡCZl�ْZ��qO<�F~b�Y��?I��ς`�#�
��b]5�_�d��|"����	�7jެ�1*��`����m� e��C�W8��䅞3���؃+[/��C�I0����č�'`���G�;m�bC�I9���S�U"hohY�Ձ�W�B�I�5q
�����f�\R��(T6a@����a�@�}��[�c�"��D;4��B�i�~�2�'a}�AR�*_�D�R��D���B4���y�G���)�O}��w�O��yB)�97%L�2
��E�%r����yr�N�>�t�s�F7;x��Uϒ�p<)��	=܌�A��M�F�z8�s %@2��Z��#<�'�?����$^4V	�eJ��DU#�H����F�!�dȻd�TM0���8V�:�0T!�D�G2l�`#��'F��1G�iO!��.P�0(��0@����s@!�	����	Nx�Ɛ���R*�E���?���$¶"�& Xׂ��6d�`*"}BA�L'r�'$ɧ�'^-��j&*
�|�h� LWEy��ȓODP(��ݢ%���l�,���7��yIg�H�"��S ��4Wu,�ȓC���8��[�(�# .\�ȓ<*��%���;T ��r�֓.:���=A��I1W��DK$S�hq����7Fx�{��0ZӴ��	S���"|�'ɸ�`��:a4�X���C
�A��'0dl �!ZB;>���*�`y�
�'� PåG����
oE<�	�'6�5{Qo�!#T%	�L�/1�,��'d���"�`��5�Ć䳢�~�'�����i��y^$������K�P�GA[E�L�	៸��I�\�2���I�$�u�%�T�#*VC�;?*��{C�[u��cj�L�C�	�o7�=af׾c�H��b �/ �C�I"�r$d�#^� � ��ś<����$No�'t&L����O� А�`Ќ{���+�'{B�ي�4�"�d�O��#�����5!e�|$)��bЂ9��Gd�����El�� F'�)^	�@��-l�e�1�8ErL�e�-����
�� ģ͔a�(�=_��ȓe"%(À��uI���A�&Ѐ̤Ol�Dz�����9����1��~�D�v����R����şp'���
HR���l�tl����r4�tB�"O���%�V<"\Y� ��B����"O� 0��&F����a/�5|$t�"O�Uqcg	/S��qU�[�hnD��"O\0+S/�&(�q�o�M^H����PY�'��ɋ�7m.ly�l��j��]��$Qc�ds��'��'��Y�t�W���q����!�zԩWb<D�Ԙ�mB�nҔ�.�EnJ��7%:D��� 
��C&��S�U�F�R�3D����Ҿeꄡ����2�4�iS� 7����<WԨe�?X�Q����'�'G�Rٶ��3�������yub�qT�'�"�'oƔ��ط/ �0�s��*� ��'�n��pG�4�"���0u�(���'B�,ȵO�sG���$C��s�<E��'�αK"�JY�Ҩ��K)r���(ǓT�Q�,�ӬW;M\k� ӯi��f��@�'gE���d�O��2�2W�@��� LN�g h �O&W�Ȥ���OD����Z�g≥U�N�)���72z5e�N�yGF�"��P
P���	P�'4�ф�)�3��^��+E擹f�n,["5*�p��I|~�$(�?�'�HO �� ٨V.H�7DE=\�h�U"Oޱ�C�G�ZU£��f�� ���>Qs�i>U�	d}���2n��+�k���K7	^4j��ᢟ�8�	�P&��O%f�!v�6��Ҏ��l���+��V� �rk
�p���'��T{�
��?f�%R��[1A}��y�
[(c���  Y�G{f�b��'����D�l*�	Jce�#�b��aD��?Q��hO�b�x�C��Z����G�)��c�"D��Цo�$# �ɗ$B�e��!`�"�	��M+���d16�lx�O웦��h�����_
	�H�C�铧 �����<����?1�O�~��d�ϣm��US��� 4x4Q��O
v�ؤ���jW̉c�=,O�� C<�b��A� ���9���4��r&�hWo蒥a),O��� �'��\�(�e�X��Yh��H�R�%��H؞��-]���)sCG^t��� $��;���A�����������䌛nnu��Xy�T�X��i�'�?�J~b�4S��<�5͐6
��aJ�X.�0�'���+ �J���w�p���-�O��K�Te�[�Q�d�ѷX�B��U�3�ēGނ!`�Tt:X�!Dƨ�(�:�(�R!7O�8�TꐺD|l�;$�xB��!�?)���h�X6m�-G$��.�g��8���QC!�d�vNr�� �ʏF"Ĺ�7Ŗ'�xR�<ʓSi^��R��5|���QV�R.!��}���u����Ob��S���D�'�R�'��I���%Q�L�Ę������B(��&�H�!��L�g�I�O�R1ۄc�W��X�v㖲y��$��.Q }Vt�3�|i���xr��o�t��O�#.�(hEn��N�\�$/?i����SS�'y\m� `:}���dށU�ؤ��'v��R��/KP�T���;a��XQM�,R��4�L��>��%S ~��:��Պ&S���gh
'{� ��n�:���Od�ĵ<a��?��OP�x�Gl
Wv"�S�lM�!(Ta҂뛚M�
 !�w�`k��'�԰q!�
?7���5CӊoJQId��#�vp��mR�	���'�pؘ�A�f�� V��<r�2
���?����hO�c�8"L�W�đ���[�>�*�p�?D�XY`��&��X��{�V��qO
@nşL�'�l�C �~��4-Xᑀ��=�z��N�/)V@�"�'��	��(���|rq�A0)� Ib��Ú"��$��B�ʃ�T4�^�q@���way��4\[�=Ѐ�V�GE,��3c}Q����+�,���ܑ	���$]�5q��'!�	�m@�d��l�*e� ��¤Zs�t�p��I�]���#h�3V2ൂF3�HC�	��Zܺ�I<G�ԅ���3���V���ܖ'����[ir�����M��@-.�舘�D���)@G\�z�b�'���)�j�/u}*���4�r�-�@����C_�Z�$����˥O�r�!��
戟��z�k޷i��ӱ����TŞx����?9��h�x7-Qd����Ÿ]��%�1�с3G!�dC(��XC��
1�b8	Ta�+D�x��6ʓp�Nl�_*bn�C	I6:�!��?A	�&�$�  @�?3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  8  �  )  )  4  ?  �I  U  W`  �j  �q  ~z  ��  ��  P�  ��  �  &�  ��  �  ��  �  j�  ��  �  I�  ��  ��  �  ��  ��  ��  � � � � '# �) n+  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�
��.B*�Z1�f��+%��O���$+$�T�J6)M3i�j�+�R!�dI(�$-��G�!P�Ȁ��ѻ*�!����UaƏ�R�2@1�O܅M�!򄕑[>J�!2��+��Dk�N��t�!���-<��A��@�uy�q�A�4�!��wI���E�9��%�k��!�,���A�k�^��Q��$#�S�OT�A���Af�Q���3�ր�
�'ؘ	Xa� �2]t��O�*�Qi
�'�\�9����,����6�D>y9
�'��a KI�}?�!��K��{%�ł	�'�P���]�fDD$P&K tsX��������>�࢓!&\0 J��]�:F��A"O���D�%5��xZGKC�& �lP�"O��c�p�bd�SK8sI���"O�a��HabV�+�'O�}]�a�a"OT��fj*6���l�EB�LK�"O�в�,1	��0�&L1y>�y "O6p�bE�jE��C'�b&��B"O�6� 6m�>�*�Ř�&vP�3"O��p�C*R�TJP@�P�LM�1"O��C1�T y�4��-��X��"O
�jQ�	�1����#��0g*���4|O� ��v��C��af����`�R�"O�Xk���f�Q���X��< �"O��a�Y`&���!O+v���"O��``J8.D����� š"OҐkqOL�y��O3yҬ�8�R�L�o�n1��C�<4½ÖdWv�yD}��M	�i��h�����a�*(�DB�I�<���G�7Zʣ��@�"=ɉ�T?Q�-Z��|�)���!F́P�=D�@�'J� rl�Zg�RUZ��4�p<����v���� O�[1c!��fn�0$��&>-���	Qx��/C�Pnp�R�BP��y��Jo�$���E< bQY�R��~���ӟ��>���۱ ��V�_�nhK�Ig�<Qm��	j�X���ߺM���R3��xy"�i?�⟢|z�!p��烑S� Ӳ�X�<���{�&��'F�f�J���J��=q`�DHJ[tOǵt����LI���hO�'y��Mh�F�X��|�`�G=q�	��|�&���5^�,�
d�I!�������s����`�)�z�PTG���
�R�d�}h<)Ħ�d<�ؘ��Ss���o�o�,G{�k�:���f�S���(��ˍ�yRH�Z;�1���O�x	�����y"A͇Y�(�1׮��t�>e��8�y¬J�;�[4��~�*��֟�yr�ϲb��#�\'o��A�b8�Py�M�^<�a'V�H�����-b�<9SI�6���ش�[(���X`��b�<�v�R�A6PP�7�$^�4͐�`�I�<�7�7'3|\� j�j�ج�ѯN�<A�*�f�42B��Z�� E�I�<��d�#L��@�É5�t��B�{�<y�l����C��T�0���"@�v�<��!ٽx������;a�$��tfJ�<ya��������6N�&��e�E�<��
|L��)�샴���
fA�<�GDޠU�>52��X2{��тvk�R�<p��.[��@U�,C�ɢ��XO�<�
�)��m{O�V�`J��Ee�<)5��$��` 4f��&���r��G`�<I�DŴ^%Z�㧖�i�d�Ä�]�<AQ��O[�qre`W<n=D%R�(�p�<a4D�x���V��A��Q��FC�<�@J<(�Rł.�𢴣�c�<�1�Ð�ZDa���:!	 �zgjYU�<����`/��%l¹!�0ZrC�X�<9�EH�K.����`D�"sz�Q��Y�<9
ԃ,�4���%��3k�(H7��S�<�⩉�4F-��T�`���+!�E�<�'�.v~�I���K�)X����ƈz�<I�e�l�����g�
��P��w�<G���f7�t13��t�rXZ�`z�<!�	02���HU�<
��!���x�<���H��a'H�F���9w.�n�<���RC�M�E�a��!�Ke�<i�/V�R@��@�ßP��A5f�W�<qg!]�On�qɅ˗ca|h�n�<)Q�H
�@q�v��͐7*g�<Q`�)iub�;.-��!�m�<q�&qP�!pC��*є��j�<��	R�|�������8�fEx �^�<�n	T}�+��n��R��W�<�2kT�fZ@�V���6eR�T\�<� �A�f�#y�E��K���p��"O�pA ��T��Eӣ*DG�ԉ*2"O�h��4X�a"+�38�li"O�2��Z�b��4���5"���"OVMK%cޭM�t��b�ͬ�����'n��'O"�'���'���'�"�'`�|A"ʓ0H`��c1j�x���6�'���'���'���' R�'���'�D<��GٛY
F%H�HVW�4�2"�'@2�'�R�'�R�'<��'���'Nx�� �����Y��ӛ$[rظU�'��'���'�'�B�'Q��'��ԫ�i��
6�Ɩ4D��Q��?���?����?1���?���?9���?a�F�k�����
��(oܕ�M_��?����?���?���?9���?I���?���l/p	xa��;I�C��.�?��?����?����?����?i���?�)�+C��!GX
+��lj���)�?i���?���?���?���?����?� F
.K�t�9Q
65�T��M�?I��?����?I��?���?���?9C�D'P5U��'�*Ϡ���E��?����?y��?��?a��?����?��*��@��}�ǧX�*g�Țí���?����?q��?����?1���?����?���B�X�ka[6�
�;�D�?q��?���?����?���?i��?�LL�p8)XF��9��@���?���?����?i���?��\8���'"i�� v��`S.��2����h����?�,O1���>�MB��_S��Ô�W$]��y�H@�<�-O�qn�x�U�����x�3�A;;���A5�C.p�ah� �����3��nZl~B?�V���m���!	֦�� ��(]�g�J�{'1O*��<�����2w�E��� _���"��#<�<��'��I㟈��6��y���l�ܭS��E9T���Q� /Mz��'��D�>�|�e����M3�'T����t=����D;�򽹟'���_ꟴc��i>U�ɘOX�|�N�%�>Б�'�:.�r�GyR�|��1��ܟt�s��3����́�UT0�T� ���џ����<I�O
��"�
9ZRr��e�t��֙���	#:"9�,4��:,���[1G�K�ĥKE#��hcٱ��~y�^���)��<!��G ���×F��~L<��6�yt�"�>�/OD\���w��iK��6Ѷ̨��	�o�L*�'��'��L� ��V��ϧ���-ɾ4�zq9�E3��q��F�u�t�'�x�����'���'O��'��H��@SԈ��)�*V��tr4\��ѪOv��?�J~��I��a�,aCh�HS���j���؟$�?�|z@gK��,:�c��&NR�h�/�*T�fIP�έ���K�L)���:�L�OD��ƅ�R�V56�Z���W'�N���	��d�O<���H#��D�u�_k~�a)��O n�[�$��	ߟ\��ǟ�9H[�L2�X�ւ$F��������v-oZT~"J��p�'�䧲�/�NݙrT�sX�1���&/`q���?�Uh9$#����fZ��X�Q���?Q��?�Y����p$����+֚	��9��U3]ZH��4�IK�Iß��i>��D�]ǦI�u'.*Tsя?{rVI�IB23�4�R��'�x�&��'��O�H��ɱx�ne㕌8C��ٺ"�	:��D�Oh��O�˧voD9�GP�VY��""5�t��'���?i���S�T���"����۷Nc���B�Z�5���*b��6$�j�<�'�@��X�I�Q�]�叒a2Q�1�	@��B�	��M�V��# h=Q�@$*��9���_�<���?� �i��O�<�'��NƆ���RU�l$�L���*���' �K�i��	�ip��HUҟ��u������5�F��L:Z��1���$,|O ��%2Hn��s�j���9U%�l}2�'p��'��l�mzީ)�A�aJ�K*�
#s�q�������Iq�)�S�N�"Em��<�Q��{��� v��Ds*��+�<���h�&��u�	uyb]�@H��̇`9>� �*Ka��Ͱ��<O\��'�'��d��4�	�td ��c\1��O��'M��'f�'�� 	R��@�u���Q�f���.?	b�V�u#�݊�4&��O�D���?1fHZ�hӼ<���6k�zL�4bʆ�?���?����?����O ۧ�Ԑ]�D%�U�C��a�O$��'R�'֖7�2�i��%�فz��D�1 ۀ��S��d��I��,����`s����p�b�?��A'
����&��Yo�th���z�IKy�O��'��'�2
x����2��	a�T� A�-������O����O����YQ�n����Ӱ^�,���!P�1�'b�'�ɧ�O��������\�& kQ�	�9�|��Ћ��v!�V�����,B�n��d7�D�<1��B�S��t����grȬ"����?i��?����?�'��P}R�'��!Z2�1&�6=��ڥ�ESC�'��7-6�	���D�O���O
L�&C��Z�`���$W�d3�����L10}v7�3?����.R��|:�{�? ���jӽu��y�"(�$��15O4���O���OR��O��?a���D��saٶL2�$�ǟ������K�O0ʓY#���|2�U�h޲�Bp�P/]-P�����+��'��T�e�ߦ�'X}�F�	X�h��I�;h�����Z#h����j��'��i��'IR�'g��)sf͓7��)�gE�(>���'L�Z�<�O����O��d�|*����"��T�S�l(��I��f�{�I��?�O[�Qsl��Z"4p��I��2����0'$���CC@�i>����'|$$���F:6��� Qi:D�� �ٟD�I�l���b>��'G�6-N7 O������H��T��Jĺx,��O��D ֦��?!RU���I�O���:&
*O�R�ʕ��9-2��	쟴9�o���'�����Sbr-O��h�nE�v��
؀|�����'��I�L��ǟ����l�IB�EѮ��� uF��M�(B���0Z`t등?���?�J~���l���w�晊�lF�5� ƹp;���'O�O1���ؖ)i�J�	�v1䔳�f�@����B��xC�:O�������?T*&�$�<����?�©E�&��!fb['\��������?���?y���d�L}��'���'@��sfa��5t��%�����DT^}b�'l��|b��p��H��_�|���q������ݿJ�F�k� |Ә�&?�P��O��$ѣR�ʐb��4Ա��#,����O��$�O��D2ڧ�?��	�"�,l�"��7<<J���B��?��[���	ş���4���yG�0P%�T�T(J�O�paBGE<�yR�'R�'*��KV�i��i�	��?)uf�>T���0�Jy���a�� N.�'{��˟����(���x�I�n/�M��Ǉ�72��k�aF�Q��'������O^�?���9 ���$g�M�@�����O��b>��mB�q+!3���6f�>$ e����`y��Ud$��
\��'b�	5)�\I�qI�)LS�0��>w�A�	؟D�	�8�i>M�'����?i���o�*��g�Ƙzf�}�eL���?�ĺi��O���'���'���<Q��\��2�(���D�'Rp8ǸiK�I�I�Dqb�Oq����X�*-�3-��Z8@�Z��"���O2��On��O��$=��%OL��2����Z,�v��8��Q���(�����Ĳ<"�i:�'����@�;o`���#J�J�Asך|��'��O�}ôi#�ɪk��(zP� +S��(���Lm�x��LV'��L�gy�O(��'�"`ŒQ�l�R/�y���r�Y"r�'������O��D�O\ʧR�A�.ǽ>��v�/��'if��?����S�T�̂;��U8�"E�����Q�*e�ʔ��*� o_������~�|��0q0�2E�¡;&1����-��'S��'����Q�jش��C(��
�`#c�S9�<��?��?��čL}��'=��n?�2�y�o�<&�����'�B�� ���������?g���<I�	�Lt����sN� y0@�<�,O���O����Ob��OTʧ]�����t��ܸ�B�K���Q�[���I��t��l�s�@k����q�	�%
r�1��l� ̣֠�0�?Y�����ʹy��?O���H*`�x)K�G��8Ͷu4O���W�2�?��L2�Ķ<����?��E�=�\������imnQ�SGF�?��?Y����D�y}�X��	9�APm�PMpT( 	$��?R� ��ߟ\$��#��G�T��Fr�8���-?� ��z��ɔ���'r �����?y`�ݺi<�铰��H'h���K�'�?q���?i��?���)�Ol���cC�=�ijw��'?2���F�O^t�'5�	<�MS��w�2h��KQ=S�N���דz(ٚ'���':��).�期���!��JE�M�F7n0P�B�2z��+�F2p-xX$�����D�'_b�'���')Z�$�>���X��w ��1Q� �O���?����I�����$f���������?1����Ş= �i�Ȝ��  ���^
q`���Ab����'�*�Q�.���a�|�^�$�\�-�ܐ������Jj���?���?Y��|�-O8��'
�βa�
M�t&�E�\`�"��q���,*�O����O��d�)4F������T�<ݨ���'n:r@��o�(�g���cj-ʧ���,�d��A3�G���fI�<����?����?���?���$��4q��YB�I�a!�49R*� a���'����>ͧ�?15�i�'��t#G�/cj���.U60�����|��'��O."�i��	�6��]�iD	)41�Ǩ�=���� q���8�d�<!���?)��?1�%ˣU�c�E�Y5j(9�+���?�����Ēc}��'P��'��3�^��IM*���9,H�"���3Y�I��0��Z�)����-6���	ceöS�����T:������M;�O�	�/�~��|�m�'zj�0ipm�b���]�e�r�'�r�'����Q��[޴:� �H"o�:Zv��K�%k<A�����E�?��[���I�D��u��Չ'q�ҥ�C���I��D)㦉�'�0�@��I�?���� �!9C��$G���r�]|xFM�S?O�ʓ�?���?	��?I�����g�h7� � ��@���}�'��'�����'�6=�rl�N�jcL���-b��y�#�Od��%��)�bm�6-`�H�Qh�3;��ǉ�~� q;%�j��1�@=p�BPw�I}y�O���	`B���F_�Nb������'�"�'B�'C�ɀ����O��D�O~��E���IBoY&^�Z����7��:��D�O��$9��Z�a�`u *�&� �t, ��^R5+�! Fx&?�BE�'F\�I,V�����f�k��qaK[�s�X���ߟT��ԟ�	i�O��]�OP�=i�C�Ke��ɶ�]"�>���?�"�ia�O��B5K�+�о4�}��k��'��'��'Qc���4��AׁB����Xrct��s�*LHA�� n;.�O&��?����?����?����Ε�]|!5.�pe��/Fy↲>����?����䧌?���7��@!vH�*�o>6�	�p�I[�)�Ӝ)WI�l�<AR|���+#&Ybdޝ$�~�WF$�"D�O���O>�*O��fg|=Z�ӗO�M�B��OF�$�O����O�i�<9�U�@�Ƀ)q�H(���4��r5f�9�5���M3����>����� O�>�H�ρ/7��sKU�ĉ�Ԫuӄ�58�`��3J~��;�E"s,������V�z=:��o���	��L�I�$��՟$���e &́@S�Qk�|� �]��?1��?q7[�P�'.�7�<�D!Z����$%RZ4��I�'&��O��D�O�I�7#�7�-?�B���^�;�ሥ^U��*k���i���'�D�'���'���'_�pCA֫<��D�G�ƹNk꼹��'=�[�h)�O~��O0��|��ÚL�r�ZsjԷGp�M"�[@~�B�>!���?�L>�O.�i0�ʂA�Nm���GJ�T��"�#@����T���4�� 	��-��O���ƒ�VH�͐fmT-P-B(Ј�O^���O���O1��˓{t���P>&�VH��-A^P$ze���<A*O�Mm�j��D^��ӟTQq�ɊZ�	QЯ�9q�hKmy��Z'xқV�����O��� Ey��[q��y��
X�5	|�p����y�X� �	�� �	�h��ğ4�O��\:�d�F�k7%^)�zARc��S}"�'��'���y��s���+�"4���>#9Rq�͖;B�n�$�Ot�O1��� 
p�R�I�F��p� .,�$�gf�G$�I7Xp�*��'lv�%�������'c�\��
�x&JH�C,_��h�S�'��'��X�<èO���O����;$ց	6#Z9LEȥ��3[G⟤	�O��$�O��OX}��F�K��Ġ�C"y�z�����l�A$G�'c:)J��&��>'f"�F��G-A��c�� @fٲ�&��<�	�p����dG��w���̶t�	�u�W6�tK �'��ꓑ?���/��4�L�DꐐqheɃ	�@4���q0O���<�vJ���M��O���E#����DjBxQ����R [�^dۓ�r��OTʓ�?	��?	���?���?�ֱ�ĥ�eMҬ��)��R����*O���'���'����'Ǡ�H��+F@j��I9L\>0X��>1���?�J>�|�BJ/��ɘ[�w����/��I�����C~��_�K�����>2�'���6���BC��2{I(Tv�ѝȤ������ǟ�i>͗'.�듇?��_�N����tk�1�$��
3�?�F�i��O,%�'�"S�hR��J&E�IL<��,���#~�6�n�O~�`��&��0��$�O��cA�D�ac���&�h����	�y��'f��'&�'��	O?b��ڱeg=ة�vd�:u��d�O~��F}�W���ش��!��Ts�g� C��P�P|[�8J>Q��?ͧ8�(��4��$H=��tcBޒ$Mpb��Q�Ufґ����?�$'�d�<ͧ�?����?��i��/�\9S��W,|(J5��H�)�?����ĝo}"�'�2�'��S��<kn�m5&�C���0��$��	ߟ���q�)���?@�B��4
�A�6}�����A�.�Mc�O�)҇�~��|��L]�e���9�T�P��"�'���'_��t]�hs޴x ��HCnR�>��%eLt�l�Γ�?I��x_����T}�'�P�`��oc���-	�2�	u�'�B��Ƒ�֝�ow������	�u(9o��r��h2�a\�$>�ry��'i��'���'�RS>���I8.Z�aD���?����Q�����O����OP�?�������V;�\#�l�,���"�M�?����S�'*���۴�y��̃�:l��IB��U�ժC�yb�æu��������O���RT�V��S��R�  `��K6�j���O����O��g��	П��	��P���f�|�Y�ܪb��l��}�����៤�Ij�	7q)����IW $�
�UON�r�AH^��]'���L~�E�O����<bޡ��'̡D�2$�ナo������?Y��?����h���$�Dh���T���i$mZ @����$�S}�'rbiӈ���I��9�#��Z���"�(ߨ�p�	ß8����e!�1�'�Ȅ��ʀv� ��T�O�W*�q �T�P���0	,���<�'�?A���?q���?1R�֚΄͠�fF[��y���DV}�'w�'�Ou�����ȝ��N���XqW�W�5-���?I����S�'Z�\qD��s����b,ř	GRq�hN��M{�O$9ĭ_ �~r�|�_���pdӊ'����N��<"Θ1��ܟ8��̟H��՟�S^y2"�>)�w�XQ2Ќɫ/��<`��^�A��0K��%�����As}��'�'䄰'M2F�>y`���T� e�t,�f2���\�t���9"Q>q�%K�B�)G� ��y���N�H���	����	���������G�'���.�&��U8r��o������?9�>��i>��	�M�K>��#ʸ�.M���P��S���䓐?Q��|��II��Mc�O�n�8��95�V�T�Z|Җ� 9p\�l��A�Oz� O>�(O��d�O����Od�r�L�F�BF�ߏvd�yX�&�OV���<��R������	x��)��4�4<�Q���:�$|�A ���d|}Z�M����S�D�M��5{% �v�r��ʎu�@��Th$X)�����#���=��V<� ��޾��lHQB��R���O��$�O���ɫ<1T�i�� nܛ/�"�����^�*�'��ɖ�MS����>��{\�!S�F��A�f�߬NK�����?y2���M{�O����"�>��O?m;����{Ep�)mN3y��`a��'�"�'�R�'e��'��ӑ-��B��3%�%BrL��at�Y�O����O���)���OX8oz���k��\E7O:�ĀJtL�P��D�)擙	n�l��<��"N!�y��A��z{�1	���<�"�'S��$����$�O��d�
9G���D�k�~u`U�'K���$�O��d�O|���	����ޟ���BH9t�\es�J�,D���0CjJ��:k�Iџ���n�I�z�$Ec�m�%{����#kK3�K���S��E(��|�,�O<����?�p����I�R$�3)�<|.%��?!���?��h���Q����#�I��0Q��e�Շ�O�p�'_剻�M{��w
�y�N�d�>@)�ݤk_���'K�'��� !W@�6���Bw�d+������h�X$̞� MƘ��'�����$�'~�'t��'�V��A+� >�
y�5FO(B�d8p[���O����Op��6��@�^�2A	�#fv'�	�.�ic�Ox�$�OL�O1�F����_5}�d����(\�*}:�J!*�j7m�~yB�Ӊ@A�������$.|���d��kuD�!ܖ���OL���OF�4�˓��Iޟ��$	�(	D\1B�
-� �@�!���4��'���?���?A1㏘)�d�Ǐ;C�u+EA<2��ش���5$�x���O��O.�DkU� ���f�ѱF��,�yB�'��'���'��I�8J�����C�:�k<R�r�d�Oh���]}�OI�}�X�O�XI���`��!�h��/�d��)�d�O��4�>���q�b�"V�|�D��.�ޱh*�S����g$S�L�v������4����O��9["D�c�-W�Hp��B����O˓S,��֟$���|�O�8�x�[i����"_ dtZ�O���'�b��?9ѧ��$VD;��>� w�}<h��E��D����$�Rџ��|b@FQ��C3�y:�R@bQ))>����O8�$�O0��)�<�!�i[�}�%MT�'����j��Z�ZA�'���'�|6�3�ɪ��d�O�LH����\I1ϛ�a�Y�˶<���V��M��O>И`HJ�2& �<��$C�?����;t,�z�l�<�+O����O"���O�D�O�˧; ���-�Y|�CQ-�$Њ�2S����ʟ��	_�'3ݛ�w��`QO���16j)Ex�m�E�'p�O1���{�ja� �
=rh|"���\�� ��:!���'��tٵ�'���&�p�'���'w0�����4,�� �K�4u�-���'�"�'��U����OT�$�O���
XnYc���h�&�P��O�,������O.���O"�OJ�i�_9.�R��jA&P��۔���Z�&T�rt�#�B[��ss��ɟ�w΅�*�5��@��وXg*��'���'�S����d,�=�z5��Ѓ����p\ɟ|X�Oʓ7��V�4��e	Qn�� 0PT*������<OV��O����(�F7-;?�����;�j�iE9[*`K�"�ci�p
�-�1U��M>)O���O����O��O�3�#�<q�����*�����<�6T�(��ߟ��	{�ߟ�� .
�?kؕ
	���@������O���,��i(TF�Sѥ.�`�;�Q�4�1GMn���DA<��4���p%�T�'�r���] ?���ڋVq�my��'p2�'+�����V�h �Op���"cwЙ�G��o��P�j�9#�d���?)gZ� ��ԟp�I @|h�H7�ͯ��aZ¥� `�V%��E�'���`PA��?�is��4�w�Vq	��9�2u�N5���!�'�B�'���'��'��~8) �7zv��p#`�h��qk�<A�w,�)*5�i��'#�8�I3QZ�ig�C�.�
M��yb�'N�	%7V<lZt~"�
>߀ �C`�K$`ÎԔ[��-`RiA.�?�d+�ġ<����?����?	S+�$���0լ�<? ��3�@�?q����N}��'�"�''哱T<�A�ɖg�н �[����$��I����I[�)
�f[-ٖ��0�.Y�\��3)�1l�rC�#C�����Vǟ8#4�|Bd�&B����፻?	А� Y4&_��'��'3��Q��Y�4):�:1�X�+)8ȁ'oԳC1����?���^��F�d�|}"�'/�d�ˇ�^�萢�7.l�)��'�r��O�&����A�׭9q��i�f�X�|�Q��[,��d1O�˓�?����?Q���?�����ا#W@�����7?	03�C]�u���'��'�Ҝ���'�p6=�2��`%�H��d�P�F��Q(�OB�D!��IM^�6-w��(q"׮>>P���,�4A�(p��� U�z�I�Q�	Jy�O~bJ�/�Tq�$hJ�T��A1F��B�'��'d�I9��D�O��D�O����3Ŝ����K �&�,��3���O\��5�dT����"L�4
�M���ù*��	< 9����s_�c>���'U�i�	B�}��C56A�����X[���	͟���Ɵ$��Y�OHRL
=ͰQ�
"J�1eʗ\���>�(O}m�Ӽ붂;J٘A�ʍ�]-���'��<���?��]�xP)�4���Wn�H���'�Fh�%�� d�踶�*Hj��dO$���<�'�?��?���?��eˍh�X%I���F��놻��Cz}�S�h�IK��/"X��sК� �i��8��R���	韸$�b>��W��r���R���j�K�@ԅJղ�nZq~�.�	Q(Y������$C>N�	�p�[�F1���2g��?K
��O����O>�4��˓?��Iǟ����+0�z1ZF͉ou��c�g��k�4��'����?Y)O��[�f^>���hխU�~Ota�Y��耹i���.,�!Q��Oy��&?��*^I��5"�7<�f����2����	۟,��������O�(!ٗl^�qJpI�$�*
L����'��'%���|b���6�|B
�9c�(�C
W�L�bl(�C��v��'�����Ԭ���V���B���k�.T�gٯ_G%	R#I�=}�)���O|�O��|���?��?>�=
A�T�5���QtBZaĊ���?!*O
E�'=����O�*�ÎO ̆��͛!����O9�'�2�'�ɧ���k�uA�9RX�]0Q�O�@�Lm0$-ǒN^ܙsE���S
%�B��|���Bt�D�2����"����	����ǟ��)�SNy��g�llC7n�-���ѡ�ék�V�p�1O|�$�O��n�h����՟�F)�)G�P�+��uT��BL�ȟ������l�P~B�Q-T�H����$�z9��3$J3O��|��h����<I���?���?y���?�/������� =j�u��Gr.�ծA}�'2��'��O1�}��.�:a��% �?E��V���o�B���OēO1�Ę3�D{���	�jHu��65���Ù�v`�	�;�8[��O.�O���?���G��$DLݟ8���a�@��jB9���?i���?)O.��'�"�'���	�F<�;R�:|@�9�A(]��O:�'�R�$�)�Z��w柧V4R*�"Q�g���?O�hhRF통Z�6�&?IB�'�6��ɉr7�ybM�y�L|��I�@�����������O�O$"F�IN������X0@쒢sirG�>����?!q�i�O�NT�Gd<�A�J	����E*\����Odʓ|$VȻ�4��d�*d]H���'Edd�d��*;�~��Fυ%\r�*�i/��<����?���?����?�f.�	s��-��)�5J&"(Q�Q���DUk}��'���'��O�rh��,����\�H������>�l듿?1���Ş1�a3&D�\�t��㏪'*\�� �Q6cV��/O���s���?	Q7�D�<�boܡE]���GY�e��5�Uπ��?����?���?�'��D�{}��'k��*�h�^ݻ�B��8����'�h6M7�������O�ʓ��y�,ǣ^�lU"k�2_��5�Ԏ̥�M��O~-��,B����>�	��`a�"-�%SoĐ /g�D��2O`���O����O���O��?�y�Ï(lJxc�/�O}6%�!'Eݟ��I��x�O�i�O0�lZA�	R�PP�A$�0 �6�����*%����̟�ӧn�I~҄�((��Ę�lHHp�n�9D�t��@�IFy�Of�'H".^,_�xs���@�H�M�'��'��:��D�O���O�˧3Y4��1+T�s!rPW*�3q})�'�X��?9���S�ďU7��j�i��:�f�A{��!Q�
F.N�F���O�iW�?��2�_!�e�:/^�z�+h�2��O��$�O~��i�<	ķiD�u���6x:dAB��h�<Q��'��	��M���B�>!��Th��j�}hr����.#K�|J*O`���b��*�z�������r(O�
�/�k���C�'�5��h�9On��?���?���?q���מG�~%�A�
ܸh5�_	e-�'����&?��	.�M�;0ذ-4�ǸoF��3�%S�����?�N>�|��%�M˞�� �����-�f��0葵�&tr�3O�p��?iQH"���<ͧ�?eB��qD���@��"Y���פ�
�?A��?�����$]}��'�R�'Q��PB�O8@t�c�&�d�IA���o}B�'��O\�Y��W���&�5�f�jb��4�EO@�FH�Q+�D�Y�S�GM�D�˟P��"+\��,�=C��V�M����O����O���1ڧ�?�w�J�>�0�\2ܭ�G�����������<饴iL�O��0f��h`�X�rq�e��W�*O��OH���O(
Dm���gP���#Ꟍ-��C�$p��@GS�/`�q���䓬�4����O&���O.�䌘&������}_N�#t��	 N��sg�Iiy��'��OG⡘�,�Z�bN��.P�1��'��!X���?����ŞV�0r�~�ء�钗x�&%�gƃ"g�@�'�Jb�Ɵ�П|"_�@hდ4I����M�Q���r�'NΟD��՟�����SyRh�>���'q��r�����T��owF<q�"���D }��'���'���Q&�B*��k�/ǖu]<5�Ξ`��摟p��lF���'��@�8�2�&�"Fd��)R.	����Ǖ;=sj\�����?�zU2���BL$Isr$�(Z!�Z#*U �� ��Ő1+�<�2K�	A�L-�CE�$��a��0��~�$̢<#N�0aT*�(�#�7 ���H�aW/n�.�@�HŠ�::�����Q"+6EB񈖏^B�C�L� @ƕ#�%N3%b�C�Й�ԁ%m_�j��D�b�4~�X-�q�GB��HW+K91Z��vח�Dt��oZ	Y�h,R��>j|(X��۞:q`�%��6-���'�B�'0Bʥ>Q.Ob�䰟 `C�$%���I���	WonE�"��c�%�`�I۟X�I�w`iP����>�xy����9�ߴ�?�����d�O6���O��Ok,Q�&�$��6ђZ�bU�ӡ�'O��Ec���	^y��'s2�'y�'�l��$�Q5��P�[�Z�@�nZEy��'��'5�'��'N6�A�U7�P�C�T�DArț ��12��'q��'���4ן(}���S�M^� �4i�0:!��×�i���'B�|��'�l��D\9'*������YU��`'N��Y��	������*L|�-�l�d�
yP�	 1K+qސ�9���)1n�qm�ݟ(&����ݟ|�u�TS���I�ƙfZ�t���&g�5mɟ�ISy"�'��ꧤ?���?yR�C,z���T��$X�كs�S�NK�'H�'����'��'��	R"X>Tg� K="ȓg�Y)B�[�����P�I���ɟp��5�@�:o���B�L��pX�Ƀ��M[��?��@�����O��c@ F+���cl�4,o�I�ش�?���?����?Y���D�O��DBz��A�5Ō��Lh(lw֜��?E�D�'!X���Ã�Z���b���*Dl���M{�:�d�O���O,d�'��I۟��{�TX!��N6�Q7��(��qnK�I�lb��L|Z���?���V�[��+r  � �G=eR����i�B�'�����OV�Ok��"U ��C�Ѻ3<�:wnۧ8i�I- $��$�h�	�����y�� %x<yc���$~1l*�C�7ě&h�>�/O��$4���O��d�8s �t��X�T|pA#�4U�<��� �$�O����O쒟1̧<��`��N'ڈD�Db�a�˓�?�I>���?�A�B��~��ܴx�`�$6U#�&R��d�Or�$�O��&>�騟���Q�5%lm�q�Z�Y�@pp��1�8�m�͟�'�t��͟�z�o�Iܓ'�^�z�� 7��  R�S7G�2mm��4��Vy��'GV�>�d�Ok� _G�%�C/[�pqsW��.S�'���ן@��T�s���
F�zP��9�Jb��{Ml6m�<��f��&Ŧ~"��?!ᛟ��G�Z{ry�3��):l�*C�f����?���76�OP��M����8,e�4�oM'Zܬ���G�˦���)�M���?��?qҔx��*�)��9jX�i֝^��L`$�i���'Z|ʟ�I1H��5��N���*I�lȑߴ�?�*O��d�<�O��*h����Pv����[��h��cP��O���~����~r���h�����(8$�#�C��M���?Y+OFU�Oi�O�5����m��V���B&?�d�'�4 r�3�	����'��d
7rczġu��"\@�#�I�V^���	ޟ��?���~Ri�v�m��$�(w~���R���M� �\��?Y)OD˓���
1A�xiFw?HJw�ك�M���?���'!�	<MU�6��?�����֨�T��\.�')RR���'�ş�A �U�q9�cƨ�9��m��B���Mc�"�'��	�FfO��{0O	~
�T	��W/7��=9��i?"\���'������9��$�@���<�`E;�k.��O���<��Fx��u�өC�
(i�ޏ%��Ad�V��M3-Oz���mڮ�����ON��p�_�v6d<�[�|C��GXh�f�'7��'��	-�9OR��i@4΀�N�6Z�T	~r��7$�>A���?!��?����?�3�#T�v�x`���\�k��*���D��b>���T����ЂY-g�J<�a%�O�x�A�4�?����?A��Ik�����'���#� n�J3(��\���O>��!h��iD��'!�� ��9OD���O��� �F�9@������ *��5m蟰�	&���|j��?�-OD��!C΁C$����ݰe θ9Nͦ��'��T�,�����ISyZc"R��do�������3��\i�"e�.a�'��	ӟ�'�b�'MR͎6;�Ց�c��_DLk�k �z�\0�'1���<��ß��'�"Ih>��
�$9d4  5|w�HD�z�D˓�?!+OF��O��$F�#��$�o���0�M����ȵ�G6C���n��X�	��8�I_y�O-^ꧺ?�1"8�q� ��B��W�XSAbxnZߟ��'��'|���y�\��y���#DFm�&�ܳ�Ƙx�ʘ�M+��?q.O���Q�d�''��'Ǝp�D�^�"���Y�eV&�LL�5j�>a��?!��HJ �����/G�,i@���$QeH�VjK��M,OT����	� ���@�O�N���t�B�?8��m�L?���'s�� �y��~���OY�-�t�O�|���+)NL���4�?ib�i}B�'&"�'�J���d�q��)���M�bH>���J�Qt�lڋv=P�ǟ�'��z�䖲l���1F��#��hX�A3G��l�����Пh�������<����~b ;�f=�ᮏ6x��d�чE����<	wER~�O�b�'��s��� �̷.�ܥ Ɛ4V.<7M�OV�DF{}bR�(�IHyr�5F��*D{�{q�]�Z�^u�VBH��ď�/��D�<����?�����S�/���xE����H�2�]&7��V}�Y���	Sy��'b��'��4�c�U�0�bc  ��|��ю�yBU���џ��J�8���@5玔B<�1f�!J՞q� �i�����'�B�'���]����A���J^k"Q�i{�����	֟�K|��V?5���P"�|)�N]3��)�"�7f�ă�4�?q+O���O~�Z�L��|�Q`ȣpV}B0�̪T|�2tB�^�f�'8bS��I����O���O�MP��	�s�~ڥMg�U�R����Ov���OD�3Ol�'�?��O��P��oΞ�c�G�^��;ܴ���O��n������Ɵ��ɀ����2��ƾ#�d0��O?1�P��i�b�'����'R�]��}�qcƕz^��GSЋ���6M�O��lZ�`��ퟨ�ɡ���<Yp�3`�D���E�`��ʆ���Q,�)��yR�'���p���?هk�h���&�R��Wh�y�6�'�2�'��L�>�-O��D�� ���B��A	�Y�2��+�>*Op�ǚ���ޟ���埸�s�+E�R`cF�I�h�e�Mk��?�6S�\�'�b\�X�i��!�FŢ5˺a��)�
����>Q�.�W~"�'U��'��P�֝�4�����B�bj�0�w.	?"�~6m�S}"V���	Zy2�'�b�'@ E�Q���%+���׍�}
@� �j6�y��'��'���'/�i>��OA��CqD[�PJ&���*�R�z-Rٴ��$�ON��?!��?��o}��D�7�0��t�v�@�J��Mc���?���?�)O��C�D�5�g��f����PB�t�h%��� �M{�����O���O���5O�'S2���D�VH���D+!�ڴ�?9����$�O,��O��'��Ά�gl��y��9b��]��ɫa\�ꓘ?)���?�$(d~rZ�|��>+xؒ>M��Ty�D4��mZOy��'J�7��Ol�$�OV�Dt}Zw��	�ԉ��F�l\�e�ٴ�?������'r�Ix�'VB���N�KL� ��ܝ=�x�0���Ц-����H�	����O�˓L/
1;�O�
T�\��3�ȼ¸l3�ie���'vrS������)���$Q�Q@ŋ6.�$��i���'��'����O*�I*3h5	�/��Xɜ����Ƿ��c��D�+�	����I�L�UJ2/~��N��'�( � ���MK��?q�T�X�'��_�\�i��i��!w�,U�ǅ�^�2I�c�>9@c�p~��'@Zf��'��i݅����=��4*T��;*�B�By�D��'.�	ӟĔ'/��'M�6]�:�	\ QBq���6���(�O���O
�$�O6��|�B<��H���Y��V��:M��R���ɦ��'=�\���	ϟ��	Tx ��g�H���@���N�X7,W�#�P�O��OP���G��5����O����/JTx��kR8j�������e�INy2�'��'��q�'p��O��I�̌=,�խ�&�!��iO��'���'8�y�����O���O2<S3������T�ѩp�v�)b�ͦ9�IHy��'	����O �X��s��=��]�9�씪��<i�$*��i��	��PS�4�?���?a�i�i݉��脵d��
�Ε�0��]B�i����O
�0�2Oj9��y��I�8r8�\�pͅf�z(�����=֛��'��7��O��D�Oz���u}"W�p�a���X�q1��?gt��&���M�Wύ�<����"������U�J�en]���Q5����Á$�M��?)��?Q��x�'���O��9�+U�.T�1��úvx`��iD�')�H�!6��Ob�D�O���Չ�>�(+P �@����S)����Iڟ$Z�}��'�ɧ5�oTSa���#�ܨ/VP�AF�C����Y�1OH���Oj�$-�dg��j��÷*&b(ъ��M�d�$�O�Oj��O0�� py�u@5F�@��!�O�}���XG@�<Y,O��$�OF�D1�i��|"A���+�D�K2��$+��Q/�E}r�'N|b�'O�i� �ybA&@��]�2H�L؉�d�'�,��?���?Qg��Dj!�)ؿ��ũ�"j:���W1O��$l�Ο�'�"�':ҍԎ���>!6�_�$�3�Z�^kP���ɦ��I̟X�'�rA)�)�O4��]EZ���S�И�rש5_��$���I�Ċ ��x&�D��ESL��D��54�`���^�Z	o�iyR�'�f6m�p���'U&?9�%*4J�cwƕJ�-�ĠT���	�d���W㟘&���}���׿Tl��1t��?�0���G���I�M���?����?�7�x��'��¢�	����1Ǉ(*�ac�s�.�0a�O�O>�I%'Ƕ, ���6�+�ȟ�2}��J�4�?����?��#��'���'W�dӒ7D��ANĹ?+���̇
k�֖|B��yʟ��D�OP��_�J��O|�@xrb�5N>-m��|�	���'>��|Zc �=��
�&bJ�$�?j�t責O�0@fN�O�˓�?���?�O?�Ha��&P�Z���� �hav��#	r����>������?���u�N�h��W�O���ٓ̀v�v`���?�,O��D�O��$3�I��|r  ]1F�� n9xm����B���'�������Y�㟰�j�R@�(q'G�?q0h�k�����O���ON$>��K|RPʖ7)Y�T�E֯M�^ �თ�6�'�';"�'̼@��d�F�,�c�U�O���ySɂ�ab���'O�Y���I��'�?���#��&jn	����# p��i�Y쓽��O(�֝�C�!��0oLm�)*�@��񄘓U�XIk�E҃j���rюcЉ9���|d\�H+	 �0pPp���|��X��8+�r�Wn�9I���)�W�Ow�8�a��z��s$i��HM$��5�.�"PK�l�3]��h��P���9�!d�A���� 6�����)$*Y��)ʚ"xP! �فP�Da1!��]���9a�M�E�ւ=��S����oϬ	r�|���̇7��Dإ-6��|��eʊg;�����J�G�J\blȢJ�ܘv�ɍ#�z<�P�_� 6�YxfϷH0��V�q8�g+jx��4�?���?A/O&���O���!	�"�J�qӃ��]�4���O����, �˰mⶇ�w8��k椃( ��!�p:�yڡɃ#'L��7@a�|��
߆k����	*�`����Q*T�D��Ĥ�BlP�I$F���Ot�=�)O��jg��K�lE����.i�X��R"Oj�������Q����<�+MI@���)�<i2��-Z~���H�v۠��a�ƍ�>e�4JT�c��'C�^���I�̧g��)kv�%�J���A�=~�P��$ �$��0���ir�@����i�Ӈ@�ZR�3������9`"��gD�S�* �ϓ�������i'��IB.Ş1.���l�q�'�џ�1����w��qԢC;��)��3D�h� '>("t"�� ��P��q���Op�G��3P���	H�$��n?���T��}�X�z&۲�y��'�r�'q�*�-��~@@t�Fo�F}*���!�9o��5 ��xcƤړ�I>
=�)�"-� �4�)��t�5����7H�v��M;%ɚ��(O�%� �'��IS0X�(C׏�py���3 "f�$/�OV���G�+�b��!gީ="yk��'�O�h�u��.��4Z0EG�_��E ?O^%@��NC}r�'g�O*��'0�EB8�o_	/��p��p ���ƫ1�:��$DV}*��c>�����s�X4[��H�z�#��M�N�VeBD���6���X�"~��!�t5�BGA&b�X�xWM�"M{ܼ)�O�����	G~J~BI>��5�Z0�T Q�І�a�<i�d��j�4�QGϐ�\;t����Q[�'kH#=�O�<�TCY2�^��8"2�@B�O8�D��O�p�nZ4�I՟(�'��'?h�b9�`�-��X� ���'��	tÞ�[����1Ov$�F@��[˚#w��9��D��O`�E���S(LL!�8�4��-^-|��C`P�a�pd��,������O���%ړ��� L\�9�)/t ĺ�aG�!�,f�L��)˼T��Q����@�~=Ezʟ�ʓ[��i�5�a�U�"�蠳m�)�>�qW�'���'��IƟ|���D��d��9D^��ܴP�`d�F�Kd�ܡ��]� H`|���NR^Ȩ�O�(�v=J�+ r�1 �%�{-���r��+$�H���ý��'=t9�3&X�,�l�`Aj 4�b�w����<�����2�ӧ(L�{��Р[@�X�l x�C�I5xt޵�C&ٌ/T�J���=� ��঍B�4�򄈦,��n���It��B�VFm� !E*Hz��9�ş-�y�'��'LreC��'1O�&a�=�$Γ�WcЕ�'C�(Ӏ�<�����O�9�A
z�l[��UjP	��䕱"��dLȐ��hi��a��)��"O� ��;��^�o|(t�I�����'�F�O�W�ؤq��)�$�K<G�@Pz�'"���֏��$�Ot�����O*�d�4tE��P�!R������GO�Q���$�ʧ���?!��$0F�8�.ȴ�bI!r�1r�� C�ɧ����;1݊�J@ע_�6�iYhԼ��'d��'����OH�+e�W%;~�d`���>F0�H�9OX��+�O�E�ՀW��H8�h�b��j��ɯ�HO�S��Ѫ/�ҝ�u�p�
��I��$!�M�9�M����?�������O��0$�>p��ᚠm���h%��J���Q9���3׋*lO�T�p�_�)�M�#$�w�%Z'�O��1�� ���D�,��,Д�A�h��uH�M}f�L�Mi���O��ԟ�ϟ �'p�����Q���Oü;� �'�Bt����*5N
��HH�]�Ṉ"�;�S�T��O�VT�P�E�u��ܫ� ��KC!�$��]��y���Q�nq` oUo�!�Ĕ Y�2�a 	�7:E�wn^�&�!�A��Urۓ���]3�p��F]�<�G�^=��0G/8(�"`\�<�f�Xò	���7!�pc�f@�<Yt�`�5�QD�7Gȭ;0TP�<���.J��cg,^���D�G�<�M��)���F�=
r�tk�B�l�<�2�Kz��L��j�~���'M�}�<�Q��(0����B�?	�����u�<�L�$=�&�St`��wJt�p`�Zy�<I�e��Kt�I$␗[=X�(uCM�<1C`X�B�0i��
�"�P0G�_�<��`��C\�d�C��v����v�<���37�����O�'��5Q��J�<Y�c��ܡ&�SUvLQ�I�H�<AFK��2L�7'��?�DU;��j�<)�#
	:cL��(��`��B�<� �<BZp��,��]@�J}�<9�.&	��ib� RI�H����{�<��(F
��(���@{"E@a�y�<!��X�8��q�C"�^iz#ŀv�<�̝ 8��(�buc�Dz��L�<�0O"p�v���K�"[�0%j��[E�<��'_�EB�xAꎪ�칱�g�E�<9ʋj�pv*ՠ��=y�k|�<a6�@g�4X׫ GJmz��x�<a�;d�2tآ�ٙI�$Y�&��M�<9t�����k��Z�m�8�9"���<�2nFC8Hȃ����N�� �e�<���`�썚�c�t���ۦ�Of�<1�g_�G�04"�"W�{G�6�"T�H����"yBy��iM�.�Aj'&D�@� ˈQrHM���8a�Q��"D�t2k �qr�ݛ$�zBi� �?D�����bD���AK1W���"D����"S)@��Jqa�}�@d҆m?D�����Eh�ܝ� M�8@*`�>D���f�v��9�O3f�0��@�&D�P�G��)5��S�K߶5�Pe�D*D��ir�c���1�5Zph���'D���⦊2h�M�B�\#JmV�Ke+D�Ȫq�ɗ.�v`ñMY�3�2x�2�)D���D��*ЀK`�U��$�`��'D�`� �>M ���"*U���$D��s ���əd`I�V5�dB8D�d��͗�L��M$J��LU:@A9D�4Y�㛩ed2�!&,��O~rd�$}�L�Ȓ]�S�'0'`ax�jT�hN y �$��r+݅ȓZTD�g��X	D04h�l��=Y��2v��� ��H�EK�n��e ��xK�aj�
Oj���#����GH/���񫜖oȞ�q
�'�©�"c4"�J	�B.J>��Ǔaؘ�j�`*扐o"22�4Iޞ0a1�� c�xC�	�3���a���8϶��f�$�nO�Mۗ(�|�S�'R�D勱��3(�5���;-�,��C�,2#e�m]R�	�m�TU�ȓ,��Ҁ�V|p��%U$j�Q���B=	!���7�!J���Y��I�� �fkХ{5P�� zn�U#�'�A`���@��@PD��c�T���'S(�0�ذ �bt� �ڿ?�ݓ�']��зD֗	'��s�n�+��<J�'{��A�:MG<��H�F
tQ�'���� ��qL�i����'I�����'���!�ǀ-;���
ŢڔK-ؕ��'��H���[���"EJ>���'�p '�x^�u"" ]
Ut����'7E��(N�O��UZ�-ƺI`�l��'�0� 6��5	�Ļ�����)h�'�\�	�<���20�$� ��'�Z�*B�E�BikT��6z�~<�M>i����j�6��@��$m�A2�� �!��D���C��Qclx3P�H6��O�;��'���b"x�� aaCU�4 �'RR ����|H�+�hF�{�cu�xh!�d%6�}� �)צq`����DyZw��Sf��
�@!�����!4WHx��D7�nm`��2�y�]c�)C��W�Y �:Ui�99�D3�c�Do~��AH?E��'���:�R!�(d�জ.�9K�'Q��C���e�Z�C��A,vW��I�'��AR�� -�`s���0<�ʏ!��Vmzi�4�Uk��h�C��}$Jp[��@�wSt��fX�*���ɒ��dy3M'�Hæ�L�/6<���,�υ͞&�O�X�XT�%��Iy��|���&a1�`�b)��6���CL*Upu��"O��ذ�E���10B���H[B�]�McJ��u/�>C�T0�h��e��n��C'�:�@!�60$��xi��􍓶Xp4qB�n�7?jp��+�_8h��O`eF}���J<�?�a���S�
�T��S"f����^QX�b%���o&D�p�퓝b����Ζ?c�H��v�� ��+סP9hl�1�$�O��q��9  �P�hҽE��dc��|�`M�ea��=M~�@/�?%>�[�'Ԉ\H�z�L�|�^-��O-D�ܣ��·O!dU��AA�E�$�QBF�Zk�}�JF��X�O���H򧌜�<��]Q�
�4Y���RH<ahY��jG@�	��)�d�S<d�D�6� e����V<�A�闗(��Z��M�S�N�J3�M=L}^�Q�2<ON�H7�]�^�S���Oة�Fٚ^�"	˴��[�d3a�.Đ��a&�Px�14�A�9`x����&Ii�Aꖧ$���	��@蒯�0�e���/���|r�2/1.�E�Г:��ѫ���D�<	�B�' ��[R��� 3SV�0��]sJ��e5Z1˥�P}��d���y�U���Z�
j��@�����yr$Вn��Z���  $)	Q��-��$�l,(%AY�2�n�9`Y(䑞��\0J@���K�0M����+\O��q	\�<;b��V��/0U�$O1v��/B�a��q�Q-  ra3�>�O�`���S	CV}���'�,�Z ��K-�r�-N>�$[�-G\��ԟ�u����vY6A�&S�9�d� �A�?�pC���(�z�HADզ.s��;�9q��X���G�T�Tl�6��C\`�C���,O�����W�׿[ᄥ�G��/F�~�Sa�<q��ѩ+�j-j�EH
,���� 7��lZ��˓h���5�yZm�&�]�L���#O�J��o��Qޤ	�i-�O\��"eX��U�&�!#�!)%D�.=�X�X�Dͫ*9�6���$�̓�Խ��+,����9ǧ�0�@4 gP�Fx�*�4�w�_�q�`�['�*�M�矤Ia��u��	�K@<eN�y�\�T&L�S��'���g*�O�μ��f�* Qp� �O�:&rA���܋��� *�M�g���� R�ZƤZQ�9�!d�>�j0�"Od�����:4be�G�o���HVMF�y�0BT�SC�i>�	�j}!�T��y��@�O?��EҲYo܄@���x��P��:�r��D�k�>����t8@����0iq�4�@'��g�$I�<�l:몴�nN�=�L�O���f>?yF)�
4��T+��̾�~rțKb�%�"��>2�TM[�O��� �Ll���'(3,O��;Q� Z3���$��Qeհ]�0D)OH���W��f͂�A����.O��؁)b�U��g �8��%�j]'V�xu�<������%)��:lg�T�$��m���*��"n�����]��]�BA)?Q��ܹ��GO�pqd=�̸q�g���f��Fj^t� L�eY�̺1��sqO��̹s�o�r�hѬN�x��H8��4��'���� J�E�G_9� X7`��
��O�h���9>�U�&ݶ#h@P���x�!\�-�Ё�'8��c0�z݅��
j��}�RmU0q�����U����Q�'��c(�(^4�ԣ�@8�D1�w� ����5;�;�I������V��
 �!8J�ط�[;��a:�n=�韔8 �-\�k�IA�Q/�����	�/a"]�4����袓� $~<�4��E�M]2��^B��׀K�Wy6t� Mםc�R���?;�V�J�F4��O����h ��O��i�IS�@R��JD'�D����=%'��#�&��;�N��N��B�����(�⟄���5 �t�ɱ62h��5CJ(!�.qY�]7��>�e�#^���{#D��H9n\B���$��8�1��w�$��Ǔ_�.#^3����L�[��=SaXo����YF�h%�"zN�g�
*.^����$U�hY�qF k�Pp�F��֏@�?�L�ZpBº(��ib��C��0<�b�ǢS��D��G;]��l�C�����Y�S���ߖ�z�N:VZ1�'̤<��$�7���ւɦ@��+��ĝ�P�3���B��0J�;(̙q��3x^ *�@)c̨5�ʍ;CP�=y�¦x�xH�	D�f�8)���7p,m�Ç�+a}�P�w.�R�݃�8A#q�F�%
�����o����$ϲHB̨PA�J��� � �*��խx�� y��B��nU)�R%!t�*�E��<5������#e.���IlzL�E�G<(q���8s6݀��*�I%jX��`�\n1OX���`�Xf�,���R�PФ�'�fQ���ঙɄ+�c�BԱRH������>���jT#>9�d�.8Q���I�xmt��N��T����x��WN�Y`��S�E\a�܍�iݵ��o7�U�R fFـ1�@ !���K^��&���'ސ�Pa%�a�gy�@	7�Ay��Wk-BT! �O��~��C=������9zZ�-A�E�"m@�uaB�H�`X�1#uT.6���vf9�S�\i ���&	�x�Ж`��pm#?I�O0g�4�?�2���\� ��D�5o����4��YP���H�tX��A��>�[��r�,�2N��PѠ��S�L��'��p����f�S�OB$���V�>�;����.�����4�0��$K§>'�z�#<O�]�7�E-G4��e�P�FN�1 �x�ց��>�O�H��s��%�VH��'Z��D�R2��v�l����-1�Ь�4�I�H��Z��]��52bdϜ��d_%B�Ι���#��4b�A�pџ�8c"SD�O*\��M�.�Ll�]���U��'�� �i�)]k�d0�ޒ�0��'+.
橐'+\؋DHQ~e(P��'�R�26�`X䫞+pOdu��'��BS��"`�)ಅЄnr���'����Fԓp��U!�C �i��<Z�'o���S0{l�E�ma ���'��<���!W��� ��a*�I��'j	���?&oT����X�l5r�'�`�a"JW����@曹Km����'F��:�C�#��y�$#�0<5���'~�æMȅ\'.��3lB&7o��y� ֟/8]x�H�=R�����9�y�N���ܻ���#kΊ`MX��y�++>z=��&��g�X�R�Z��y�L�?[L�H�D��<d�tl��N�yr̀��4��$ˡ��X�����y2mJ�"�X@QM $>��j�lʎ�y2%G�_P�˅��f�P��Ҏ� �y�("{�l:6n�)?�	IN��y�$���2�N$~@����y
� ܌��G9I1C4�U�,��"O��QV�յm@��(C3��	c"O*qQ�2Ȋ�� hN�s|j9�"OA�D�0���H���҆"O��x�۩l^H0¡5k��P�"OX��FB�&|����߂m��t�5"O@��Iτs#�9S��
&	��'k	����	�`�8��U'aT�	�'�F�(�K�VRw+�#�Tu��'�� �*���Ћ�ˀ6!tx��'�*y�K�8M��	f@S��\��'/Z�#�cÁ}̸�p�R���̉�'��ܐ��D&w�"5C��`�=a�'�� w��$Zm2�G�3Q0		�'5��c���3
����A��l��'B��h��N���B,M�P��A
�'� ���
c��1���X���	�')�	�#H�*YA��Y�{����	�'�n�"2��L��R7c�(�0��'�T��%�j.��Uf�t���K�'�xkċ��"�v�"V.��Z
�'������Ў�zgh��6�����'mN�k���?V6����L��"��`��'�����#Ƣc�^lY����H�R�'���h借�Lʜ����J #�p��'���j�j�'�T�(�(U�x3p��'�dI��8|{f��>�H|��'Rn��gOܚz� ��R�5�`��'l��X��ڌމ��W�5��yB�'���2WZ���J�Z�.,[�'�8qÊ� ��� z�I!�`�<�q��R��<�%�*~ ���\�<�a��3.� ��㊋C�yǹu�<)�#���rC�w攑!M�<��J<����eOq��Ã�Iq�<iG�B=]xQ:*Z�p���Մm�<�e��3�,�Cu@ϱ9�<\sBM�d�<U��+a��K�D�za��G1D��37 �9S�0̑�5�D�J�.D�T*��ˣ?:)b�Kʣdp�I��>D���`Y*l���r����\�*>D�88���%AVxP� �ߔ:����&�=D�|�Eʄ4r����dߐ�3�'!D�4@��ND@���cH���^���?D�@@�H )�
�E�/�HxȦ,<D�8I�	H[�$�`��J�$�kUb:D��S�fXC��4�p��4��i5�"D�<"��K�b�1�BI�:o��X�/ D��!��Mx�B3'ۆRr��3$�!D�l��X4>�
Uɓ��*Zz��em:D��O�0;aD�F�D|��Q-.D��bP)�%�L�ZF"�Kƪ�h�(D���B�U�\����_��FS�:D����~�Z�P���ug3D��(a���r���%h�
��QN3D�֠� ���Z��g4+u /D���!S�< �{�)ׯ �V(�. D�4b�nG�K ���@G�L�f)"D����ϙl��B5D�2I�����!D��kDK�C2�t�"�0K���a��?D����@�� ,��.d;��Ԡ>D�p{7%��u���"5G�I�d�=D��QSe�b��Ф�sWz���:D�t�� �w�V�pƄ��v�:��"D�� �����Q��0�"�>5��t�"O���C���L�s �D�*@�$�O&�=E��+~*�#�23a��x��W��y�\�&���P���%���h���(OT����H5��#&iE� ����� ��!�d�%G��e:2'@<lrp���3u!�d&#riRoڿʜ��GB$0\!��>���2`��O�����*i[!�D@�_Ø�kY" .����d0!�DkZ^����0�@�1�E�<#!���q��]�͋9`��p�$M>u	!��8m�����
���#�@��!�D�	��Q�d

�2�f0��a�!��[�,�|��UĊ���)�t@(�!�dͅ_�Z|[�K�a��Y; �Х
�!��
�(������
-����&>�!�d��'�z�(�]e�T� O���!��'��S���.",���aV�/2�C�I@i�s�J�4ev��T�ֳ�6m-� )Ȁ�z"	qa�"^,v�a�4D��3F��h���I
9�V�K�J=D�D(����EHZ\�4}��d'D�r��tA
��7W'�,izJ&D����M�C�q$,�f��9��%D��*��S
��\ �	ʩ
h�����$D��@���U1xM�rg[#6h�ѱ�!��oZ\bԀF��B�t0°j�d�B�ɞ9��})BQ�vn�
��X4?u
B䉚x��_>�� X�m��C�	�;�>�ڦ`G91�I��!Ԫ"<�C�ɜQ��pi� �$s�� J4 R�Xs4B�I82A���[,`W��[E`��gH�C��N�f�K���#�|�x�02�'�F����P�X��އ����'��5�F�]������Yr^���	�'(h����!5ָ�'�F%8�� �b�fA3�k��D�N`;�'��D�ua�3je��h�CB�0�	�'�t0'�r��� ���MHp��	�'��M��F1A���B@C>.P���'hx �O]&1��ͱ������r�'n !��D��@�
肥�'&R�Q�']�|Ch��G1~�z�#�'���Zc�-�ɚ���!o��)��'^< �ïH���ЁiT�w�P܈�'�P�c�d�50oBd���s"	�
�'-*����H0EF(m�� �FQ

�'���eO�8s��`�6o�6��	�'=� ��,E.)(ٰ4�Nn��X	�'��ͩ#��&B2p��m��z�͙�'�\�!�ķ'�:�r"B�zn2Tش�Px� �)h�*=Zv	&�6��'����y�G���%Zc7$֠�k����y��F3:�� C���j�(i����y�5Dn�qTy�r�[fm\�y��J�,0�)R��d�r��`<�y2��d<(�,]�%�<�Ł��y�n�5"� �b�N��v�c�o��yK4"� �N��daq���<�yRD��V��<�rc�(BK �Bc�5�y��g�r�Q��٘O������.�y"�ym�P�E��{����sH�yboE�xqysA()��|sI
��y�j>vF������.Q:"J�;�y
� J1�vl�F������1%^�l�"OR����A�U��L�1R"O��;��z;~�)��Ė+�T)��"OF�ST�ʈqd�Q�.P�hҞ]�e"O�X��	>1�,]��J=mĸ`"P"O�e�DNQ&3JL�*Y�I�jT��"O��WA	!@|���G�1l�r��e"O�1j I^)]��R(��1��q�g"O���o��,�ƹ��ĉ)����"Op}�Gn�*(Dx��`ŭCo��W"O��fFǾp;���&��pQH��"O�����N�t�����J�	8>���"Oia*1n��M(���J��h¤"O�$�bɉ�V�x��jW8ḧzC"O�� ��:1,��Y�C�zXr8�&"O��P�#5Y�� 0Ç�fh�2"O����-W2:89�� jL"Ը "O8�PVk��r�I���A"l-Ј+"Op��@	�<V�갓�F	�v�y"O��@�Cm$��vc�+��I#�"O�P���I���8c@۾`��'nqO�ţ /U�X²U�DH��{+�a�"OJ$BL�}0���eI�"�=��O���	�'X�.�r���>:>(�E�C9C�!��=,�8�0nZ�;Y��AC�'	�!���B#4$f�y��N�iNL�"Ob�
p`=�(��`�y���@"O2i�cl��M�D���(��vRhA�Id�OGB%!D �8����_�~��91�',8\`��G�w��2�m�2le��C�'��x*��8F- |"#�׾d�B���'�8�� �F
:T.T�uEǣ+"�!P��(O תR����QKɯf,�#�"O�U.����5�4�rMC���:�!�<"T��A5�H�ȅ�Q�|�!�dN�5�R� A፯�$�HA[�k\!���x�@Q���M	\f� Ӽj@!�d�	kW<���a����A@\�D,!�D�&���qh�9�	/��X!���+xl�˕�F�
:ҎҺ!�!��Gx��2f �~1J�-G?4�!��8%�\�⤂+o0�Q���P�n�!�S�}D�	Gb9�HM�K��!�Q6UL��;�hA��`�IF�Eh!�$�1��Y��,��ՅΉ�&x�6"Ox9*P
 z�3�䎌V}�Q��"Oа��̜�q�@�QiN�	���"O�
g�U�k�0�mf��ehU"O,T��vT�eJ�*�d�r(a�"O^��D�\�b��=����X��M��"Opi@��I�4$�ے�&twtSV"O���R*N�:4������@q.�!�"O"}z�)S�|�2	�ȸp� (�"O�q���'+Ȳ@
N�:�Y�"O��b#/5p���҈Ѿ60F��S"O!S��B�� �e(1|,@�"O8X�C�A�޵%(�I���"O8�㔮�!D�B-�&G�\�̡�"O|�c�U3C76<����[�4Qb"O��1��OGCh�1�&�&��(�w"O8��um�#m�$���D?X�TKV"Ovh�qc׎~ �U"��L��� "Oљ@�ʪk �2��5�JD��"O`|IpCJ dj����!C���1"O� �� �L;Z��1e�!�☁�"Oz��3�2y�1�Bǟ����"O8����A�����H�/l����"OX�� Jא1�N4���gdtU�6"Ovx��R�@��d�&�)S���"OJ ���9�Ҵ��f�21V��`"O�m
0!��u�� ��D(�	�"O��9���*V�Lb���%&�yu"O�p������R�n��Hr�"OPm1��U{5�A�pM�7c,�RU"O��C �
�!�,U���!e(���"OL��kV����4L�ZF"O��X�\1Ć��M�hs�I��"O�ő�&��?�e���$�3"Ob� ��V
�jŢ�ΰk�!Pr"O�Y���Ӆ^��3H�2P�L R"O���
PF�R�h������"O��c �J2�A�!�9-��+r"O�!�MLm:	�ao˭q����"O����J�q6~�SC.��\%�`0"O�M1W�*}y� rM�	����"On����y��q���߄2 ���"O�|��R5�n�QM�
Iy�Y�"Of]�b��m�&՘PM��q�ʑx�"O��2��;����N�u�5�E"OhPy�hް �mD))����"OT("d(��b�1ɛ�Z�2QS�"O� �r��<�,��)�t�U:�"OjMCVʆ+D����1��SE@�[R"O�Hs��˶*��X�AN6-;vqi�"OJ�"��9J�+��$�d��"O,�s��ē>�$�@��>䉈�"O$�@AO�c"��Zbi�6Nd�g"O6\�6锿_�ѵ�1 (8b�"OP�BG�1�4�Q��߭]�����"O��aH�	�8-��2��ȱ"O��ʴl�'a��� %��
��7"O�9�o�6`Ű����чwMp$�g"O���4i� 3�:�Ic!��xKpH
�"O�0:��F�tDi���Z6�1`"O�c#ه.s��˅M�f'L�;B"OH����|�aB��,km��)W"O<��%n�LM�M߆$^R0�#"O*	x@�٨�Ĩ��L�>y\N� �"O�P�-[�2����]�gW�!kd"O�%M��|�px{��A� j�ՊB"O�E�g��%(�<�"eF>	,nl[�"O��"�N�T��H��i�b��1��"OU��G�1a2����ڬH���P'"O���7+�(I�Xe��t\�9b"Ot,��צ�y�"X�!ǔI1�"Ot��ë��8���;�g��Y�HEI�"O�0R5ˁQ���Cv��7g��	�"O��82
]�mD�` �N����9�"O `�&��P2��RT�D�E`��w"O�\fe_����k�O��/�Z}�"O�\�C�ޘc/�$��+S�V���#b"O���.�p�O%�hIx�"O�H!�LS)TIE�WB
@��q�@"Oҵ�&t�إ�@N~U��"O�����ݻV�����HZ29�\Q*g"O� H�M�00�ǇH� �N�A�"OR$#M��$�1�B;x*�-	�"O*����4^uP���
 K�"O� YH��VqQ@�`�l����"O*�CŧQ�<i�Ub�2�(8y�"OB́�oTTߔ���G��jX
�"Olz�Ē����2g�+�� 1"O>@ �GO/�$s�5B�=�v"O4�w�[�7�ػ�b�E�HH��"O�Æ(�nT��;�a�QJ���"O�����\3 �3�J��34�I "O`H{��L�E��43 T9 �"O�ē!��D�l`2%L��u#�"O�9kG�~&4*�-��(�"S"O�P�C�]_�E��"8�N���"O0�X�	�~����L6O �-�&"Oz��쟞 ^`A*�4[����"O�<�b��p�.ءI� *W0qc�"O��rE(��=d$鲓���Bl�4(E"OX�C�/�B��(1�A�����"O\̻4��% ����� � yzL��"O�,��nV�Xc�[�w�n!�`"OP�ae
��b���P���u�ba�"OFx@���9p�UzR�U�JM.M�"O��)�C����! H4^�h<��"O�ܱ$j�X�^�b!)ޔ�Q8�"OРP)��/V�� ��_���"O��ʣ$��TMp$C�\��4"O�dZ��N0'��h�i�9b��"O��Хd�<w�L�#�T�X��;�"O� SG�ػ(6h�#�@Q|��"O,��A	άVH�$+3��0FN�-��"Ot�K���A�4���I<\5*t�"O��SFI	N�P�ǩմ$'
3"OxQ��	�#5Ь{���� �K�"Ob%DOњT��E�0p��l��"O�ԄJ�!������5�n)�"O� ��	>�� �V�=	(�%��"O��A�UBz��'$�Ql9�r"OB���6>-��ɗ�ڨj7"O
!�TĤL�J�A��!�d|�"O"��i�=���>��p��"O�11KA0V��a�OZ�7�xe��"O�T���)�D�"�M=��,�"Or�᳃H~�P֍��k�
�J�"O�-�Re�Z�T<kЌ�>��]7"OJDk�;4`j	xd,� Kt��"O"�;�7CY�|�P��<v���"O>��e��o{�HX�Z�T/x��D"O�`�"M�"����T@[+H \�3�"O�$�1)˗y�s��շF㨠yA"O]�ahL�Ѩ���.ćU�Ь%"O*y+7�_�	����P8��) "O��Є0�N��Eh�U�����"O��c����3��J�f�-V*�00"O,̢����4��,y�σ9ɀ�"O�A���F�2�ع��EԔI߀��t"O�h�K�]���N��Hbj�"O
hȱME�F9�%��`P��@�"O�`ՒM��]Y����V�ܕ��"O���Ehĭ:�����A'2�ȡ�"O�e5�	�`��<�v �n�h�bW"Ot<5"��q^h�	��H���ɓ"Ozy���=��E�2(H�.���f"O�	���h���ض&P�U	V�"O�$�2OZ8	���F
<L��"OX��&a��Th�����U�5� ��"O� �d!��-��a��ܑ�T��r"O�ʠ��oK֑��Ę��8D"O� ��Hک<|���L ���6"O��+2@'+*!;5K�`�6IK�"Old2 �w"P�s���>llɂw"Ob��͗7����7i�`/H��R"O�X��7|�JyB�匞l8��g"O|1��LF�d���z�Z�M�d� "O��`7h�=DkZ!�O�O���s�"O��Y6���|���"%�z��lʥ"O�U ���Y�~���D�##�hQs1"Oa"���Q��\��
^EA�"O$M��l!����� �ru��"O���'���]fN�����l��["O������ ��$�'�ު;Y��YU"Oh`�@�X$v��DАFO�OE�S""O�Q�qb�8o��z�EY�U(��0"OZ��A�Z�,*E�BF	��"O�L���U�*����㐍`�NM�"ObX��c��~,p��~bL�"O����.5i�,I���AV��A�"O����H��.� )�A�A PLYq"O����N����G�rk��!r�|��'�ԩ�r�Y	��I
#��#&�N1��'�z0� Q�{8"" �7����'H,��mS�rBvAz�'��,��-B�!�4O�63��	�'��t��m��=}F�@�R>�]�'D�XC֡E�)���g�ݗB+0��'P�z��O�:i��f�ˊ4@(���'� <
��͚F`R9{W�\�%��U������5Ax��c�=�Z���Cv�!�W�~������L�4���
�!�Ē�i<�l!�J�"I��pG�B�!��[�>�I�6�7>~a�V'S0�џ�D�ԁ�9��		��ȡx���)6�y�\+*�<�&������W��+�y�2�*P�a�OwU8'����yr��d�B�	cb	�Đ[v/�y�٠K�P F@��U[�mӥY5�yr�����[DgA�N�&��R �$�yr%=r �|SA��;N	,���T�yŧ�V����oڙئY7��xb��v�t)cN�s����u�F
ZV!�d������P/�z	.�*M�'�ў�>��Ɗ�1"$� �֟4o�e�%�#D���&+Ԗ,0�b�-.h�Bq�"D�(�"CїE�(�C R."g�T1��!D��Vfܭ_��lp*�"n
��$�>D��3 �:#�|�SJK�|���s�9ړ�0|����+�� �&`�p�7�o�<���C$`4�d�!mz�:���� m�<YrL,,�1��r^f ���h�<�T���l��Lu��Xc�� O�<1FiO�^<a��\6��%bI�<Q���("���1�A	K��#cI�<I��H�{�2 It�V
	S�aB��@�'=�	Z�Oe���T�)B��e�P�o��T9��x�iG��D����-�Ȍ:W̞���x��X�=��������y��r�
��p�!��X1!�f|XaaY-1��s�(Ɲ1�!�DR�R��*�M�G�����:!�߶@�t�y@�8`*"쒐늑c:!��|�MB�� ��YB��Ζ(+�'���5�)� j�S��Of��8�	ч1����6"Oz@çm�9+P�qF��HE�2�'���	}Q�h�2���\�sn�<B�8C�I�+Z���[X���"e�	�C�I9L����d}7PH��`)<+C��?F��!�f�-��l��V�B��,(ҰI�����,4i�0I��B�ɤh}<p�ԧٟ�9
���}��C�	�~������J��g�Q-r�v�HG{J?�K�CW2�,�e�+T!� �C˷<��_`��#��]�~�L$#6�JI��ȓy��sT���tE��_1|�p�ȓ)@��)���P�v��ti�*�ZɆȓ/l%9�KT(,`����h<p��	���d̓m��dY����Ro6|�sA��bN�����	���O<�b��>��ȓ$��Bd�%p����6�Μ
RE�ȓWў0���G]=��icb5-ά��j�n(���30�$�)�b���W��0�D�e�Zq�C!Q/��݇�NR���&j¥~�B	�e�Tf
���7�����	Q��8YE$XiG u��i�p;���U��IX�I�	bI�݇ȓ��Y	U��3~�|��Gib\�?I�Z��0se��7H�b��׿,O:��ȓ��B��́LF�Z�D:;�>���#� �IMV�gR��2󋙲%�rq�ȓ�b�
#�\�b쑐h�?~0E�?y�Y�dŘe�5�^�9Qi&h����	�<��NF{(���BX^A�%�Cl�<Y�1K�J�,ߗC����TaL��<��~��j��~�?��q�q�Ņ#�b���*�yRL[S��]!�$e��C�3�y��c��B�.�8n怼�ă�y��/>*�L �A`� A�b�F��y�πj�: �3U,RX� R���%�?Q/Op�O?Q��H_U2H��e
.6Hiw�h�<9���M�����N�x�c�b�<�ABP )G,��	�%�b�P�jCu�<Q��? t�Ҳ@�9j�X���Bs�<�����(��&��=JwAům�<�cI%o��[U� ��0���ZOy��)ʧh�T��Gꅤ^�0����)!@xɄ�Ix�'��y�S��): ��+4�Y�,ٸ(O��=E���!q��xJT'�6 
}�G"D�h���z��4.K>'iH�hB�5D�H`GLT`IҗJ	�*&HAs�5D�̓ᧉ�g;�9�a(����)��2D�d25A��Y����Do�8�9ʰ<y���ӯu}���
j�F(�1�֔F�.C�	#F�Z�saL�b"��+��N�C�ɷF�I"$
T8���.�'��B�f-�qR���&_�8��v�.�xB䉉GƦ)�%GDx,�1���TB䉍s6�2�(��ww,m�e�E�R=B�I�İ f���0|�vl�r�@C�ɢS�D,��#�>hy�:C�B�I&+�����@� Y����旐n\⟈�I[��~�4L�b�c�����ѭ'2Ѕ�*���QaJ��Lq��2�*]����ȓ.'\̨c�?NΌ�6Û1�|�ȓy��� w�V����$�01y��ȓf�~t��Yn���&��R,���Ɠ>Ќ��v��U����ȮU{����� ��I1�ͅ7s4%�'d��D5HW�	|�'���	��a�)�nI�Z�#ۈx�'*a|b��%�J �Mߢ���B�_��y"N�����;�&�� ̛�ْ�yr��*��T����.0�� CD"�y�&U:�ȱ�&�*-� �a��_��yB��5�����B��#0�&�y"�.��JcB��"�Ǖ#�y""�9*��$�0�f|s�a@?�y��N�>�Y3�ވ!:v�z�ꖂ�yr��������: W�U;�k���y%�/��-�ņ�-e��;4��y$yf��pk�I���hE���O�㟢|�N�j�l����Z�l�XiIE�<���U��(�[�.b�@F�B�<!�M 2�޽A�!��(��k�z�<A�Ŋ8{"d���=a$�(ÊJu�<��i2�C�ܻb��b��U�<� �/% pr�Ahzd�"P|�'?}00N).����t	(~�x���=D�LPp͋�d"b�SL��|�p|���-D��s�A׼3��Pf��VD���*��0|�Q��6��U�T�K����TkQN�<�'��(a�u҅ ��v��`'�Eb�<Iu&��2��@�!Y!�$���M�`�<YA�P�zX(%��)`�}е��Y����<���3NTUs���5A��Saf�S�<Q��,C�>1 l�Yl���e�<���O�+%H���? ����'Dߟ$��	n~bC\�4��ID'�r=J<Y�*�>�y"W<Q���k�>!+�)К�yB��'($�Kp�Xu�"��i�4�y���N\�̴֣r�Z!��QG�<9��W]8�ݲDB�[ZH���Wy��'h
�R��5B���ۢ��5&�M�
�'�^y�R��>!��I�I�K���
�'�f����MH�cG�Ld�X��'���:�IE�Er��ã!�Q4p��'���z��ɺ/�֡����)�~1A�'��0n�)wS��pԎWf�x��'k�8�H	
*h�Sϙ�Vy��[N>y�����O.���eۀW�M"g��w?� �'�tU�-ԃh��2S7��@���8�� �S�5�T����V��y�h��^1��O"�=�}ZTB�+[�xH��_�mb�&]D�<����-*�8�/<_6�Q��[�<Qw��N �E9��2F�k�k
ş�G{��I��k(C�Ḅw����h�v$ʓ�?	���߶������ʼ��㘿2�!򄋝����؝��iQ���{B�$G�����УNV{r�F��3�!�DZ�i��`�H�"U�A�NO��!��Y�2�x�`���sP Q��:�!��?#��`���N��̋�b�!�W0Ly���B׶��RK�O�!�ЋQ�d�y��%�\=C�/�
+�!���c��`�l��2���;�U�W�!�Ęr6�Ia�"������f�]&u�!�$�6�|���`7��D�g���'�����.^A�Ǉ[�C�ֹ��'�Q���" _��`���B h��'&f����ޟp�%Y!&�/���M>9���i�4_,,(u��A7v�xen��O�!򤖓�z�I��$8T��B�!�� ��Ha��%[B�9�XG2��"O���Fۏo��T����7;��if"O�Bt��	�`8��_OV�
R"O^x�sk�?H���Q 2B��p"OV-�Ca�G�>�!�i�#AC�8��Z����}�S�Of�}�W���LU�D�a\�K0�I��'����̐�U��l'ѥG�����'?�Tq����3o�A�D�c���'��ĸkY��Qs���4@��'�`u!�D�oFx�҂��FR�m��'�Ti�S��2��1(�#�?�)�'f���'R4A6���������'���B�T�85����u^н*�'��X��D0)�*��$l��' �J5�=+�hXq$��q5����'��k'�Г��ѵ 't����'qp��w`�j�#�g!e�|�+�'��y#�!�z* ��ۈ[T�("�'Jt ��9
��'�+��QB�"Or�#��zg����L7�\�5"Oґ��Ƥi+�q˱�<7v���"O����
a���D�O�Ҍ.�yrM�ր�:�GU���\�%^2�y�*�TQ�����c6t�F��?�y�a�{\(���8Zl��p�Ί��D%�O.iK�`�(�"=x�JxP1�S����I�,e�vH�V+y�D��-LB䉊y4�ѥHڿ,������� �4�=	
çK�l��n� 9\ɹc�I<]4�ĕ'ua~������r���*$@�mK��y�ļ0�-�s��Bi^v��,s�'�N\1ā�)x �`�
ͅf40yK���'!<��`�aXp��LUp��:
�'��ch�	hV%pl;��x	�'%Jh�q�+)��8b��X�Z�8	�'V�:���&3�U	ECzA�j��y�-Ү^�
��`F\*9��%��y�'։H��*PX4,��4{�)D��y�k�#Y(�u����U�4��� ��y"�(!Ib-��P4=����'É��y��V��f{K�5S�]��bC�yҦ��Q
�牾A%N]���D-�O�@�"Զx�Eᅎ�6;�T�A�"O`*f��y�@B4��v�lS�"O(�06EZ(W�~Q��_�@j��A�"O�)� �5�@�
6C۠S�P��"O�XV� �p�P�p���&,��9��"O��
��ɨW!�4�A�U(c*H�d"O(���H��T��,Y��D�F:�AG�'�ў"~zj��?:�E���O a\}�׃�����0>I��I+
��xW�Ĥ/P�uK��XA�<��Ê�R̢!�� [�Q�^{�f_U�<�ů�5HU���� �V���"�c Q�<�&M�J�ְ3囋�L�2�M�<�D�4�dE1v
tp�EBV�Do�<��G�4e��ik��W���)AF[d���hO�'�n��i �?zJ�i��œ���"O(Ab0O�D�����d��a1ڽ�U"OL�Qɓ�R���ew.Z�ٖ"O���"힆RʌJ7�S�> 2�%�S���9���gi�.�� ��!v�!�, @^\��a��G���񀍮M;!�[5p��C'�]�'�V���OùzB!�'&t���TSo��)�и!!�� �|�b�K(5�Q��/XW��xҔ"O�I8ӯ�AҐ�ⴎ�6Z���"O��X5�^�;��q�%�+57�eJ�"O䄫��.PWN���.t%Dq"O��jD&�"�&R��$�"O��H���Y�HYW�ץ5:|Ò�'V��2=��`Sv)6W �	k�	��H�$B�I�D�ɠ#Jf��Ί+S�B�	�!���s���h҂$�B�V�r��C�ɿm�:Y̍ ޘ�c��Q� Lʣ?1���V2Y�%!$BY��4��0Ŋ�`�!��9��I�F,�m��JVC]�]!��͠4��HHsO1P]�|���J��	^��The��<t�q*J5�����'#D�0�嚉͒�`e��"HT�Qrj!D�y�dX�`��DHDf��*�+'�=D�0��◸)P0����61H�iG*?D��7eF&C{�@�:i���"D�0ر�^��3���//��D�#D�,��صJ�J𤤆�]%����"!�d$�O �0�%@������&Hc�d>LOF�#w��J��y(f�2i�N��"OR�f�����*D���"O(���jP��NP�.��k&�� �S�	K�����㝏���r�2C!�dێ`�6,�B�Q\�r��Ĩ��0!�$� �p���D>z(h�Ʃ�/j!� &\���E数Cg���Ǌ.d!��YF���は��do��C�gL�P!�֊�$�f���eq�E&%G!�DF�,�k��B �I;V�:wFb�	o�'��@äU�j�>�����(l���
�'��4+��)[����fJW�#�jD�ʓ$��=�	W�+���#U�Q�	�'�ў�|bCjG��: �K<Il��@v�D�<ywn�b�J�K�%N4r�|�%��H�<y$W�H,���{z(�-yGB�	�UOj�`�}:��Q�H�e��?I����.�΄rx^�8�Q��!�d��^$E�+؜k�ś�AL��!�D��uO�,��&/�5g���[�!�d�*�1@Zl.�A�v����O2@H�j�U�ZD ���%j�l͹"O����ǔwC؈���/�N�"O<e��-C�=������3r���"O�uJV)L
<b��$f }}.�x�"O�}ѧ瓧B��<9��c`��b7"OT3#K�u2�;��]�(^2��b"O��I��V�iQ,�s" �3�����"OVli5��tL�F��&y�V�Q"O���-V77Ѻ�3O��[ q "O`���`�~�
}P����D��y��'��,�RdR'���pPΉd�R�j-D��K�m��tL�Պd%�2=�"�%.D��P�
�:�L�d�͚9���K/D���);��yD�� $阦�2D����$֬]	���`�W�y���0D�L&K¹sH<!҇��>o�䓑�*D�챵��l�Dj�'Ѕe�FE�fn)D��0vn�53H��Q��;YDDY���(D��e�N�<�(i���Qb\R��1D��jf�Ʒ'�|���m�A���/D�K�$�!l�s%��/|��h*B�.D����Ǫq�����N�LՌ�P��!D�� DhC�"1x�Y��/q۬]!�"On퀂�عBׂ���D�>�� 6�|�V�h��S�~<����#IY�4��a��A5�C�ɜd1�7�O��詢$�%�C��LE"�1��$�x�i�iީU�B��(�U�V�\�a�����(���B�	�*I���HםQ���P��{��B�	=u(da��[[��(`����B�	
V�~����˔
}�`A�J�DڔB�	4�r���l����z1MA	h�����	�Q>��uC��A}j�x��P~��B�I%rf<`���5$5Q�?q��C�I5�r��c
>h�
	ؕ&_ �xC䉭)�F�qLX3uc�0����5ybC��+!�����W[��PO�1C�		zb� ��lB"��6(�	B|
C�I"��
s�	
�f�@��XJ�B�	u�ع��
RI��M�IQ�5xC�	�nY�+3�A8t�^	"BE�{�C�	ɩ5�9a��4��.H�S�.C��7r�����͙M��GO�U��B�I�M�b���@+.0P"1'_�B�I/J�NlHBц^Ϯli�.M9��|F{J?��
�R|��`�.
�ÈP�f�>D�����[��`�"B����"��&�;D�pУ(C�Q����Nŀ7��S��8D��Q��@���Q�*��k���b�+D�4AFƐ?a�p��s�c�!$D��"��*��RR
_�5��%))"4�Haw'�VW�b0���������DD{��)p�`B`���e"w��,x�ڹ��'D�d�vo�_��bE�:d}��J��$D�P���<0*SF�}C�rDI#D�h!	R�*ֈA���� ���5c;D���"NL��jK(	<�I��/:D���#j�Ot�U�'H�/S��U1p�6D���r�²tXk�n9��M�T�(D��S�'��Qi�K'���iG8��d'D���nC�7sVA�b�H2�T9D����\+U�M��D��c 8D��c"Ԇ1���4�Q0��X2�!D��B����+8�i91h��wȆİa.>D��8�G�kW&���,�i*'�;D���qk�#�|8��Ԩ{2�c@�7D���3# �Q��"�֬x�E2D��B�F�RW���V�Lx���0(4D�ȨBI9@������&0:֐��4D����`ו'ð�P��M%����.D����/4A ��X 	�,��K'D��ڇ���,i�h�s
W�_��PB�%D�X;�`y�j�S���A�l|�@�=D�����f�Y�7�k� ���7D�`�AI�p��1g�W8ZT��;q�'D�غ�)�(F(�,Sӆս*�(8ƅ/D��[�'C>Mx��r%M�<��T1�b#D�ȋ����⨉��8�� �bL?D�;"��W�&y�2+�\y�i�c<D�h�!�ɴ{3�]jw��Xi��#ï;D�r��9`�(��\m��H��9D�l����`�c�.P�BQN�M6D�p��fݔI�H�U�Ln���b�4D�D�S�BR�q����o�x��4�/D�FH_(��	8�
�Q�z��8D� Xfj*Q�����0��!E�5D�� $ū����Nz���"C��&�T"Oļ ��"5q��� J��~�"OPeq̒yd����RZ�N]y�"O���f�*�J�%͋�k$PmB�"O@���*�V� �K�'A���t"O)��\�@�޼Y�IZ�m<�DJ�"O��B&�[}*��ǿt8�y�"O,��V!ǅp���@Wn4�6"O��
��?�J� �o�j�e"O��5���T�$M�Bn�?
(5��"O�`��2z��Ԡ�M[��[�"OrY� �Y�:��㔁��a��"O�jW����u�dkJ�#^*|H2"O����En��c�o�x�S"O)�S��H8; $R2�&�;�"O�}�"͇�Y����6cݜY7N���"Oh��eK;#�z���"�-yF�:"Oވ91C�7cP.��D����@� "O6U��`�,"b�l	")� M��l�"O�� &�E��AP��6,�> �"OF� �_4Z�4x�� � ��c�"O��:#I�Mײ����"���e"O��#�R�G��%@b��?||�Aj�"OԬc��F�n��g[�L��HB�"O�X���.��{�G�s���f"Ol���ǡo+�E��  c�x�"OȘ�C�tE���&ѴU���c"Of�ȁ��+UX�2% %�	w"OT���ș�`��de��4�4"O܅B�d��7gX����	�B��"O<MIv����ċsE�0l ْb"OB�� ���4^�Y`p�)U�>��g"O~ (G���X{����ă��d%r&"O�d#�j��-�]����)��|ɣ"ODY;�2d������;��E�"O��Tϥ<�xP1� ���HT"O��� �V�>�#"��M����a"O��"�n!!$ô���#��p@�"Op�
�A���h @�i�4X�6-�o�<�a, %�0\��+��${�)BE�<�1�8Z���e�B�1^D�ʠE�<�� �, �t���$�&���j�nD�<y`	 >��	u戮R}d1�M�J�<I��Ԡv��
,�n!K �`�<��)]�:�x��3!�: ъE�F�<1�W6Ph#��8����m�N�<i¢�Q h���@�C�r�h�H^L�<���&��i�.S��иA	AJ�<Y�`� � �ѐg��@C�(Q�N�^�<	"�G�A�c�&��S��a'[W�<Ad�[�Ba6H��ȵ�� ��DM�<���S�N9X�y�� .��e�v&�H�<qd�ͷ<�Ö�&�k�N�<�sG لqQ$l&+��ʰ��F�<�A�P�b��Ea^IY�p����/B!�D \���d�9@��3"��!��ޣ%�6p�f�>*>�)�fօB!����`�6.(�Zg�D�a�!�$\�<�帠o��j����Hf!��P�-J��(�Sx�D�d��;UW!�� 
�@��ِ	��Pb��P�\�!�^�; �u��D��,ٲ���Oz!�* ��)�C������4Ӛ�!򄔭��Q�O�,-@��ۄr#�C�)� $�KAڻ/��Q�<(��$"O�]20W��bU`N�)�	�"O$I�녜&�Ѣ�G,JE��"Oly{ �ħx�& "V��k�tx#"O����U�>��"�?w9Z��""O�M{�j0a���ǇǠ}4� ��"O^QI`OE�5@� ��k�-r�"O.86A�1>=0�ɣ%"�ؠ�"OX<J�I���F$��.� IS�"O*�`b�ɸf �H%Dح,�4;w"O^j�'�%���1���3}n� �"O���`Y'Ak������teb�8�"O���0l�*����j %bLA�a"O�`-�<x"��7I�h%��"O@�Q�X�eq�a�Ɖ'=�AS"O���!��¡�wϑ�s΅��"O�tR68}ȝ��#�;l�T�5"O�:Nr�T�N�B���J��y�)�_bj���K���rσ'�y2�/����jR�}&�	�0�Q�yR�Q671Y����K��`&?�y�m�MxΔA'A��E�~=q�5�y2b~��=��&�=CR��N��y�,!$c����m
+��PZ��	
�yB���̙&�^uG`�	��?�yl�T���iP�W�ZX�2���y��¦�$�����}��1
ѧ��y��I�,�R�@QF��q ����Z��y���
DS�����J�k�V��Gf��y���!%�ɩ�h�f=&l;� ��yr�H�
�=�7��>^�t���H��y�j�,ˮ�zb��^Tzf��6�yr��:f�ŠVD�V6@@�/���y�$	t�. ���8LP��"F���yƖ4^	@�إ��ѪIGpD��'�h�:UFR8�I��`FI.f�p	�'�n�*���6��	���	)H0��'r�!ۆ�H:g�V諱D� r�p�Y	�'dF�2UϞ:d�ޑ1`��b��Q
�'�<�B`J�Y���bT�m����
�'yT��U�ɘ	*�E�a%�/;���3
�'�h�nR�T���F�@a�`�	�'��Iv��>q�$�q�'61?�D��'�BH�w�U�-�Р��ΰ. D��':-�F��n�V�k�τ1(�"��'�.t�#D۾����K������'�> :Ņ�uƴAu�IX����'�r��f�C/�ĩu&B�VnF1	�'fn���1f��l"q-��I^VL��'^Xrk��.]��\0Pc4�'�����hg�qb��F��Ia�'����d+�2J�h��W�\�M>j�'��8�HY��@%Q���6����'�8�W꒝0B� 0-��1�:�'p^�3A�Ց0��ɲ�_�%��	�'������ɖE�RqүH.,$����'*n,	g�е@�V�a����r�pP��'���H7��1s⌝����$�����'�$���0E��03"l�#X<q�'�8M;w��V��Hv"��(��1��' F�4cs��ē��B��	�'���ˆ�N4%�5ڱ,��\�	�'�.�!B��� M��ƛ� �]�	�'/n�� ��-<j ��ҸK��D8
��� ��1k�L���ʕxw ��%"O�����?y�h�J���nEh��"Ol|Zf��,��!��Hb�W"O���$���/��jœ�w���d"O�\�"N	�R���cU�W��V!b�"Oi�/ؼl��lQ6F����"O��C����FB���fKZ�Yc�"O��� ��;s��X1c*˛Pd��"O�Mz�c�>Z�.��JF  ��{�"OfM �ϙ��N=���SN�2U"O&�DڪY�z�Ѕh� +�0�B"O�@
U��x����*\����t"O���&�^�+^x�A!�*�ِ"O �	��سb���Iv��&pz��z"O*(@��_�_�)f�W`o�A�Q"O8 ���}Y ��E��(��Y�"O\0�Ӭ�k���Ҕ�M��[�"OP�xD/�N<<�t"�`O�@P�"O�8 E�-�Ȉh���%�&��"OH�Ц�dm���v� 1�P��$"O>� ��Q3ܸ�u�M� �h���"O��!��Fd��	
�5�f�[U"Oh�[w���
�J�FK7V��i+U"Ov��� ��ơ��G�J��S"O`}@�k\2*5+�E�=Z�ɣ�"O�9�A�*$�r�� .�4qPR"O$rAE�2,"4(�'����p"O^`yǎ�C:����٦SR��P"O vg�/'��1�ŏ/����"O�U��R*^rR�0 ��	S"O�Q��:�1�V�/!�N��"O�p��2���хB�ppS3"O����A�j������Z�cTa��"O�Ъu��6r!�r�A�MN�#�"Oĕ���ŏg߂�0֡C�e�X}c�"Ob0�#,)0~�����a�ڜ�"Oj�x'<��ʂF°xp�i�`"Ox�&�݈
�ĵ�+�gf����"O�j�JH!r�D�	i�4<c8�P�"OH���J�O^�{MP�9^���"O
��я#��5����=芕"O��J��W�f5\m��+��L�ܹB"O�1�O��&Gt]�P!E7x���"O�U#C�O�z�ȂU��(�T�C"O�2u�
W�R���}��ܢE"O2��bLL��
��‏��R�ha"O:IA�EP="����i�60e��2s"O�����4bp���]_��2�"O� C=n�P� ��AO5<q�&"Ox��G�#vzl`�k
2%� �""O�Ⱥg�!{�\�8�ꘞ2P���"O��3�ޝ0*�\�����\��"OJ��R�W�7�)TIP��@�j�"O��bu�߰|���z�X��"O�}�%�X�-��<��
�C��%�E"O
���!!��a��bH8q^�� "OJ�``lќm|�s$�F�Y�	y�"O�PGl���F�3� ý �:�#@"O*�zc��x����E�BG�80"Oj��Q�9�.�7�ЌD�B"O($Sf��� #���8�0q�Q"O=��BǕ)�<O�t��}Pe"Oh�3D�#8Tp���%?|m�%"O틆#�6���	��3�"O� �|�a�B(l.����	�" ��"O �q#ڱG�pYBG��S� �)$"O�H��?WV��t$ݔ@�|X�"O&ݙF���*]`3��eE���"O�pha���9yX� f^7X�l10"O�5R��Ј5���0EN?�$�1�"O�P#R���n� ���6��)"O�CS �>`�fK3�ɷ)��x�`"O0�Q���H�6��G��W�q%"O������G��r}�|���B��yb��2,T0kpc�D�QA�lY�y�?~YN��3��&hY��KX��yP�QT^�I���uL�t��J�4�y���7^�z̍fT��K�y���-��"V`	c��h�m��y"kD\���9����b稱�eB�y���B�$'�XEHL�E�S��y�B;dđx0lN�J*HA����y�ˑXh�+A$Ï?�jT���y�#�9I�Z��#��&B\
��H��'" F�"ov}�V��3g�X��'�D�+��6r��(��[�a����'�&)9@+^y�е{�GLf�]��'6|���
,vt�z�#�����
�'���(ׅ�P����9�� !�'�Y;��Kj���Ӓ�F�+���K�'����b/~�H1#�)�5 a��s�'� ��`NZ'^�!a���,.`x
�'tVQ�`��*��]�8tHl�*
�'PD���߷?�Rh��
�zWN���'�ly����b��C����@K	�'�����O����Kv�I�x�nEx�'�Ha��C'Ө���X"rblQ�
�'���*�/�UDР,B�x���
�'����Q�0M�,@.�|�� I�'���p#ŅE�D��G�J#t���0�'PHⳋ�8&�&a�W��b�����'�
0��b��,x���I��h	�'�}Y��ͪ&��d��s�L�)
�'������6 @r@c�qG���	�'�R����=
d�-��
�>!��'�1p��;�ll �R%�H��'���。y��ܛ��� n�\��'���@D��E����iM�x����'��F�݈L�hkwm�m�@�x	�'ބ��VK_�CY��yv�>q�B�C	�'������4LB,�DU��X"Ox*¬?#�`H��A�bb"Ot�{�/�҈��'��UZq"O�a��A�*�HǦɱI����$"Ol<��� s[���bOɣv���B"O����`�5!�0�%N�9<!��"OX=*PNGN���띧W�L��U"O�!�aLG�N�lp��@�l�Q�'"O,TP��_�Y
�����)�J�*$"O�H��.Μ7o 9JaA^�����"O��jF6$r�;�ϟ6	��y��"O�8�FI5h� �[Ce�%t|��p�"O���%������0Ik��"O�Ak�I�WB�<(�IL+Wرcf"Ol���͗0l��ay�bӧVP�"�"O`AD������	!��D���"O�+[�@�K�%o���W"O6q�ѱ"n���ʘ=g�l���"O� �ҡ�T���F�Y�Mj��"Oz$*�@A� ��q�$$��"O��i ���Ur��ʜ)>�2�"O����-G����[���"Ob�c4!I3F�lkE:GN�xr"O�dYR����|�cP��|;�I g"O�L)Q�Ԕb�Z*Uf��-�`"O��HPa��,�h����#`51�"O0ݫ-�5]l�p ��J G���"ON�ҖEֻkJ��b[� q��G��y��X
&+�,Rn�R���h��yB�ڪ!��@�X/R�"��c���y2#����τL��mA����y��Y�P��Q�΄@	��t���y��+*�>]Y��%K*B���_��y2%��k��x��"��R�L(r#����yR��6v��qĀ\.4R��E�M��y��Q�
*!�蝎|�Dp�c�1�yҫ��1�j%��ȯp>�t�S�Y1�yr'��m����%���a��+�>�yr�ƹL�"��NT�Z�����=�y�F4"zX�x�C�2W4�l�@m�y" ��kR����JCHբ6���y"�L�)���� �)E�
i��k�y�!/h�(�a��@�J ��ش�+�y�	Ԝx�?;�|�d���y"H�(GLU�Ö0�bx�T*���y��^��5��N�+N`c#&Pn�<AïW&o��8`T�>�Ti ��M�<�3ڍy_��GF�Q�r�1�*J�<	�`��Pu������H��Iq$�}�<��lFSʼ�V �t<�q�D�m�<ْ��+ �VQ��/�Խ Ņ�^�<Q�@_X��հ�ê_�e��l�]�<a�蜕/n9�O��]��0��[�<�,��Y�|�R ���>�ْo�<eaN&�(�!�
>�̫q�@c�<A���E4�]1�ڃ><�xC$T�<i�ߧ0�}J�N��j`�ea�d�<Q�K>\#�S��3qn�I�X�<��=kR�uKS%B�,�z%�MQ�<��,�3$��mF���h2b�
M�<Q1,̴c�����
�q*B6��S�<1R�ѝW��2�e[��$ήWܤC�I�.�\�iDx�:��@���C�I2Nz����A��6dv�Zco�,HZB��8M­p&)� �P`��q8B�	��eK1�ZY1�)��#]�q;B�I�k\Z0/@��b`{5%�'�C�ɴCs�f��}�U��lݯG<�B�I�A2�9�g�(�*hRS��=u��B�Ix����̜D,$@�Da�E�B��3sb |�c�[ u�M�T(؍r�C�	��gE�j��I����&�C��.M�8��0�N�@�D����F�hB�80qh�	4&ƚ}b����=%G�C��.[�� �/C���F�5��C�ɕqU�y�Le ���cE� � B�=u��i`����B�<�#c&�:*��C䉠t�ʨ@W�בV����+I�|B�	r��+��C��J}�ui#`B�I& �D���ɼj:z! F c*B�� �^����$Kݲ����
;n~dC�I�?��=
&�=j2�4�V/<)�HC�)� T9�	����T#�l$�s"O$B7c�2}t0��BC�#xW����"Ov 8$M���#c��JI�50d"O�Qi�
z�6А� ��gH�ę!"O�m�"�35��Z�A!G�#"Ohã߇0Y�Q�%f �);���"O
��p�Ȫ/'x��Ve�w�,�QD�'��d6d�=��W- ?�d"��L�SF!�J�Fh|��c�^�^:" 0�!4On�=E�aҸ!���Qk]�}�Xٲp ��yb��,zrD�$�(wc�dr.:���>�O��"7h�!z�lĊ��_���0�'T���&N8�n�9<��5joD?I!�D�+S����ŬT��.�mY:,!�d��d���d�J{n�[��C��hO� )I�m�:��#�?d�eK�"Onx%8�ȡ�5�م.��9��$,lO�xQ ��	�L��5�>$"O4�H�
K+@��(�D�j��݃4"O�+K�6p ��&cE=��J��'�\�dQ��T�5-t�z���2lO����V9a���S�A=����h+���S����d�%l�\Ls�)�"(ZjY	��!0�O�=��j!�D�D�=e��'�J�!&< riXZh<q�`��F�|yFG�[x�#�Gmx� �'���{�4#Q�F�C@��dݚ^�C䉛�E���ۑ#�:H*�BW�Z��C�I2���s�Z�~y���B�L� �����X�t��h%����r@�*Z>!��"]p���I��ZKP�w�K �'=ў�>=ZDM��z�\��愺VB̄�5ʔt�<����t���V����5bTg���'���p!c��VҔ�C ���7�D��e�<D�$���K�3���)�զ|l"�zH-D���2��>\��T��"G�F-�$"*��1�y��i�"��Z!m7��-���K�'l!�dɷ#�zڡ`K55�Y�tn(�!�	��RS�$]��a5.�?M!��Z�<��PN
��$�n�/{/!��A�+f��@Gc�~u����͝�/!��T��A�F�W�$̠��R�!��X�2(>+��P�Q�<��f�ȿ~��yb�;6���Qc#��8�d��@�12��C�	�(.t��'Z(��2@��kª�O�=�}ZWD�G�:y��6`ڔɳT�]i�<	#�
<8T��pO��C_�0pF�j���=�B"�B)sq��	9/���C�c�<��� ��,��E�	V\9�%Ǔܟ,���$QyV.�;IX�s0�,8 a��?��a`�5f��A��qE~���`��1 $��*�{eGTm�����Y�F����	Z�E�
��WN�)�����Mc�.�^�d�@��/~lH�J�`�I;0Q��>��(]�8��iABW����ۃH!ONb��ɹQ�L�a�h"�~�+��B��9r���Gy+G<�J����� ��c��׶���HO���< �	��[q��1gn��f�t:�A)D��g!�d,�E�Y�k�H��',O\m�~�>D��Xs��=_ ��P�,�=[�L��<9
ߓ[SzDJaK�/r��B�\4X^J�$��A��4�,1��C4(�Q�T�V Z�0B䉣[���p�,=����G�$���?1�Ig~�`��8��&�3.R ��F���?��n����k�&z?��#�ʀ9 � "O� .	��#T�69��C�GPk���1�	�P��>��wh�9
p�	1 ��	�`�k0D�t�a)µ.�؊��	����6A�<����Ӹ+��a飄�% j�q���یUSlC��#4s��+��ѩ;�����a�P7�#�S��Mk�H�I�>���гM0Nܺ��Of��'�S�'90�F�e̩��U)zҸ���4���ʕ�E�֤���(-� ���u̓[$�=�R@ÆDӼ}��ܤQ��L��*jڵ"�g_D*x���8(^�&�|E{���oK�D� ��䞾c� 0i��yr���:h���d�׋Ym���F�̲��'�az"��a=ƍb��A�:�q��С�y� �n�4� ��}}�d:�B5�ybI0�>,�G�Rrs��H�#��HOޣ=�O}4-�Qf�+������3�R���'H���0䒞E��)\&,M�=	�'�<�¡Ɨ��=���_x�8;�'%��˓�Z�*��Fn�<��ы�O���d��7�Ј�6��'��I)�C��Ug!�Dٱ	%��zG�V���l"a!�dJ�m�8'"C\��1�֋D?S!�>?�ne8e�œ�H5�p�[�!F!�$A-P	��&��w� P�BN ~�!���eS���a�7q7��a�.'!�]rv  s��M/�J}	���1�O ���/z�����6[_���e�!�d��KN����#P��85�R�!�$�3GgF1K�̈�eL�XJ��z�!�ԅf�P�����v>-�b���"!�$ól75�낻w������=ma}r�>��)&����բ�K����t�W�<�Ɂ�~QP��.:x1it�T�'��F{��n���4���o��XOF�zu"O�YIV$ڜ%�f1[� *LZEh"O�U�&ܯyt�r��s,�z�"O �� �Z��-�0��M!��"O�3`ܙ;�1B�O*l�%"O�jqDŶ,����e�ܝ}�P�J�"O�`s�L�>xbm)�F
�E��Ò�@���	�U��A¥OuR�x�LχC!��,y���Br	��6l[�L��=E��'@$i*@�{��u��@I
Q��}��'a�}�D�Q�^h�ipr�3n���'�p�C�k zDűA��;#�5#�'ɨYFa��;�U��/R�:�a��'/�!�QF�*�	�$&�83.b�!�b�>qI<a���'�uPSHW$Wk�u�� ��l��y��'�O1��4��d��
dq@�'�<���=|ON���CX����/ʰ%ZF+�S��|��'���M���HbWd�~����'�
��q��5o��qBw�L���	y�O�$#<��+��h$�l�����%YC�<�4.�!J^t�x�@أ <�K��@�<�fm(sK����
�4�P�C��y�<�g�ҎKR��5��0;d	P6�l�<p����aáE�l(�!J�`8��$�P�
o͂��PM�7T�$a�W,-$�p��%t-@'�X�'���`m��(OT�=�O���� �
.M״Pņͽ5�9�
�'E�#��Q�8�X��Q}�m�
�'Bb�MW�y��؋�FąLU �8
�'�\U�Ҩ�4:RT�a��M������'�H]���[�p������a��� �uQs��0Y����
ʟe�s�"O�[��H�r�.Q��韊V�t�2"O*�8W#�*u���ʄ�7q̭��"Oƕ���d�"]x������u�s"O�-��U50fD�x K[�n��"O�]H��9_�B����9`6��*OP���ρ��pP%!4��
�'ȰP�e����G�՜��LH	�'v0��I�
�4$1�n	53K�,P�'TX<�B�!�8�ԓs��3
�'Ǝd"�a�
��i#m�$:r�9H	�'D�Sq�(X��ybrh\�+��p�'���Z�@O/$jH�K�#V�'n���'�v��O���h�ۃ���8�'��0nF�^�R6cU,����'x���dȊ6[�8��E�ڤ`�'�̙E�P
&��|���9q�$(�'w�x��� 2k�@�.���	�'���Z�̀+z� ՛��4 �1�'���e�G�<�����˸bX%"	�'Ofi%�=Ԕ�	A }y�]C�'������o$0���ؾE�X�
�'��Q��ם����T'؁u6.�Y�'�H��b�'.�t�r�`ŖKb��'�^m�f׼dC��y���Aˢ�J�'���{���:�����8E���b�'U~(#���f�1d閺?ߞA	�'g|�!@	�8X4`�0��I-/$��'Ora�箍��蕘���1'����'冔S�N�`���D��vyS�' �5��ة�f�Z"�?��8��'� �F
Й5Q�-���/� P��'�E�7�7�D-�q�Q,�b�B�'�X���bC����wG�� �>��'�r��Ad�4Z��w
��$B�'��@��D$ත�yb���'b�������k�l�rh�~MnpA�'/D�� �P��qS�(/v��%��'�v�q]'U�Z�` ES�f�^t�	�']
إ�:0R�����]��9	�'s`8d�� (�� A\�P-4Պ��ty��#��5Ǵ(�tO�u��d�*�u�lu�ȓa�N�q&�A=]s&��K�2�ȓ�t|� -�.����� 豇ȓ1rAa�CB�� ��D��v�"���`wҹ�஘ ��l�2U<m�؄�r�pcX�`K8��H9.L���_� tc��НFB�5��١=��ІȓH6�8�!��:VTi7�4uP����!�t<�d�JܬI�k�l�Bl�ȓm���"�A�l^\���Ð�9g�����m�F �7j6.�M) ����t�q2�<<j���
����ȓ,�\�I��4�F����Ue�2 ��Vg�+�6*�J��&���Jm�ȓO&����M[(&y�l9#�]�Y��фȓ8�Ҩ(�C&;��)�2��d����ȓ{�f\Z���D���ռ~22��ȓKD�&��390鋗�Z;}B���h�řq��\aE��D�ȓs�� ��-_���K> ���ȓ�T�JfO�{����d5&��<��c��8���U36��K�/�,'�C�	�;�x�ju(E�d��p`U�x�DB�)� d�k�ɜ��|�Sg	� M~d&"OV�P���8Hu�䀖%r2I	W"O�����v��X%��o9�(�"OPp���H�lđ��� w�%�"O�����-[� ¡�34��XQ�"O��Ad(�SSd협�؝9�XY�r"O�d�tE�#�
	ڔ��=.�X�""O<�@����F���j`�ˋWyF0Y%"Oΐɢ'�7��h��~T$e/$!�dF�b�z�x�W7Y��Y�R���P�!�$U�"�^A����%�b��!K�a�!�H)I*"��uN92�ഹ��^c!�Ě$zʲ)�Tk����cV�9r!��+�X�*5�'G�`�Ҵ��fz!�I	߸ ��$vi��B&��;f!�@� X�l��qa��k0�.*Y!�$���mN�3��1m�%4!�$�%�R�Y��̜v?F]�Ṙ� !򄀡lM�щ�
ΌA��0�@@��O.!�$S�U��FGO�wc���ӯ	4z!�D-8�p "a�F���(���54�!���q�8���!�;Zk��Y҅N1Y�!�$�|���PS�)X%X�]!�Ć10���&�ĻL����2,!�d��Q�ْ�@�b���hÔ:�B�	$B�m�sH�ø�J�O1#�B��(7�M�C�Z�I�r}�#��ZC�D�4�wC�
+�t��1,;J��C創|�)��M�e�~q)�:�!��k���)�b
:"�lA#��A8!��ع^������ĵIc6�Y�W�k!���1����!�(x�d��'�0�!�$�t�.�³�P���a�Хj�!�F��a���J�'���3��K��!�۫=�M(4ꙏ]�`-��"ȓ�!��G� �h(���9-���aB+ńC�!��1+;�\ [7D���6��\�!�ރ^|�]s�!�v=vij�!��
1R�V���č�PJN9��S�au!�$I�*���j(��ev�C
�!��<e3���R���H�E�9�!���&r,<���ĺz$���Q}�!�D���P�Ё	�bs��*!���<4�ܨ��M�$6��CZ!��"_� )�lCT�Q�[*20�	�e���r�'by�6��}E0��U
�Q�	�`�VL�E�ڎ��A�T��M���ZFC��T�8��J�<Y�"�y�z,ׁ��>�l���H�;��b�4uS������2P��8;z�L�ܺ���aW"O6�Kb
�3o�x!B6k��HT�$�9&�)۶/�e����I1O�Q>7^�pKHM)� ��XBV�W�+<`*�$K��x���Zz>=+aDLd!���Q�=Z�0��GS�A�X�!�yi�I�aw�L9s�|Zw���*�$�3e!������X&,�
����h���=(�h!&'Vay8=ㅍΣB=~q�w���
u��
��S3_��(�׆~�<�O�#}� hƝ#��)��oߙ��ՙ�%�d̓�����%��
�r�ybݓX���9Q�:������(�4>ɚ�A$����Ѯkz�y#ɹ.axr ��5��I��ǧ\�`�Q��$	 2�	C�ɓa%l`��6�r]���)פ	:�9��
��9�T�6{����u�T��2hl�Q-Y�Z����g�L�����Æ�݀�AaE�xw���,L�_5lX�q�\�ّ/Ozŀ�%�bu�)6L��(��QTfR� �V��dC�*��qA����NmH�'ܧ�� ��I%�`��$JzU
Q(�pd��1B��L�T˓?ιi��4 ���PÂ�	����O�b��'��;���?g�|�8��	�
98(�@�ؾ�wfYP��&I��-�+=4��ʓ�*M�G Ǯu����Ó ��� ��m�t�CC�1**K)�<T`�v��81��$���!�q��9H��Y�K �� ���#Ĵ/Wr�`�T=�Nl��	�81��A9�J�+�(��ET��[ĨP���#q)�?�H8�E��@�m�K���N�;a(��d��p!$	7��-�8�"�F6�&���+<O�0�r@�2�2��s���t�0�%�tTi`G'�}aA�F1]�v�1�A�r|x�H���3BC�)��$?�����b$����˗�V�.�q`��N̓W�&�A��	u��i6YZ�vQ(u������'y���+�X��X�o����'�
1 �*�9/!�y����Lz,�Sh�<����9L��t��?�ZȠ@��.|�3Dʟ͘OȊD���
LH<��a�q�pUI�\�en�0+�'](������9���7�.)Is%�+>.�1`�_23�fl�Ш�7]*�����Oh�W�V3U22���l�59���@��')�  �N�t0�9�E,�"�<���ǟ�fuʕ��M��K��0�iS�Kq�i9&�i��	DlQ�Y����e�R�4��!sd6�	� ����G�`=�7� I=��SRG̐��4�؆H&�,BF�]�M��⚃�yR-<jM�U�ٜr�������g���ړ�Z���m52}>!C�lX?[y>��9��i�@%.�qj�KF/�NC�	>7gz�`5�Bz�j��lM�<�[#�V�" ���VQ?��9�l�����_�TJ������7,�~>�{R�J�L�ٷ�K�����H'c}��F�&r���an�O�|"����>�������c6b�ʽX�� k̓b�ȱx�΁)KV>e��>qɟ 8��M�p�Jdhħ[�s	
��R
OQȷ�	�m
�QCF�ɭ)X^�����,cϒ�f ��gq��'Ĕ#}�ep�����J?"�S4.l�6u��/I� ���B
QU
�  4���<�h��A0Ra{ү�� r6eRXQV����bC�[����d!.$�em��M��̇�G�`PS��/�jp��Q�<!j�o�ȹ2$�*P�4�;ņYv�{����n�$ �2#}
w�܁Y9r�)&I!H�h`�C�XH<1g@�z*��D ��HIt�ӞQR���"�IM �I�E&eEj��~r��0��0��*9� P�C�;�yr�Y!N�^p�C)u`5���	�'���l�:ԀBGV�zY��ir�		Z�=�E��n�գ�`+�����V�l�TH
bbaN�ժ��H3f1yf��:Z����D=R�����V=-��9w�_��APDF��j�G}��w]D���(_�S<(�hT�p�[+m�(�C�f��X����d;�ɫ7A X)E�(�0�EG��˓I]-�@CA�pҧ(���!��<I�L"��G�tl�B��4�S�~V4�����xB\i�G��*���O���@��}@8'?�p�3���@-B�2-\�f=��c�d6���Obe�
�"tsX��L��F����F�B�"���4��?Qg`���||���|��i�f*���)F|�,�>��殟`��r�v�x�L` A���.b ���$$�ɛ�t��1��5�4\�B�Ʋ�{���� �H�ҧ(���A�c�*���A����y
0"O��3W喭&�:]��ɕb����Ti:��I�`����t��*;&h�U�[�j.%j�K

M���dݺQ�g �B^۲*�8:r���훅�x�^��(0�I�!���`!���S���O@l��)�~[���aɏ�lft��'�� �l�UₐKФ:O��0A�t���I��1@��''v���L�xˤ�R�-,w�aӌ�$�OH�����mڦ��Ν;4o򨪱EȦ_��+ab�	B�!�ϋD�p�G	U��mHsA�	��������q.�B��y�,��:�l)x��Lw�.IB'�:�yRNJ^�ݺ4
ޑru~Јaσ��M�«���'���%��3�G)��2��\2��dw���'q|Mdc^Y�LA�� �2�4�?�	�sb �	�@�zU��ˠ����=D}2��x�}�桛��r�*Q�C:I!�d���x�<1a�a7\���bң:p"q;�(U{?�����&��e���ٱbwD���"�B�ɩ^���Ke�1O�$�ӆ>
j�B��,�,�Qm(5lM����\�*B�Ip����F�"��%B�Z �C�ɿ�@��V�^�.��jKA��C�)� da�q��=�D��Sh�(&"O�E�!\�,��,R�00nF"O|A!$��ռ]󵯀�A3��P�"O�G�#��l�2kL�X,���g"O�PI���U�a���W�d$��`"O���2��}L�<A�AI���D"O8�G�Q��H2� 9n�9��"O|�jT�� nV~�#�ǩy_�L��"O��J$�ڧ1����d�p�]�"O^�����4��ae"�o!� Y�"O ���Ć�͂L�҂^�k���{"Oܕ���	�y����%`A.B��X7"Oօ2(D'h�1�7��>��훗"O�3G
�7��[�/�=a#��&"O*�0�g��:,)I� �"OhB��Q��`��B#��h�"OP�1�Xt��]S�C�*�1p"O,�cE�]?���c?�Y�F"OpUP��ޞ-'��ّ!�9�5�'"O�0��G���u��.H�i�"O<Ћ��N@�#��cx��"O�٠�^�A���BA��<N����@"O<dS��Y6�:$�� �6<���z�"O�QH"�_�,�y�o�J|Vp5"O&����<�Ps�� �L(�d"O�,�0�y�N�"��A:��5�"O�6/�8��x&�ݘo�X�M:D�xAWgEQn�2w���5E� [��-D��`P�Xx���M�������$D�����,�����l���lps�f"D�D�B%�5�\q�t�P3r_�TP��?D��ȆT%[j��]?�h�Rf�=D����E��p���+��7?@$óI8D�8���'��a�CP7����cF;T�􈦤�=�(�^�/"�a��"O��0�L�77���M�7<,ly�u"O�i�CF>|��1�B�I��e"Or0�q��[��+��ƈ,e *�"O0i�E	u>���E3��]�U"O���4-]`[Z1�6͏ fH�""OR\he�VH��}�w��eD����"O�؈��C@���7&�>����7"O�h�A��ڰɧF��<��]�"OR�	#)Q"E�j��`�Nc��D�"OtD��HRvؽ�֭�)䨚�"O< �T��K�� 2�ö?�}b"O� ;sɔ!:�3D�ƍR��v"O
����ލE�
ԹkE�g�>��1"O0��#�2�y�e�ܖJ��d�Q"O����O�*0�6�a�̸�0�"OZE��HFwh  @�k��܀C"Od�`�U�h�R�!uΟ	�.h�p"OtCF-h���L������"O��h#gSN�P�!e�%Py��p"OR��R�*iC���.�5I�ލ��"O0	��j�)#l�ܣ�n	��͋"OvH�s��4����@ʘ�M�.���"OlIc\�d�P����JU��)C"O `��&ߕ<e�M"���(�{�"O���P' �>?��QF�En�̼��"O�}3�e�6Qx�ͩt�)q��<�$"O�M)���/B
�(6b��0�,0'"O��xΛ�_%z�� �n?p{"O�M�݇#f�a�&[�eK@�d"O� ����HϾr)���5b��"Oĝ
�Bn��	��#ڨU1�8y "O``��B0a�v��6c�!{[����"O��Y��1�`��<�|��"O\uX��}�,)��C�X�*�I�"O�rue�w������R��}�""O&� �cQ����d@ߪ{�B�r"O��)��!W���T�WB�h@"O��{��By���B����`��"O2����Y31�L��!�>`�"O��P6ꕷ4�DX����K�*T0�"Old0��J�%�z��q
�z�|C!"O���e�T�2�բ�Y�!���9�"O恰2i31�"�*P���u,���"O�!��ETU��53$c�"yzpQ`"O,�q�R�2��A$6�ô"O�1(��R�;q��GG^Y"O޸pr��)?0�H��m�B��l�<�C�E�8DDk��^�\�BjYj�< ��'�<bb����Pw�N^�<���7�p�6�NK�I8��U�<���%*��K�۷��k c_�<��¥\��a�d��&&i�e�D`�<$J�YbS��Pj��'@�<�c�"�NMj�hB��ۀNKy�<��݂.�<Y�`�.H�Gc�m�<a� } ��Q�J	k���d�j�<�QВ;���0� �bMR���x�<�g*�>_��z�Z�l�61���Q�<YO�Ts~�8�e'_� �+���D�<��C� x��M�f��[��G�<�c�V�[�u�@�F�t D��ERC�<iUn�9�LثW�܉�N����t�<9��ɳ#�X�c��H�f�E���w�<!0�]I�����0p��J�<��.�#f�l �m�o�L��fA�<�s�B,Q�0���
�1G ��4�YW�<C)�%Y�p�NR3~�xҁj�h�<Y�(P��p�H�-{$)�*NL�<���X*�$q1	E�*,��!FS�<���R(�f<h��'��q�t��k�<�1K^�F8`P`�,x���#��<D��h�C�\��:Ti�7Ӓm9��=D��0��O,_����'T>SLi:T@:D��e�F�F%J��S)ķa������;D�Dy%	��:��بT��Q�ԅ=D����K4d�8Xr˖8q�"���i$D���tbP�1���(�dS�g�z4#D���Dj�(v)XE��d����!�#D� �"i���pA8A�բ@k"D���lS)
RnE�WM�
�P�;q�'D�(2T��+ϲ=㲅��0$�"D����m�� �.����ǖ(=6İ�#D��P$�77w<\��V^�>����5�O\�pd�`���F�1F=��Q¯�9`���a�'��A`�N�W��uo�p���Y��d�IpP��ӈ-�Ӗa���H�AR������3����DN�`��� &�@$p�e�΋^И���)�c�
LWڗ�P�%�9}�SLW`4� E vtP\�`H�D5�#?�"#�)-
���b���&Ŝ�[���o�-X�)�(u H�kք��U�H����.=�=��![#|�U�@��-{<�Ɇ���m��|����B�/}2Ā�(g`P0��T�F��c��+]�T�Z!F&��(���gg΄cEk	�঑h��a���+XM��P��"E|�P��04k֥��T��;2�V4Y�ǟ�q�8�JT�A�I�F����:#܈;� �%��M	$`�
����L.l��E��A[nӊ@z�,����vX�Dr�q��h�!�a/��I��!�D*G㜱j���X3�Z��4lt@��b̟(QrP�	r�ƥSC���!�m�]��2��q:� ;�a�t�jV(��P��*D�s�h�5M��$����S-]�[ղ�ns�'"�je3�(�#k�L���dΚ�ʄh�a�7q� )�hԿ�x��1	�҄���<���С�)A�	�Po��q��A޿F* ����g��I�a����k��I%�ׯ-m>��%gӡ?p����+�O0��b�U\�؈C���3@���# �10d���iM9��9S��; r�'��C�4s�O�����C�EN��]�@a��	��8"0
X�#�z��"�
"��4�ӡX����(�M��g�M�����F��!��,<O
�R͈!\���1�9?��"5\��J�ԜB��$��ճ`�\�}�e*؁2B���E�D�d�DlaSh�PΰQʳ�6T���5�������G� ̠2��K*X?�Qy0�>Q55�gy,-/(D�&K�0��=j��^/�yb��u���� �ë�,���KիD�$�b����2�*�j��e��%�Y�(A7"2`��	;Z-p�ɇ���#g����
E���1,�*~�!�ݭ!̀z� �#ka���1���
1���	�$�Z�.�q�NV�(��N�3�"H�N̆}����$���y���y�P(���"Xa�-)��:+�ٹ`JP��=��O�QͧQ �<�dj�zB�YI+x�x�	���L����WHGSb��t�i��h�m�!������3y�0+�<ӢBq=�O8�;P�U�b6�� ��&Tp�[�DΡCX��`Z��H�^��☡s��q"V'+8u���"O(��oq�B݊aI�Jq�!R)d���A׊Tm�D#�g?Y��A�<;z5�e�Z�z leK�g�A�<�n�
��Q䇂a>��I��8��m�Ij4P0�'.1��M	��`�7���\$:A�x q��"B�w*7Y�a�¤�9��� w�ɡd�!�$M4X�N��W�0!��H

h��OYq�m�$��x�����<�@ܑ�d_#bN��F�E�!�>Ss:=�a�Y�sd�ZgF��;�l�EG��*g&��tg���p��ؓB��th$��`R�ȿ�!�d�Z��hAu���x1�T8O�T�DV���N�J�Ӕl%��gR\8���X�ab�4���;}���	8��ؗ��I�]c�!8@:T���:�΍�]�@S�aOx؟HB *N)�	HE�N?;�p�Y�2�!�4� �`�9���`���/�t`���`��_���"O$�3!.�D[­	�MB�"A�ܙ6T�d!�f�5%�9S�>E����\��H�0����녹�y�)���9RT$D�b����D���F�'�@�S�E�H �ϸ'o6颥�ֆ	��q��[,�r����>j8��u(�����o��K�d�� �)z��!� �+�O
`���6 hћ�N��{��1G�	�8��o�;��O���"�@>?F�ţƭV
����'�65�B)��P'L)vly�!+O@�`PE0nv^�J��|Z��[#�X�2�m�2&Q��P�@QW�<q�"N�iF.5Q�ϫ5�d��'�����5�l��w!K�g̓e��pz�Dý@���0���z1���Yy<m[R/	���X�*�"�Q��I�$��B�I"�l�	w�r?��Zpo�_�pB�	�^���@��T7jfp��\��tB䉀��D_�L�}�����.B�	&I�bC�!�c��V*[�pB�	�L층�2�[l�DS2 �'[�C��5Q`�����СH�Kr��C�Ɍt]��DO�t��
Ө?��C�� *#<�{�'Ĭq`��cȝ�N�B�_~m�҈A���S��X�,*B��pZ�&ݧ<���'��(�,B�	�G;�l�a�X�(QщN�2�C䉼.�yA����98%�6 C�C�IcA�%�d��69Fy�t��
�C��v���'�=�,��S�N�B�)� ]a7���$%h`�fg��WP����"Od�SAŉZD`�藇�kS��f"O�tK�)WR,��LM1!H�\K "ON8�Ѐ��l`���j�{��E�"O�U��l��oF�<����h����"O�!���.R���qt�@��ۇ"O�0If�*qA>��F�M�_��yg"O�l{Q�Ҥ)tA���B~kF�ѳ"OfL+��L��R&!�@�G[��y�&��/� �)��aIb��!��y���PX{#��*QԎ�3��^0�yb�q�n�F�šO�<�`�^��y�B�X*�ٖ��6ikb�����y¦� 	�I�7�ֳ?^�"g� ,�yr�_�����SA�^�̜���L��y�	9~���p�^G&�jE�ѵ�y�����5���"�0 �k\��y��I7逩 W���^m��R��y�B�y0����	<�<������y�aƸl���{U)�1-�5�y�HN�_@8@Q�<kZ,xҦ��y�e����ف��]r�̫�HG�yb'ֽk�T2�H��V��~�n\��'8,u��$��,L�`��qX$���')�5;EB/_6$�3/�l���	�'lJ��b�:I*ĩp�ڥY~]p	�'��9
vhR�}{�i�a�j�03�'�M��  `��]AW%W/o���J�'Z*)�l��? ~�)�&g�n���'��9��V6f>���&AߑT� �C�'2vd(U��
8���[��J��'�6`
e̝��ƹѰ#�9<�,�3
�']�=Y�	�`�q+ЂV�<�x��'0l ��ɏuu�͉w�D#0i�I��'3 ��9?��v���0oz��'_���0ѹz�:��d�T ��'��03u!_�C]PPE�ߨJ>�A��'�����+/\�H�T�B�NhS�'�L��'mO�6�����Ak�&m��'�����	{�v<bQ
d�f��'�X�bF��Pwv��3Gd�����'���c��!a3�\�'�\K��a�'��`��&��R��2�.U7C^�|��'
\h��#BJ	Z4�OjW�q��'�$s5&�
%ټ(�fcӮ��'C�H��{���ŋ8�� ��'��mZ�&{@�Fœ9'��i�'���k�#*�&}a�,p�'��tBFF.��v��u�$��	L����Fұ4@�F�G����L�7LI���ȓQs�\��E"0`Xv�| �M�ȓ*8BC��F*��t�!�]|\���qb��Y l�K���A�ȓlR<}!&Ţ{���H�|��Նȓ|�jIA�Ϫ��ɗH��|��\����~_� �b��?_��X�ȓ6�Р򧏕eO�yiGȍ=e��8F��S9���H�Һ�U��bB�#���}�c�5��O�R\�ON��Q3Ո������"|!^u�*OV��JN<���XM��|J��W����G��|IT�[2�AΟ�Pe�y,��ה>%?���4a*4IP
Ox��ç@G��@�)��@����g]=~�II>�꓇�(�P���ߺڞ����B�<}i�R� dy�ޒ�0|ca]����6/�9�r��� 2�K@���o�:����+���|�H~v.����a�ٟn2�����S8b�j1p ��)ۓ͆�l*/����� \���a���i�ǃ5��J�O�!mE�|0v��$~�I����ʧ;�zH{$�7I��%	�H�0p��+g�l���'T���Ԋf>	CoωH\|�%�)T�Γ0v���I-k���M��?��BӃM�bM`'+�,2F>��P�1��&W�-�ᓼ>0�M`R�C5M���{���g���O��[��-�)�+8F�Q�3�Ly�\$�TR��I�c`�؃���S.u+�q(�%�j�e{��	�/���r�b�0]�ɺ?Jh}a��7�g}�T9&fP�Z7��8B���q���s��#<�zV�λ��<���BR�5�`�C�e⬫��v
� �&���&Q�a	(��[�X � @�?�   �	  �  �     �(  ?2  =  %H  :S  _^  ti  �t  �  ˊ  ��   �  s�  ˰  ��  ݾ  ��  m�  ��  ��  8�  ~�  ��  �  O�  �  ' � � V �  '' �- 24 u: �@ �F SM �S �Y �` ,g m �w � �  ֖ ڝ � _� _� �  x�y�C˸��%�RhO5d��p��'l��ɶBy��@0�'�F��L��|�t���pd��46b�Z�4?NNqhs��|`I4jE�M�6��"-_�7RN�wk��uGjY�7���
/Y���F�6=b�l��wm�u5�@%=,ĥ�t�X*v�"@�#�0 ��'��O���]37�,����M3����U�̳��A#['�QrDM[Q��=�2�I5'�lÚ8+J��E�Ql�6�\<9I��d�O����O����.~� "G�zʤU ug�%w�����O�RP޺/�pʓ�y������?1e��RfL��篅�t@���ɮ�?������?)����'��$��fe��"�[�AߜXJ��[ !򄟤Y?P�����{ʠ�z��+K�J�"~d�CP��(e2LIcP?���=O9�)�7(X��yr�Є:���1h��(w�HBĭC��?���?���?����?y��?i̟����Q�T����H6&c�hz�'w87����M�ڴQe�I��M�i�6�|���WW&`�sK-n�h��AfىzN��Ї��j�4�rt&��,`�O��f���d-�.���Q0ϕv�Dʃ*��p���I\����҈iB�R�x�4uqNN�I�1�aD�<��2��h{�_�b�u9�1l>$F�\�L�|��� 10C`x���Ȋ�9�"�G{��	����D�ǢյO�t�t!ʌ��=	������oX!VW�=������<��)�?�M>�������`������j0����*U�<B䉵1x@YA���X#N(a��ԃ{/�C䉉"p�]6�ψ���e���0��C�I�_[.}"���̲̲�-�3t��ğ�B$�#����V��Ir��#;��N�F���^	�^T��↸6D�z�@�5���'>a~¥ܯp�xd�5k��9l	 `#3�y"����a咻�xc�&0N�C�I�C�L)�a�Q�Fr��2��FtTB�ɫ�E�P�	�$���J�?����x�����n�˳H�	���d�4���S蟈��d~��K�}�ɋ�l�H=T�0�y�藻g4^x���P�Lɰܪ���,�yRM�P��*�ꉅtİe3�b�*�yrF۲���(bJ�q�4��y$C�c��A".
�jdԂ������VG��(���:D퉲? |��ń�72f�1WV�|��֟H�I]�)�S� �Q�	Z����җグ �B�?e�P#яG�-��)�`��M�B䉬D3ĥp6��30*��9&葭��B��-P���KG��"ОѺ�+N�32�B䉆a~�AX4�T�H
s%�E���OV��>�� ^�Tl��'fR���[�~��S�C��l�8�ʹ]%[�����ͧ<C$����Ie�LK�Y���HH�[��¢;xH��I4=\X��0�	�Q���P Թt
�qq���!U����Dֆ��'���'\F��Ua��^LAPT'g:� �\���I|�S�O�p⢚�/5`�I��B��x��.�"�]�r�6�x&CK22F�q����3�?	,O.T����O�?�����˧l]
�$�d��P���lVޟ��I� =���3I+�)�'<�0�A.ǌ7|�|���Z�p����'-ܠ1��i�S�Oņ�u��
�.�q2��!.Py�OTU���'pr����� ��ݐ�%+Ntt����.[��'D"�'ݾX�AnŔe̐hq�(�m��$�F�O�8C��M��xQ,0}��Ի�{���ʌ��O���'���/
n��6��?!�>�Ӓ�ѻϸC�I�s�4�c"S-LzE�47��C�	�@�0��hS"�ᯚ�K3PB�I�7�
�� �&o�D҂ϓ�l�B�ɲ3Ӏl�P×	!Q�D���R���˓ ّ�"|�s�l�Ԅ��&T:a�#b��l���?y���?H>��Vi�����<������b��z�	�f�!�ݔ&��!���A+^���k��\�,���9�O�%��H�,N�`C�g�iK�U��mz��'l��'��)�<�,�<[,����`�"I����yb���+Q�	�a%��tV*5�6�X ����&�'m�	�1��	v���A
�Y��EL�ߎ-��$��?�L>����Ԥ���O� ~�{"Y�@o�IB��'$\)���'�4�[����O(�,8C#�<er�ѣ%F
2ax���?)��|�"��X��X����y�$�&��;�y�J�s�^���L�r���g�4��?���'����a!%0T���6��O��L>qAN���'���'<� �lQ�r9RU��K�7�xE�5�'��B_*̜a���o�8��\N	�鹢�O��S�M�䈙�	�<i��[�]�B�;n�s5H*&��pЯ���Π3���z�'�}J��Ѝbrp�(Â˧<�&�'�����~{�V�'�2��4�'�\��bH�}���Kr!�S��L��'���'��'���bF���g!�%7��Ę��d�g�O�TaBD�	A>�z�E�70w�(xf�iMP��b2!d����<�	k~�"I&H �� �ƅ+� ���XCvD�O���b��	:�1�1O���/�_�V1y�mO?=�f�z����	�J0a�)�3�e�` ��
-(�H%(�H��{,�D�O��Db�d��4�<���p��ױ����E�
?�ܐ��'#ҩ+���k�Z���a��-��`�,OP�EzR�O^�U�pI1O�/:�Ęi��`��}�t���\���4�?���?Y+O���O��Dϛz��U34 �*z+0�����38�x�	ċ@(SP˅��p>���;{�<��$��ޠ;�N�d:���Y�y�Ђ��	&g� E�&�A��uHu��EeRP���PG�)��������	��M�����O�㟜�)�e���j�^s,ѣ�Wx�<�6L�'����M �ޕ"�oJsyr�'�r6������'��)��>��D x�卢m�Ҵ[ei+� ��������Ov���O88P.շ$��勅��<PǕ�4`%h�"�N���i�z�`��mO:��{�뜼~�2y"�͖;�ԕ�k.u��HVZ}��,�e�'�&���?�Եi��i�OR�q���WT��$�7bn�	ٟ��?E�l̘<�z�H��H"9'�� ��M����?x��$���>z�Ƒ�q��N��|R�'�x����U�� M�hX�4
��lN���b�O��'�O$�p��o�0�F�L&~��Q�"O�1FA������d-;�|"O�0@��/Mx���,W�6>̼"O�љ��3p8��b��4�e*�����h�U��#1(<��ƭȺYY��'/���4�R�d�O��8�e��D�:hD�z���t@����<p�&��c��jѫ%]D���z!�a��+����}���!y$��ȓS�RI˲oD
%����C�!G��ȓ7�I��� �'�bt���U*+�≖'�`#=E��B��*^��8wF����Q3�+���g~,�D�O�Oq�<�B���.��Ze��2ffԅ@�"OH9�W�;�h�����*T�Mj"O���tnX��ҍ'=FVܻ�"O�=�wC��M�Y�D܌}&��k�"Otx ��MT��&�՟uxh� �|�K*�E�J���=��`#yZEs����0fj,��W��֟���O�����>Jh�Z$Ky�uc"O�]T�_�T�b8�Ã�{��!Zr"O�h*�e�!"F�T�Q�dw�4�u"O�LgIB�wa�Q���-][�L��'� �$��+Q�%�2(K~M@!�=Uuў(rP5�'(P�\ۧd�:[#�c��Z�S���A���?1�pj �ST�m�fp��h�!K$樄ȓ"k4ɐ���&6rx�@��H!���ȓA�vݪ��Y�4�H`�S�Vf�m�ȓ/֬�텶,�.xР(*�PD�/4�'q�J�k2�e��B��r%�O��+B�i>%�Iޟ0�'Y��{��w�B�PCh� BhD(0�'��ase�&H�>)᢯GK28S�'�~x�3�
C<d�7�T-� �p
�'����nȁ^t��F���J��	�'��s�43'
IR���iV�*O2aGz��	�{��d�ͺ|u���M
z;�I�I��Iԟ�$��>5D��S�^��D� 7�8,�T�$D�� $��l�8�0���^�ur�"Oxh �
fڅ�.O dct�i�"O$�@Ch�%\�H���MD,jP���t"O��`�/D��u8veX"/dd��|��'�h�L���g^��s'�*,HNZR��^����~�Iğ���O�PyfCKB�h@�3l�%����"O��Z���HR��,|g���"O��	w�N�I� A���įwg�0 �"Ot,�
-s����Շ�jTHH"��'���Dφt�������uTX�J��L�A�ўD)D�"�'r��RJV���ɀ̓3�@DR��?��C؂P!e�B�xl������.׈8�ȓ2"����͐"?�R�x�����ȓ�T� B� �x���e�#b|�Q�ȓ|�i0t��__�����ʥ{���ER./ڧ`/nM@ ��9�9(@
�Jo�8�	�{=�"<�'�?q���Y)i��r�V�0��2צ͏y.!�{�>��(�!�80!6&O85-!���h4����[�]�\<��.�)'!�L�C�H�B�K
,�t�b�O��n!�d�8�@y1�Z�<�6�`��Xs.�	�HOQ>�j���Q��`s�(^	Kԭ���<�t"�?Q���S�'"��Պ��H85�@����`ppC�)��	��b��>��`[�*[:��B�I�F+^Q�5b�n^��z�����
C䉒4�k����jf�,h�ņ�C� ?�5�p�4�dE���7�1O��F~"ĵ�~�D��D�(M�e�ý$�sc%�?�L>y�����IJ���B��5l1�G/K�B)�B�Ɉq��g酌U�}!��^G�B�IV�����-�����	�A�~B�	�<�Z�#��͟LF
��t��o� ����ş�Iu!ȃ#ü��D� *V�2V�1ړ9���G�$ڥ2{&)����k���b� �6k���'Na~r.ȧIc Y���A5�a��&���yr*Z�����:Ѱ�X$*�yR�S�hi#��o)`�k "e�ڼ�ȓ*��`
2���[��`��Z !OJ�Fr�7ڧw6\z�n_���0�Ȁ 5�r��	("<�'�?1�����$K�h�T�ʒ:��&iM'7!�ġq��!��?���mՌ:!�$G�p�f `� �� �+v0e�!���U�P�ր� Z��A���4nN!�Dˁo�p]�c���nt�(�W	ύP�I��HOQ>�i��<b�e+ro�k?��b�<a`B�?�����Sܧ\�e�F�J�\��E 2'�����ȓu�Z���M�Q,����!��J2V����<���B�>ĸi{� �U��m�ȓq�j�`��?)������*G�Ԇ�7/R�1���-<E�D
SzA%�����Z?VB��݋wߢ�������iu��~��|b�'���O.8 ��Ä<���+ba=zN�@�ȓ��Z%��$=���-������m>��y�"
�+�.�괢�5h/�ȓ`�j�i��� ��阮@��]��	*�?����1m�}ؗ$ ��T�0��J�'Վ[��ɘeۺl�c�̃0��(y�f\�@N$���O�����'����H7[��#�mER!�S݆x��܅Sy�m+�I�j�!�3���26OS(��H�!/�!�D��Jm�a�U�D�c+�4
�џ$Њ�I�[���iD�P,4�Z-��J�_�"�&�O��O��d7?q��Wq���&dM(O�m�F�Cl�<�.
5]^�	cѪݬq6���a�<� D�r �M �)H�i'Rv6��S"OT-I����y���ϢM[P�P�"OJ0q��	&n֥k䍁�5KH��Z�������G�$s!�Q(@k��W�K=:˓9^�P
��?iL>�}C�N9Q� �,�ڜ2CkP ~�j=���� �oª��H�F�l:�t��\Ҝm�"[�"�|�pWL=+�Y�ȓ=��XJ_�P�BE	�7bzpPQ� =D��Mc)�p� �dd��荹G��'�#?�)\?�ņ�3vuBo��B�t���x'����w�g���/���&!�ҀTb0C/�!���_�p�x5$�DD\���%3�!��=�đTg�h��D��+|�!�M�K���0U+��#�����`�8\����OZ�7C������W�M�A�8��v�	iz"~�Q��V(�4C��g�FH�+��?i��0?�e`��- �����E�L\jؑҢWc�<��B�2Uۥ��0SF X���]�<�T,ۻ~�.�R�Q1h2���\�<�`dA$g^�R���*.��("�X�'nb�}�D&^t��ץ�RZfx�Țٟ�7��|��?��O:M�����NQ����"\�4"O�0Z*�Wc�8xsK"O���#�"O��R�V-D~�tf昰p��R�"O�uJg�^�qo��٥nQ�X���"O���O?1����F��\x�R��+����/a>���c�CN�֨(5��4@�p��4Q���?�I>�}��`Vd1�@�6���'�x�<)b�
 8�x�r��v,R#LN�<��%A-.�l!�ܰo1h9	��_�<YfԢ`�lE��n�#x@�X�k�S�<�0��j]�d� G���4��1C�M�I��Oc��O��	�	�^ʈ�F$�j}�{$�'��'|"��>I�`^1<R>����P$�l�"�K�<�-<y�����BI�l���C�<yE�D��]
�E�$-e���U�<1�׮VM���h� ,�05qգM��,��<��DPdiʐc�p8��@2r@�E{b�� ƈ� ���C˼KKP�!(��W�N �r��Ot�'�OL�H7��I��	!j"��"O�m��Gt�`H��FN�k;��*�"OJ���6
U��dR�O�N�W"OD`ڢ��Ʈ�!$$S+g�[�I��h�<ԀeL�j0X���Bړ(^ْ�'�8�S��4�b�$�O��7hdAL�6A�����:�b���)6�Ke��Z�� 
�"SZ�ȓ��%��o,�V<Z�F2)�j��R��U�3�ʁg��ةL�Z�6a��Yʺ��p�Y��ԙ%ǄJ����'��#=E�D�!R�i"0�ޯ]�����T���d�@t���OƓOq�6X��"��AifHN%Ѧ!��"O��7l��p&��[`�AS�"O:�s�'�ly�@�����*C�sP"O*x3�˴'3n�R�j�w�f\ d"O�öd�xs��q$H%O(q�|��7�k��0�-�ĩC� �U�h�Y���=8�h��~������O�X�a��|>�Bf�)qX�S�"O� 0vP>Px��C��:M�$,�P"O>�##L�!�����Q�_���"O�����\�HcL|D�	1&��r��'�n�$��:h�5�7#��3d�Awo�3�ўh�TD1�4&�!�)K�9D�q�R<������?�i�&�0�@@�6z~�8E&�
���-���O~ ��@� TG�Ti��S�? "�٤,V{ �)vG$����"O~�{2i�-!�
�ħH��ta���	�h�̸
�e
R�B�1Х�0Ē���'�x\ۊ�4�����O��G���yg�L�Y��ʒ�)j7f-�ȓ_w}���'�I"�$��8�H��bO08�p�\�q_4�6+Bs�^�ȓa� �r�k�nl��I�mw~���E�y0�m�.WY�]zs��?����'D�"=E��-�':���1D�?I'���RK]�����v&�$�O�Oq�����- g�\F��t4@-�2"OLRsG��hP@Pl����q�2"O�EY���2�ƌ�MC�ei:$	3"O"�*Ղ�zLtseKN�b6�y�1"O�� ��+�l P�d�x���R�|2�2�=���:h���/\�yЪ�H�[�ԝ�	X�	ݟ��O s��|`aXCލ/5:9"Oj�y֠��%��l��"7X��I�&"O:,p�-_'=�.mxB�AH0�!�U"Ot8uj�8q�V�9��:?�]�V�'*��$K�;r!�4�֓.��1@��r�ўh1�=�'|�І�A�f&��U�lU
��?��z�>�RD�38v�x�U!�4܇�~_��e�a�Ѹ��q��هȓO����Ƈ�}S�X�(ԇE���ȓ(A|����j;ll E�ą[���G
-ڧm��u*P�U+����M?Bg����/X�"<�'�?q����� `� $M��0��,����e0!�DJ<h����cC�w��ȑLl�!�<��mJF��2G���(M�!���bni۱�A4-`�у#�@!�D�?�d�;Cf��x��� ���D��&�HO>���&��]Z�,S3�ML<�r�f�0*�%S�y�n�,R|��	
|�����'��F	�,9�bpn@ �J����;I>)���?����wG�QxD�`�\�+q�����F���`�ƋK=}�r���/E��O�`�c%�������W502˧)ZвC�g,Գ��˫x�(G|�AE�?����ODlQC$��O��!w�UiN�.O0��D_:M
\x%J�(?̕uh��t��}���<y��Z�G��B3#�1�:P����Wy�ڬ�yR�'G����OjeY���[�l�Fe���]X�-�O���&_tX��/��s���)�'Qj\Q(W�Hj5����^�mht9͓Z�f�ٵe�
yx��E`����%�\�
8˗%e��,a�gP��yNC�?���������d�4@��oe�X��M֣`tP4:C�#D��:uNϞ�f�&r,(���;ړR�?�q$
ܿ-�t�h��$
k���K��D�Iܟ�d��?�M;���?������O�����j���p���JN:�8��U�L#�q�I�P뜜��F����g�'�I�C�-CBm�"*�F���h��׮�2���.�ת���ɫRP2�Ɓ<�pس"�"$�<�>{*a�I���F{�:O�(�EGU�s?���ʅ/��i8"O��v�؟Q�j�����?��)8��'Xp"=ͧ�?y/O.�:5��'@�!������ b��rr�xn�� �	ԟ��'��'0�ɋ"⹫΍4Bi~I��)�-t!`a���;3��c����L��� 	��pb7f]>�Ak㤜:2@��D�b�š��/ ��D�b����d.ڸ#d��DI�I
������	G�'�d���D�!*D}� !^�_#����'�lb J� K`y3��R�L��,O��n����'h������~������F6#����'���71�m�vnZ���d�O����O�����&�c1�×��4�܉8���8���QƬы�r�a�&s.J �ج+�Z�sJ|
ӧ��d8 �Qȓ�,-�8Fc�s�'f�4i��?A��Dhݔa���"�^�C��%�"��(��*�O�m�c�(H��䒢 !i<H4c��'ö˓Hm����O�8ZE5	��	~��'Z���h����O蒟<�$�O��â Y*:��K6��R���	]���[���:5'�8u���6o��'��OZ��ks��"yVb���i��GH��'���۔�K�<�VYcc�V=�?�0�O[��!R%̩u�!�F�s����/�O���;?%?�秀 � ���H�c�������
�(Q"O������$e{2�B�x��08B�ɮ�ȟ�hhr�Ϥ{"�`Ɂb�c�]3� �O��$�O�aC!������ݟ���^y��'f`Őr��&#ހ�� ����u�T}i�
2L� �c�<���I�q���@�e�&��=Ӊ��>�@��O�-��^ÐtA�?#<qF��&�R�P2/�Q�^���o~�^��?I��hO��(�FU����1;"����Իb��B�I2.������u�Bt��FQb�h��Oc�����'g�I�p*�Z�
���I9ǯϔqBx則�U�M[���?9����D�O���`>�:��Ha �4��,ߵ��U�W�/�Ԃ�?�0�
ۓr��!�Խ
;ޜ(��GZ�8��%$�,��К�A��eia{����?�S�¨#�Ұ�#F�dlh�Sg�4�?����.�8��C�J�F$�*@.Z<e ,��L�1�gB�2�M�"��EQ^����iR\�@8�'}��R��"�����c~�!�d�˃�H� �Q����?���^KŪ�`�r�Z��O�C��YrQ�՜Q0�qÀ'��6��8	1G*[}$p�i�.�<P���ʉs¶��6g�?Vb�����O���O���l>��/�c���d�;n<j�S���O��$9�)� r��\�9���薁* � 
�i��	�@=����E��L�F��'��S�X��?����?iI~����D?Y��L{�υ6}\�qϖ�Tax��'|�Ov=!��Z����dL5k���P��|��O6�{��d���b�`^�0�$u���I�����\?���`�T>�I�,�E��L���ƉwZ~�IDJNK~�!}Rb���I;�ħI�.<�hT _��H���d�\=�=}�̭�G��'@�-���O�]i�u� N�>�TM���ܲ��I��	<���'���.�Ը���Z ��gU9��<��a�'=hy���M�u��e���M�M������^����_�*��FP�5�6��O�lڕV�h؄���I��<�rF]��v�o&��O��G�T�G?��l���"�A�eh�W���	���ҧ�9O~X����0���C �D�"#��}/�,��&	2X�'@콠�Ox):��Ҩ����d��n4.�
@$��^"�J?��!�@~ʟ�d�#-�����N��C#�&6�1�
�bD��Q؟��Q�W&I�$�4j�"k� ���'D�L�ED4I� MX#,V4��q���dӂ�D0��I��O��禵��m�m�5��8���*Gp���$ ��`��y��M�ë	�>@��B�˅#(Hs7c�^��W���OZN�ч%�!>">x�(Oa)�р�'�v(� ,΍=�|����N<W�,0�
�'cjU�Q{��q�K�H#�'[�eC��ţ,�<JUܡKHx 
�'���as�)l(�ZQ7R�	�'�N�8R��q�TXqI0��	�'�<��g�-��mk �͢F����'z(�����~И{RK�D���S�'�����#��&��G�;C��,��'Q�D��-_�8��3�B�5)U4�X���ON�D�O���O.́�̋C�8(�t̞-@��p�U��柜�Iɟ��	ҟ�������͟H�SB�� �(��B�O6G�<Q���M���?���?����?����?���?!@�2��+S�Q~kȨ�A
%M����'`��'D�'s��'���'�Bg0
ݎ��ʈ�s<�`1%�
6K 6��OX�d�ON��OV�d�O����Oj��Ց;�l��R�j�<BG�I3YqqlZϟ4�	؟ �I矀�������ԟ`�ɉ���MK�\�td�C��\%:���4�?���?q��?����?���?	�i�t�"�"Z�X�Bp8Äѡ���f�i�B�'`��'�"�'���'r�'�^�(�lC�Hj��#*�K&h=�W�oӂ���OJ�d�O<���Od��O��d�Ovl0P��P�d+C��`D ����玲�IП|���d��؟X����p�	ן���I�:}mp�ѳ����كa��M���?���?����?��?����?Ѧ�ζQmdM��I�	.���Z&՛��'Z��'_r�'�R�'FB�'R"��	Q�b�(�lK#|h*��2�M%Et�7��O����O����O����O$���O��^m��t� YYt�#@ $Z�=oZP~��'M�h�O�d�����r"���6A��6lcZ���'��i�Ħ9�_�fd"�$G�?��ݛDټ{�F��I�� Γ��$�)�(��7m��8��c� m�	۵0wi�t/�O���?s�1��|B�'>yR�G��IXѣQ�rZ�ā����D%�$M`�'�?a
� ,��-!8��Zq��[��p����B}��'x"6O��/5+hEb��#q|,Ԛ�G>r�T��?��(�'���������ӱ2O�j�ϭB�s�Y�"M&�H"R���'L2���I̎'��D��ԋ]xN�bK�O�,�'��	��M�"�O@`�Y��Ok3��yBM�"{Դ@d�'I2�'4r�Z�|������̧4,�Ķ�(}����r��؛�LͽC\6}���	ߟ��'�1��(KE�~��8�,0✕��U��O���?	��$�C}�Z�T_6���T/V8ꓪ?���y��i�+ٚ��i��Z͖�@���%M�&�`��'�j��Ăǔ|"Z�41�Q%:�P�FI�"l�f����R���B�O��	���`c��N�}JqPC�W,6�`�$�����?9�]�t�	��0�.X�(���E��`���#.:]9ҤAĦ���?���!N_����3�������.;R���P�G<U��
��ߞN��d�O��D�Oz���O6��,�'t~8��πT�\�����R���O�D�O�'�B�'UV7�,�ɘ_� ���W-wҒ����Dy��O����O��$αwH6M.?��h�> �e�ʠc�(��	�V�4Ic!CD �~ґ|rR�pDx¨���
P�썊��1g���'����?A��?!ϟvH�h��W�r��PD,�t� �\�ڭO��d�O�O�'V�VS�H��*�\�Q+��t-ʱbkũK��]mZ������VY��'V�'�*�B:À	KaE݉������'�J�ă49Y�<�����2��'���U���ܴ��'�2�:��-Q�t��R$d[�l��	���\;M�7������]���'��P���?��?E!��4�����w���� J�Oʓ�?)��?���?i�����PfzA�٣u,Y�E�^�^�8��?����?IO~�Q���>O����C�K VP�@���q�N|�D�'M2�|B���
��N{�v�O�	�HR�H�x�*�]c`��B�'�$=`�K?QK>�,O����O��8Q�Y$k���1����0�Hĺ���O���O��į<aZ��Iߟ��	#q��9�!��Ja&�pb�\�y�@a�?y_���ԟ�$�!���=1�f�Q��k:ڴ!�ddy�F��7��@�Q�i�0�����'���^,_��YY0�Z�N� X��'��'���S�<��ec�A�e���
����A�̟İ�OH�4��f���l J�̌���fs�B�I�����̦��۴L��H�'؛���t2W�V���ߋe_��Nݼ|�vq� �X�&�֠&�d�'���'��'|�'�D�&��{�lu��J00*� �Y�2�Oh��O��$5�i�OHM�Nu@�KT@ԥ��ʓ�OD}�'��|��4��+O,	0��8uT� P)_5A�MB��i���I�v	r(��H'���'��H��N-m�"�����2tk4�'�R�'���'U�Z��®O��d�LJ�	��kT����)�L�/�b�ভ�?q&X�H�����Γ>��<���
P�k� �$@��u��&ŦU�'� YK'�O~�O���(d��4C��X�`�0���^�x�2�'��'���'���n��Y�`L4F�4�� E�X�����Or�dWW}"^>���4ܘ')��'E��&
�L�'�.N�K>����?Q�J�05�ڴ�y2�'jR��1o߮����z��I���".Z�������4����O���Q!~��R�JU�S��<�D�t�s�'P�X�2�O����O���4Ҡ�Q�X�>q�.�Zr(}�B�ny��<����M+�|ʟ|-�E
D�Xl��iQ,��[�hT��W]D�4!�I�����Q�5���O��C��X��go�S�%�¹��'���'�B�'��O�剭�?�0�O>�xQW@P�}�S�Ժ�?����?�7�iw�OH��'�E��8�������ʚa���p�'|��C:?l�6���:��'��ɛ0[����N�T��X�vH����P���	�`��Ɵ��	��X�O�P��N���x!��M
o���Z������H�	_�s� 
�4�y+�J����Y]n`3&AX�/��i�&�O�OD�]���i��$�.��U�Ů�7j���
�.M�)"hܓ]�`�	�@��'��������4(PV\R�Y*��psf���D:�,�Iџ���󟤔'g���?y���?y"ĒȽR�K,e"<9B�����'~��
���wӐ�$�Ѐ�M-"zʬZ0eH�l��ǃ���ɻɆ(
��o||і'��tI�՟���;Oح�֋�4s�,�[�ƭLbz$��'��'q�S�<)P�I<��8��#)��9�G$I��l��O˓Y�6�����ͻ�o
:��8�����S�R�
0��O��oZ��M{�ixj�`G�i_��=�݀e�OR�e{wa�^��M�e��@����@�IKy2�'R��'�'1���f�t4cd�?w�nա��(��	)��d�O����O
����D3J�r���E�j^�19�	�|9�'o��'Lɧ��'"��$N�M��%�KT�kuFW>�:�F�i���]'�8���O��O�˓,,ɱ�E˨� �.Gd]h���?����?���?q(O��'=�� P`Y�� )�&����&�^�rD�'�:7�6�I����O���g��C׌ % d�X �<$��{��64?��Y8�֣|��w���C�qzl�&��o+�h��?����?Q��?�����.��$i�i���׎��>�f|cQ�'��'ʘ��?���Fr����x�����`�q��!�5I�	'q�'�2�'y�ℕu+�6���~�8ŉ��˄q�ɰa��2�~b�|V��Sٟ<��֟\AU�4g �����,�������ߟ��	my�L�>y/O��D=������X*Л��K�uy�>��?9I>��ܽ�@�@2JY�x���(�ؕ��]0	�px"5�iO�ʓ�ڕ��� %��
��.2x8)�t̓ r�3"�ݟ��	ܟ����8%?��'l"���;D�t�A�Y5 ��1j4RQ� ��4��' ��?�$��2�`:��Q9
` t����?���s�@ܴ����B毱?)�O%R��P�O$i
�e@#7�l����d�O��d�OP�$�O~��&� ,'A
.]b"�]=~.�l!�kC��d�O��D�Oܒ�����͓5Dѫ��)�q�F��
(+p�	ݟ�&�p%?xP�즥��b�@���$x�\����)ۜز ���&�t�'��'c
�r���,���ЖᑊO�����'4�'R�Z�X8�O����OX�DF^��uKi�P��틅�\j㟤©O,�d�O��'��k� B�w*`R�jZ�6� ���Cfy�I�i3T4#����4�L�P�2�	7_
�2L^5\Ҁa#V�u<��O����OP�D7ڧ�y2IX����@��.
ًÏ �?�0Y�x��ܟĈܴ��'g�4W]�� ���Z$)����#62�q�Z�nZ�Mې�G��MӘ'rR9gj|��Ѻ;ŋӐ/�*�X���E��r��FH��Sy�'Yb�'U��':�瘚x�H�)��Sd<1`e���)Or%�'U��'�����'��@��l�&$h$z&#�N��� �>�e�i�&6�HC�)��;�n���[�DC�q�QYC�`��c�f�O��hJ>i*O�(ۂ��(O蹚5��7.�`����O�d�O����O����<i�^�x�ɯ|��ݓ�Ri>$�q�C�GU��*�M���O�>I'�i)7����HX��.c��{�N�&,����F�7m!?1���24��9��ݼk�OO�����0閷;����5��0���P�I� �I���F��n��0�9R��F�`噗P��?9��?y�]���Iٟ���4ט'�h��ᬖd(�
�DηC�e���x�'Gr�O�xl:�i�	�l�n�xtxxj kƫ���0��J�F0��g��_y�O�B�'6R�αuQ�X�#ZS��MAP��h���'v����d�O����O\�'}\h�A'�P����'I���'0D��?��4<�ɧ��ɼ3�~�2�Cɉ$Hƫ�6��:��-����O:�����?9�$����rb\M{4$�	���'Z�Z���O���O4��,���<1b�'�v���V�4ji�6���J*B���?A�B��&�D�`}�}�*�A��j�،.��Q�GÐ5,G�nZ;�M����M��O�xr����O|������:$x���N���@`_����'���'���'r�'d�
����(*{-��2��ʹ^U�1�'x��'_���' �7�{��@  #���jJ\�@�g�O��D+�/�	CR;�6͸�\�AK�CQ�!a�͙�\Љ���O� �X�~�|R\��|ᄣʧ ��,;ա�:(68r*�ʟ(�I����	My�.�>����?1��d����ɍ�A�x�*�.[|8Mяbį>���i��7�{�	=fhF�B��������h�>T�P�'�:ܐo�I�PYp���KƟLpW9O�X�̋�<�>�{�+�:ia&Q��'��'���'f�>��taB��&�,v<d@��hm,��	%���<ѡ�i��O�����a�I�!��(\ <c�˅9"d�d�O��d�OD��S``�v���jpN�~R ���a�R�:qL+�� F��'�l�'���'���'1��'��[t�E1Q��QAqO�+10���[�x��O��O<��7�9O�i���9^�N�]/v�aEV}r�'hr�|�O���'.��S�M\ lN�+RNY���=�r/A������,;�J�4��D!���<Y�k�
��X�'UcCF��g�O��?Y��?)���?������\}�'6�)��A�q�����MI�O����u�'N6�3�	��$�O���k�@i�E�=` ��" �ٚft85o�/@60?�q ؼ:Q�|��w-ι�P�K]����=Jq���?���?A���?�����@s�;����H��(̈ڂ�'���'�T����զ��<��6l�N��#���f�:��E�Pd�ß����8s�eM����'��YÑ�M�:|v�@tʽ^f-4胰��������4���d�OX���=��-��-ڝ$s�Ƃ��TE����O��S������	��O���9�f�x��D.ɔb�p�*O4��'�2�'�ɧ��]gT��ׯ��b��DF�4)�tFOF�07�!?���;�	l�I�$q��a�ndK�)�-<����	՟��	��L��L�Sqy!�O� �-�(d)F��7���T�����'��'�N6M0�	�����O�`�D0�c�s_�p	5�O�����Bml7�??���I�c�c?���l9����N�-���B@��O8��?���?A��?����';����d�=.�\ˇ��2*o<들?����?aJ~�_Λ�4OfU3&8Z8�<����2A�N�� �'�2�|����D����O�M���J�el�I�#Α�o��X��'��[��u?	L>y*O��O�-��]�*��a�.[��j���O����O����<�Q�4��ޟ��I��ژs�HQ+�����g�?�bP��Iݟ�&��3b��f\�P�I\}�"��ǈZ]y"B�>q�<-�f�it�i>)���O��I�W�D�B+F !�.��0���J����OH��Op�$<�'�y�ڃ
�6�0DNK<~<>L���?�Q]���'�Z6�&���?݀a\7r �ڀHǧ��qchKџt�	ϟP��sɊ�m�P~r�	�����"LQm�'{�������V�n �Ɣ|�X�4�	��������	ǟx*�D=d�*,Y)��G2h��Sy�f�>����?������<5!�>2"hp�h��F�<(Q C�>!���4��C�)�S�q4��f� 
��qQ��� 4|��$ٖfv�:���`o�O��L>�(O	�j
�X*�8���	N����O����O���O���<QBQ�<���B� ]R�K't�4Ui��о3f>e�	"�Mی�M�>����?ў'��z�C�7l�X�*�+z"���<�M��O�m�G*����4���1�^�[���{g����ʂy��Ղ��'���'���'�'v>�f`�>SS���ߠ3#��/�O����O���'���Mӎy�E�T��t�.W)w�Z]�2������?���?�ĕ+�M+�O뎜�Sj��Asb�&J��{���=o����f��t&�T�'���'�B�'<iv�O� G\��/�V�\��'V"Q��O��d�O���<�Ǎ	WE��7�#O��Ӈ��cy2��>���?yI>���!Z�&�'���A��8 ��A�ǜ�e��lJb�i���?�2��OГO^aʳ��>��	�b^�xN������O^�$�O�d�O����S�rQ���l�^��0��-�?�)OƝn�Q��Z��	Ɵ\�6l�0���@%�z6�P���ݟl��e >9n~~�%L*M$H�~��D�M&�����&[��h`�a�P�'�R�'	r�'���'d��>\��s�̚H�`L0�������'fr�'����'¸6Ml�Li �B)T6�l��FI|��ҵ��Oj��(��+�� @�6m���Y0�T�]���I���&vr�-��ON�����~b�|�V��Ɵ�Zǁ��Ԉs���mq�G����T����D��eyr�>���?��)��,"��:B���jA�T�@�z�#�r�>!��iDN7��u�	�1m��!��:3E���5�C62���'��x�-+��4c�O�阞�?9��o��R���	5��!�K�S%�Z�2�'���'*"���<� �4OX h+�$�C��L���Z���s�O��D�ON�lZ|������ןm��+%g"(Qv1�Q��?����?� �i!>�ói���O�@	Dʳ��]w�@L3#�T�e�"�\�E�m�O>�*O��D�OF���O<�$�O��*�����Xy0R�ۡ&.� �<q�R��������k���l�vg�m1�� ��K�ZMX�8��dCɦ�ܴʉ��O���S���h+�݋�n�{�<���.��$��O�U��_��?1G%�d�<Y!�C�P��nH�\nv����"�?���?���?�����W}��'���e�����P� ��-�#E�?��i��O���'�2�'��dQ�z J	�#���CLA5z"��ó�i���1��J$�O�q�(��%HFT4ɜt�(�z2 ����D�O��$�O>���O8��/§>�B �ŝ!z�V�rFb�A,ty�	�4�I!����O����1�<QR�]�h��lyw�^zJ
CM�����ll�T���'E>6??y��U;=����ƃJ�Hk�!I�"��	�C�Ot<�L>,O���O��d�O�dؤ�������dA�K�2���.�O����<�X�X��ٟ��	g�ĀD>X/�L���$G;����#�
��$�T}��'<��|�Od��>&�n�jd���D�Y�Mf�Tcb-��������6T��$4�$�!)��㔎��F�_(A|���Oj�d�O���*�	�<�s�'aP��E��T\ah�W
l��ݠ���?q�hr����\}B�'?D�⠅�0U2� ݳ,0��sg�'�)�->H��?O��d
~4�L?牔�� �0KR*F#�5P�k]0@����By��'��'Q��'W2�?�Ц�J�.�̚�^x�x=Rto@E}2�'�r�''��5nZ�<��EEl� ���82PlX������	P�ڟ0�	���H��̓ J`�)�L�-�c��8(�-��A�ẟd$�������'p
=A��E�c�2h����QUJ�B@�'2�'�rP�@�O��d�O~���ip�MI2ύ�p�x�Bsj԰%�P���OFHm���M���x2��-��L��M�����K#@B��'�d�3���D���O&�iЩ�?abh�܁�C��6<��/�}���e��O���O���O6�}Ҟ�� :t��Z+U���QWNКό���'b����d�Ǧ��?���1�,�c��у#kb,�v��dU��b�?�vLmӠUoZ�3lnU~B��9֬`��$zL4��DJ/.h��ֳxU�����|"\���	ߟ��	��H�I�$� �E�-�lsB�2e�
��sy�ϯ>)OB��;��>K|�-�'TMFxc"�F:]�x᢬O�<l���M[��x������J�l�����U��	��B��@t�	�&�X �'��%��'~N�i�q��$�����b�'�"�'���'��Z�b�O���yl\}daI��!�c
9�p��^Ǧ%�?�Q��K�4囦C�Oƍ�#cÓ0L������Nz���^:y���(���Zp$��$�Q�ʼ�HX��蕥Ylڅµ�ȟP�	ޟh�I����	Ɵ�E���ΰR%�(y f��3a��$"]!�?1��?!U��	�d۴��'|����aۮGgZhA�`�&��	�O>A��?��W3v��4����x��b�Y����k_#Y��5�G�{��I\��|y�'���'�r�o3̩���s��9bG�w��'������O��$�O��)�.L��덺.�:���X��'����?����S�)F4��b ���7XҼ*1fΤ`�b�A#��ݛ��<�'O�d�IV�I����Ѣ���,��������Ο4�	�(�	\�Sxy"��Ox��wG8	���Q�~1�)��'u�I(�M��r�>�ջi5� ��!���3ͅ�1,Naؐ�j�6�oZn�Ftn�p~�a+��Ӫ1&��=�ݙE�xILmh��7H���<9��?9���?Y���?)˟ƹ�FW�G�t���G`+�m�To�>���?9�����<郾i��D�=\�!j�a�!|����5`T�p��6���a�N<��'�R��1v\}bڴ�y¥Yz�:��W-Y�X�28�e,�X�����ʔ9�i�O���?!�f��ŻP�(3�`��H�[^�x9���?���?/O��'}��y'%�C:%�m%5{,M2�<��O�)�'���is(�O�	���?���XQJ���RtJ'�'�2˘�jJ���,ť���������NI牓bK��[�:��<���������Oj���O ��-ڧ�yR�4 �c��**<�s�H
�?�AP�T�'��6�'���?��ׂΩvb-0�X�`��E柜�	�H���	�� o�<Y�� *����~�T-ذ6~p��.&X!mf�Py��'�R�'[�'�R�Ğ ��PK��9ia��+�Y6*~��:��D�<�����'�?y�dN�o������5����o-"H�	�MS�i��O1�����%aY� ҩ�<<��$K�N�(z�HP.H�	�d�I
5�'���%�L�'z��2BEr|�!JD�M �N����'��'b�'f�S���O��$� n&}`�aI�/Vz�(�fQ>j�X��YǦ	�?��Q��ٴ%��F�O�a7$W�#~B��Q����q ��[.U�v���)vTiD�4�)b��v��g2؉q��3f�ȌCP��O��d�O��d�O��d�O�#|b�l�X���r� \Kf�5%������ퟤ��O��d�OԱn�J̓EJ����@:G%�)� Y�"���IL>�ݴ8F���Ox���лiB�$�O�,��gGZ��1sӃB1	N�B��D����2=*�O��|����?��s� @[ #ԏ.Lhp�l 5�T��?)*O���'Z�����OL���H�V�DT��!_?~��-O���'��'�ɧ�ӀBB�D�UM�(��M�F��1�F�&d��x�.��R�����?��Fy�Ʌy���b��c�]	WHO-�	���'���'�"�'��O��ɷ�?9�E��4���2��@��ğ0�'�X6�"��0���Ot�v�Bc�"�ʅ�,Fv�j�B�O(��!u�7�:?�;T�<���O���5�j���Oq�T��DG�� GZ��<Y���?���?���?aɟ���@�Y�PH�gi�g�ꥒU��>����?�����<u�i���׈Xu 𚔧C;M�I
��Ӕ-�R�'z�'��Os�a���i����(U6��
�$�hNµ�be��Q����������O�d��H�pC��,A��r�U�#����Ov���O�j
�	�������A��b1T�7N�	~j���f��4�����IL�"X|�'�Er)��3Ԃ9�$)�'2�����sS�&C0����~�8O�XJSꜳ nP�rC�ܓ/?�MC�'���'���'��>E�qO\�7ƒ��T�w�Y�$��I�I	����O�������?��� �ٳ������i��kR��ޟl�Iߟt���+6Έl�v~Zw��crߟ&�����L�*e#�)�*l���8���<1���?i��?I��?9Q��iP<�J�" ��n%���'�b��?���?QN~���=I���M	�!�у�FI6=���T���	���%�b>�X��ъ�|�EĈ�,X�b�Eqndm���`�(��'��'W��7|�`Hp�ޚ����&E
Y�"h��՟��I՟��Iҟ�'w�듦?rL��=�����C�'�ze�� ��?!�i1�O���'��'.�D�mL&�)d�/T� �
���[� 8�t�i%�	
N�n9��ݟ<�����Z����l A� N)�.���O@�D�O����O��+�g�? h�%ݸzc�@��S*ʸL���'Q��'r\���ߦ��<)��Ŏ
�ڙ� �6N�@m�SM�j�ޟ8������'�ΦΓ�?U��R�[���� ���@�!���0�饟 $�������'�'_B4��k�*nYK�e�1vD�qiu�'��W��ɮO���?aʟ �&�
k�N��tK�'v���� Z��+�O���O֒O� ���E,�A�h�����Ja��/W���ne~"�O�^����N�j1z!ė�m@�X��P�$t����?���?-�M�M~b*O*-�I�(b`��E��R�|�GH�g�H�$�<	�iK�On�'��$�=P�-�4b�]S$C�,��'��X���i*�ɫGi�A�	D�r�p8����.^c�)r�aE�H��Z���	ɟ����p�Iן<�Oh��3� �~,�I0��P'��9�U���'2�	�禕ϓkD���D�_,i��<�D���86��	���&��'?A�I֦��Cl|s�Z.+�9z��2<���	0G�e���O��O4��|��C�|�	�f
�9�� �)���Hy��?���?�*O�|�']��'cbgJ
G25٤e�
_����C4`�O�t�'�07M��uYH<9RaR��Lh����vd6��������3����L Ȇ�������"Ȑ�I�y�ax�D_p5�ၣ��V���O���O��D.ڧ�y���m!�	��)�PL�yp+���?�Q���'G�6-?�I�?�w�$��K2��3lՋ�A�ԟ@�ٴPH��gc�0sGf�x�?R�Z'��DqҶ��kv�(B�G�0تl��
_������O����O��d�O.�dҕd��hh��~���CTe�I�(ʓ2N�I��\�Iߟ %?�ɉ�h���BΞj_R|a�f̬KR��[�O�Qoڷ�M�U�x�Ot���O��u�(Ӂ)U��y5��Y HƇ�2	�4R��xRnA�r J�	gy��P�\�l��ӃW@�`c+��F�r�'���'���'�������OVm��b�*#hH��8Q��L �G�OȤn�L���	���I�<-U�N(S��>Y�q@K��%k�����h�
����T�i��}y2�Ow󮞨&\ ��nC3���3R&�[Yb�'�2�'M��'.�ᓫ\��A�Pi�^��\�S'/I"���?r^������4�ٴ��'�>�� E�]6�:������M>9��?��K�,q�޴�����ؐ�9NvZ\����'&��0C��

 ��I^�IDy��'s��'.�ͻV��&j��}/@y�$Ş?]�'��	����O����O��''��$8!�C�4u֍�Ы�s�(�'����?Q���S��� IK���c�u`uأ��^����./�����<��'m�t�	E�ɷ.6��:��B�D���X �Gנ5������	ԟ���|�SFyZ���1[0�;�,cQ��K"�'��a�b�dp�O~�D
�>�����-
�*T�F"����D�O:��hn��Ӻ���K���?���ފ'��X�CE�xL�m2���O�˓�?a���?y���?!����ְ16�d��i�?�b ��X���?����?�O~���S���?O�愋�� t@rN��=� ���'��/ �d?�I�t]v7M��:��"-��򂨞*k<�tI N�O����BX��?��-���<ͧ�?Q"���8VX۶��7f�"j���?����?�����DB}2�'Vr�'�m�f��*K��M@夝�h9��YP��MW}b�'_b�=���nМ����MRg([
���wo�`& A�Xu6�����ßP(1<O�E�Ӧ¼F�h��Փ�����'xB�'���'��>�Γxg:L����'A�`�X Ě��8������O��������?����A�&#�� ���1k��&
�9���?	�����3,Y���А�GU�����D1���=sԊ�Ud�n8�D��|bT�x�I�d��ܟ���ʟP+��п(���aOE�V�|P�doWAy2��>����?������<IU�����OV��F��`��27��$�M�ihO1�8�kw��?"�aǊ1{P<x��I�_�҈��i�<�X$4M���'>A&�P�'�f�h���Q�a
�/.kd<ѐ�'��'���'EB\��k�O���x���^7@D�m�%��5�������?�bX����۟0�{�b����L�q���w�����J���'/���f�c�O�� >4ڍp$UJ�鑃S�AR�'\"�'$��'(R�F��t\�M�^�$���w/��$�O���PL}�V��ZٴƘ'Q��"��HJjQ)���6�N>i���?��?%ְ�۴�y��'ˢ�"uH*_��4[�+�iy�I�^L�8��䓤�4�*���O��dA6i��T�f���WkH�!Q�������O�ʓ.��	ܟH�I���OW�ͨEă3\X��T�/>�T��.Obx�'��'�ɧ��m�ཙ@'_�)�f�����w%�Ы�/��{:(7��Ny"�O������O���˴eD:t/:rW��)�e���?����?�������� ��,l%�͒���)�4���O`˓]����W}B�'�"#�q��`	�D�"�>0��'�-�"p/�V>OD���q��h�'��$�N�P�6e��n��'��D�P��<���?I��?���?Iȟ� FiH1�X�ck�a5�޲Dr�(�c�>y��?�����'�?q��i��%1��p�H
3Bp @##�B��'��'8r�'��a "8]�F2Ob��E9?�P�S�ġU�`E���OX��@��.�~��|rZ����͟���x3��W$� ��Kp�DƟD�	蟘�	ny2#�>!+O*�:�4Y�$���~�x�^�[�&⟘z�O�]m��M��x��B�a�@�� _)���S��I�|���r�H��C1�'?�j��'4�ϓ.p9Ҁ*�3NXtj��ݙ"��������	����m�O��@�v\x}�"�܀�\s�J�?�b��>,Ol�_����s�uL����K
kT0ȣ��;�?Q���?��aŬ�{�4��D�=�l��'�b� �.2��,���\�E���2�)�ļ<y���?����?���?�W�W�M��=�(D�@���)�"��n}��'��'��O��LB�5�N���)]�|p��I�EG6b� ��?����S�'B��}ȁ�8�&,�Pf�7��|��6�M3�O���]��~�|�^��YsO��o("a�O��ɄM{���X�	�(������	py���>��bp���kW	2h���r���j��X����D�o}�'[20ODI��MUv�e�ܯ7�X�K���Uy�����c-]RQ>��;r�����/��`$N ��(y�I��P�	۟��Iԟ���R�O����Aa�!Z=�mC|�
����p����ĭ<1�im1OzM $�ɇi�d,�@Ñ�!��|���|B�'���'e~źƸi��I�^C �֭�,6)���%A�_��P�Ͷa�2��n��wy�O��'�¯l������s�E=Ӕ�����?�)Oȑ�'�R�'�?Ys6�?T�[0@�0d*�Φ<��^�0����d$��OnH�T�����ION�:憎���&�[P~R�O3����� ��'7���&M�r6�9ʗ
M��5���'���'���'��O��	%�?)���5D�uR`�ײr�2��U�󟨕'��7�.�ɱ����O�
7��2��X�$��� A��OR��#X�7)?Y��*i ���&�� ��,9k�j�?�X$8�,֥�b_�������I�4������Ow��r��E�pH`h(����p�R�CwT���	���p�s���4�yRa�h� �a� 	m��:W��2�?������}����4�~���2KY�kY0`�zE��?9�D�~����+����4�����'n6�Iq/�O~�8jP�P�Eb�D�O��d�O:�tX�I̟|�Iϟ C�Ɨvv���&׊9�`�����a��0����M���i)�O�@��#ϻv�bV�]�2�@\���<���J���4�r->��'������y�E�s� <���;VTh3�ȃ�?���?����?	���o�pr1(�' �N���兎q�:�kGG�OB��'-�	�M�b�O#��u���
`�wO�����&�''J6-H̦���4*$�[ܴ�yR�'�A��o��?����U8��]F��G�0X��┲r�'��	�������͟��,2!��o�6J"s����R�T�'���?	��?II~�ՄQ@GJE�5��A�Kӧr1�!�w]�,��4d��vn&��IO$�&o˽{��S�Hv��ypKkR�� q�+�!�O�I�J>/O�D�գ�[��j�BC�c��S�o�O���O���O��d�<�^���I�b3	HLP�U�i���1Q��m�I��M�� �>����?��'� $W2J�
G�SU�\P	��)�MK�OR�BB�a�E��2�:�C�L�>tb�Bs��n�=#��'2�'�b�'D��'9>�)�A|3N�;Ê�D�.M2��O`�d�O^M�'�I��Ms�yB��>���s�x�f�����>v�'�7�NϦY����J l�<��tJS��4,��̓�JY0�8��k�u���ͼ�����O���O��DI�2j
�A�S�Kl�,y��="l�D�O˓Z��IΟ8��ӟt�O�l�wi]U|]��mJ-<
��P-O���'8��'�ɧ�S?=��$7H[`�B�æ��f����B�YR�N7M*?A�'aN�	h�	07�8�b���k8��Bd	 �B��	�����	n�Sby���O ua�֌B��P���#KꠌcE�'�B�'D6<�������O�Ճ�Kу]I�A�� �8Lj�Ɔ�O���%[(�6�=?��R�#B�c?q�5��{�.|T� e��� �c�O���?��?Y��?�����I� ����V�ղ<ښ��`I?����?���?�L~�,I�9O�����C�,0���_5p���S�'���|R�����nܛ6�OzD�f��&�����+ИX�
!a��'$�j�]������|�Z��SПx@[�
T"-s2�-7l��¡���@�I�����ey"��>i���?y�.�#�l��������s�]h��>!���?�O>!����\�z�QD^����u��$�O� �D�ޡ?�@1;����S9Cz�
��<!��E�(4�0Ջ�r˶��4)��\�I̟(��͟�G�d=Ot�����zL؛�ꀛm+�	v�'>������?Y���
�Òn��f  � �jѱ^_(D��?i��?���M��O��v,���z\w��M��԰R��F���R�O>�.O��d�Or���On��O
� &1���\��Up lָ����]�8�O���O��d=�9OZ@xTA2r�Y�!�.���P�D}2�'���|���;P��`wON�Frx YE��=��!�iL�ɅV�|�O�O0˓{�E�ł��>��I�FW�f�x��?����?A���?�,O�Q�'N�7{���d�(9 �t��
$WC�o�`�tҫO��d�O�扬� ��G�
���ti�d|jeq�hp���4;\�10k'�'�yW�ϊT�\eQ1l�? \��u�vc��'5�'���'���Ӏ!3 �Ss"�52��
��&SB�d�OP�N`}R�ܡ�4��'ќݰu��y|!��,w�|�bM>���?9��^j�z�4���T4T7*��	��w,$p )̞z��J��O��~2�|�W��Sן���џ�ӆEoh�A���ړϾ����ݟp�I]y�E�>���?1����3$�"�Z��X		:Ti��܆I�I����O�d?��~��1�Ԉ�c낞 q�R�(L�!.��s'�٦ݒ+O�I��~��|���uR�y*��rF�p�O����'Y��'"��P�@��rH�P �H!'^�ӒgY�!�T��IEy"k�:㟐ӪO����=h�L��E�>�t�dbQo�f���O�M±�w��+S�e��F/�S�NVH���Įs�R|�`��b
����<A���?���?i��?�Ο�����'�̉(��Ŋf��HRcJ�>���?������<)V�i���^�|Qp؉�#nVn��(¾[��'2�'q��'t��
*�v1O��H�E. ��I�@f��DȨ[A$�O�2�؄�~R�|"\����X�OJ:G��8S�J�>Bx��A'G ����I�����[yȷ>����?y��S�x���>r�4���7M̕��̣>���?�L>�7c߄B���j�*�V��q�.����Ѫ#`X���.y����|2eN���ϓ0��!č.[ꨅbUO�0C�ru�I۟d��퟈��j�O��D��^f���A�pcd���K'��>9��?i�iD�Ov���u�� ��(5�ԉ�����2�(�$�O��$�OrL��sӆ�Ӻ� Ҽ��� �-�<9��인*�B� oJ �'��I��0����x����l�	�@��Xa�E�: \�Ȣ�[9Q(�8�'�`��?a��?��`I�]X�����=m�hq���8I���?�����O:  &-�B�2�Wa�&bLt�7��^^E �O8�oĵ�?�@">��<���5WD>�A��T&$�6ݚuf���?����?���?�����$Nj}"�'��8AܤH��	���i�p����'��7�?�	>���O��dq��y��a��Y3��L9�y��C~+<7�&?	�A��>dT�)9�Sۼ�EˮX��RtfD�TSD�r ��ӟ����T�I�8�	��G�4OW8<�؄!�-l\ɚB���?����?��U���'�46-/�I�O%&|hG#�E�qwٱ �
�O���O��:7W*76?�Y�,�3����Ex`�i�،��Aa�O<�SL>-O��O.��O��5o�J<L`�!H�l�$�@N�Ov��<)�[���	ϟ(�IA�t�˿q!���a@=l�`G/ ��A} ~���nں��S�i޾�J���"ǀN@a��Lo�<�ӡ�	ktB�HГ�l�S��2�GP�	�94�T-��A����:Q��}�	˟����(�	L�S`y"a�Ov�F�!.jC� :6ǲ��''��'P78�����O���$I�z�S��U�@kӐo�a>�m`~�d�?I�|��ST��+~�j�nD9Gǘ}��%��;��d�<i��?���?)��?yȟ���NQ�Xx໶��2�F]�P��>����?����'�?q�i���
�e�8V��u'6^O�ֵi��6�z��_�Su�N�lZy?ђ�21�� 1�)ߠ>C�Y0$�4SC�B���e�IVy�O���Ҹ#k��u�ۅ^I|A���:|�'�"�'~���$�<���+�0X3dI_�B���[��e�X���)�>1s�ie7mPs�i�u9�ix��yӎL#.��Q2T��aC�|yZX��F=?�'7�����:�y"E�{-ҷ��|EY��?���?���?Y�������w�\��ʣK ����b�'����?Y��5y�V��矊�pc�
�� q�<rԝ���j�������ߴ&mL)0�4��� �Tr���'�uw�_�Uܦ�+c��sw4�JH�&������O ���O���O��D��(����f�d�ڦ��2�f�E<�	�����㟈&?����C�X��!Y�e�-����I��*�O�%oڪ�M��x��$��.F)��P�C�[�<)��
B��r+����$�	������OʓjxJ�B6gߕ_X&@J�a	]0�t@���?����?���?A,O���'��Ȑ��(�[��h�&l-��X��'�,6�/�I#��$�Ħ)����'
����$I�C*����Ʃ?�v����Y��M��O��M���47���ЀW��´i����S�B==��'r�'T��'=b��-7�zX�o��T�nٰ&7U�J�$�O��A}b�'8Rf�*c��y��<ZP�@�a�bCr4�V"�d�O��c�0�w�v�x�4��G�6��T�aF=j���i ͐�p�~��h��xy�O���'��� @�Ҷ��Ms8̂���~�Ӧ�'�"R�(z�O���?a͟�MJ�ٱz�X
���?�n��[��r�OF�$�O��O�')8�e�Ϝ�W�V�{�O�"^Qb��b�X�-n�B~��O{n����?�l�PV�Ӥ��#6'\&�l����?���?������DW��:�Չ-k]��߳6��1�F�OP���OD5o�~�z��	ğ�����Q��U��k�$=�&��Qʈݟ��	���l�l~Zw��i��۟��'`@V%�1G�*}6�-pN���젉&Wg,�2�ߧ�|�h M�rf��E� i����M��Ɯ ɧR!�ꡠD'�6������~��p��ͥbD��� 4}�ى��ȶ��X%e�t���Hvb�Q�s� �#��lR���sĉ�[[*1��)�*"���!�%�{6�)f�$��|�3K�Xn
lѦ!��hvѠb+� 6��y3�,fؓl��=ư�W�=�� �U�7��ɻ���%j�;��6�o��!��B��)�Vx	�柪 S.ꒈM-d����Ͽ:t���rd@�$��d"w�]*�K䚠4k^�*�J#x;�%A2
M;¬�Vc8؅��(�v����Z<1��׈r�`t���Y�����a�+ݲ|�G�E�$z�x��J)[�̘f�0�*c�E���Qc�?���	ŎN6\xB�&�6z`�h`��d�Q T&~}*M b��5�a��Qt(��%�*B(�b��4i��A��ڲ��ԮE2@A����o��=rBx�0���O����Ox�'3���|�<���%	�~�h�q��'s�~��?��h\��?9��?c��A~����i~������?��?��W��'���|2��ۜ�)!�Ú$f��᭐-#��	!^ބ$���	ן���w����>���Qd@��Y�2��L٭�?�Y�ؖ'�b�|��'��H������,�T���lK�C��e�!�'������I͟x'?}�'Co�J"-ʷ���3f%�e��L�	�l�Iޟ�%�h�	ޟ�����[�DA6P\�x����Dv�i��`y��'"��'��O���?��i��W�u"��I�+��Y���<q�����?y�KS�5��y�b�=(0��wNR/(�HL��GR(�?	��?�*O��d�J�T�']B�'[fds�B�U�J� "�T�Tt:آ�]���П����Z6�����{>ٰĮi��\��]����g��O(��?����?����?����򤒧f�"%�f�`�V}�Emġ	�4��O��(2�D��>yكc��^74�R�׀dC0�p%��O��D��i�	ǟ��� �O2�%�ء1X�>g���$r�Ah����Fxr���O���ڵR[d�23gZ*}�ʄ"m�����͟H�I���	�Of��?��'�"rAG	nPhP6皞�F�Q��"E���'���'���,�2���l
T��]/p�p9�'���'7����D�O(�O�q�aGC�^�̫4��1��� �<ɇ���?�+OT���O���/� ��"[^9�⠆+E>�1W��؟)�OV˓�?K>���?yg���$6�H�*<�5`2 ��f����H>���?����������Aq��Elkz��@O_��?))O���&���O���X�ʰ��#H��e�e��I���� �>�ʓ�?q��?�J~u���l:��k3��?}�\`�N�>8B�'��'9�i>��Ip�D�!W 1�u�n���hC�8�?����?�.OD�DU��۟��;����Fƞ<]�$��!|�Ν&� �'�"�'V��y���`qJ!�V����b
�C��^����%�M[/�����O�L�'a����d��A�N�% �e$,x������O��>�	4��J��ҥ�ĝ�x��G[�=�˓�?���?����?!*O�:&�}1hZ=�ܔ�!@�A�V��'
`����Ӻk�8�i�N�x͓U�.�4��՟��	����	CyʟZ�3�ȵ�j͞F��1õ�ύaPf�f#��Oy�6O����ӬF%���A�,M��Y��':b�'��	P�t��0O��q�
bAA\�\����P &���"#]1O����<��'��b�
�[}�)�����Ƶ�������O@��?�Iȟ��P�>��@W�c���SԫA�4p���q��?Q���?�L~�0�Or2t����<1��=���S(g�\1/O���O��O���|B��l8 �w�:�P
���2J�p8O>����D�</���$ޝ���YbA��O[����ѹ(K���%��񟴔'%:��K��r��'S�&�7�[ Y��a���OH�d�<	/O�˧�?����yW$Ϊ,�x��akۻ9D��M ����?�/OL���I�D^�8�mI�^A������!Q��cy��'X6��|Z���?Y�R���랸\Q��2���ۼ52&�O���?����'��{̾��!�	$�l�e�>a�D�s���?Ǽi�2�'OR�'
�O��
1�6���ɯ!��8`4KC�0��'b�'�ɧ����j�(2�& �냸C�0��Ӏ����	Ɵ�����ԗ���4?�6����Ff��oK�5�aoN1<N"<�I~����?���I�<a�F�?e�`M:�J1?�@*���?Q�������!��Q<cb$dx���1@�L�L	]SH�O��$�<���?�����W�~t�D�d�E�{Q��C)?q(�d�Ob��3�D�<�� bhw�ݝM����%��q�R\��'�]�|��ޟ��It�S*��S��*
�HRa��o��'Ly�'�R�|Y��ǟ! 	��Zؒ�k߮<�����O�Ky��'�r�'/�OS��'�?m%O�d��6�F1	���?������OV���Ovh����擿b�,�i��;D�q@)B�(^�4��ȟ��I]yB�'�\맾?���?)��Oa�P��� @2�t�
���O���O � �;O��d�<�;\&��e��-�p%�1�Ԝc�V��I\y2�'̈7��O����O&���q}g��S�ТAo^<:���Ȓ@�8M`��'����6��ģ<Q���nL�J
���%F�������D�?��WX�f�'�r�'tbe�>�/O*��p�B�2J`�1f���u!��@g)�O���45O��<����'Z����B�v�V8R`��{�d�Hׇ~�����O��O
��'��I�X�Ft:���� [r���*�6)���	ɟ�'���Ce��$�'�B�'#t3ǣV�r!W��`�]��'=��'�>ꓻ�$�O���y��B��V�ʥX�`K�e� ���'k�I�'����Ib�'g���Ŋ�$]*(kf��C�L������D�<Q����d�O��d�O@��P��-�VM�f����>����� ��$�<)���?y��� �db\��Z�6IR�DS�Y����?(O���<	��?I��tU� E�ŉq�]������,��!�	ܟ���IBy�OA��g���%D��`2�U)Y��L�k@�����Oy"�'�b�'J�9�Ο�牰4��
�HQ�g)fT;1�mD���Or�D�<��7���ΟD����X*"�W�@���P2ɇg����#Cy�'#r�'���'#�'�C36�3V�T�Ya'�Y�B�rS������M����?���?1�\����@��h0haAj_�G:�d�������֟d�b���IQy��	LS�aR$CE�h��M*.�+�R�'�R6m�O����O��ĆJ}^��h�ΜBv��� ��NI��l���q�.���O�RF�_o�j�E�&l�$MKC_�7m�O��$�O���x}�U���	�<9��x�$�bg.Q4��'G$�'�bˁ
	�O��'0 δJ/x��C���Pi� �8���'d�,���O
�0���vR\V!x ��mU�#˓a���<a���?y���ɔ$Ir�<3�`��!�ԯN����E�'���'��'���'h�"U�)v(�!�x86��w"ɂW$�R���	ğP��J��3���DA���XqQ�G��x�	XFyB�'R�|R�'Lր�~҉K'%�f`���1-(�ʐ逫����O�d�OX��d�$>-�bO��snQ���zV�P����,��U���(�	�-n�e�IL~�+��=��HɣC�#(�
�������?9���?�*O��dRa����H��d���&�р6^�5IB���L$�0�I�� ��E�$�H���̈ .U��BO�<�2aP���O�ʓ�?���i�����\��1��d��O�Te�����M.r4b��ʀo��'�rc��y2�|��ɓzviq7�M7BOI�%3N���'��6-�O����O>���[�I���	1��Ek\��Hʫh�,�$���`��ܟ�&������T��S`�"�p����.#b�LJ��iK��'9b�'�2Ox���O��H�Ra�@B�w^~ƤL���5�ą�S��<���?i�w_�F@+&���8O@�H! ���?a��O�'���'��'��3�	�O���p���,TH$�_���HI�X�'U�'�r�?ہ��?kZ�hr��9Za�4��OH��>������?���1S6R�BD�.Ԕ���L]:�����<�*O>�$�OH��+��B�?ə BR�.<`���ƚ� �<����?�H>���?��,��<�����3��y�3J��N2>�+��;����ON���O���$>�����C@֤*��ޤ�����d���	n����		���{~R#ڽ9��
M�Ggf��&�ո�?��?q,O��d�v�����ɘ �Bd�2�hH�E�Z9OW�e'�L�	������<'�`�'$��PBPCó]"B5�b�Z2
q�Iey��'1.6��|r��?�FQ��6C3��@k�'��=��"�<�+O��<�)��@""�T
��"�V\Y�V�?������'
��'1/1�4����A��O�6����\�q�6��<�������O��M�,�J�����pp���P�^���'��	�`�	���'��8O4�l[.1�<�z�%I��<�b���O�������O4�$�%�f,�VA��pG� +n���O��D�A}����'�I�
�nm1½�EN�$p��@#�<9�ʦ���?���?����D[c��"�a,*�6,�XN��	uy�'B�'��'R6O���QhH/�N�C�	n"��'zx	��O ���OF���Ob�'��ĭs*�{a�Չ%���-��?A��?Q��䓖?Y)O��4�R�2UyѦU�#1��b���ʓ�?���?�K~r'Z?��I%Q�5��În�6�K'$[.��H�Iӟ`�I��6��y
� ԙa���hBAN�8${�l�5�'���'���'�B�'��'y��'���E�9vK�MA�B�\m(MK��|��'l�ɺ_&"<��GV1��Sr �4�x�ɷ� (|hٰ���=#
�t����vbP`�
,��C�'�u�g�����(.�8�/k�a@�j�-�ēOV�d~�|�oڋ�?����?�����
T%�%�]�\�R�F;`��?��K�lM��!BT�CDfu�iE���!�6l5X%ۯ*����%�'K*Y;7������JBR��(q"��I��\8�ֵ�8a@��	3ڹz��͂9�H��AD�Da>Hp֡ %eZ!����6	l���g�m	"h�`��2�0ʳڀ�5���S�
_��[fI�	NΕ�f	#9�{*'	�̡;�eQ�]�����	���3�O�56>u{�Q8:�,1%�|���Ȍr:X�VH��yg����BϞ0���X�N�\�n�x��4s]ؐ���:@�ӥN@z@m�ğ�lZ+x��`�VP�1c�HBJn������H��;a��	�b1w*�Z��$�`G�,+����0��hA�!�Y�P�k��]�
SLC�{��E��EK
\�1�TF�=/k����P��dQ�22�'��)���>���>�8�)SČ�!��y�ъY�<Io�>˺0r��JFrp���
W�'��~J1I�5��8"Gΐ�q�<�h��S?���?A�F��$?�6�'�B�'X��	�h�Ia�
�$E���`�&ѳN�r�}o΍��a�����'��) �Eͷ#h|8�����`	������	W��i�Gh�3�I��sdn�\�(G�ˊ"%��Oڵ�!�'-����	��"F}��'@H�n)���$"Od�{G�R9[��]�!�0,�~8z��O4$Ezʟ�˓l���w�� � ��N�S�ҁ�e�I8y���'Wr�'��I�����|���&l��G2u��l�A����hq$cʡbQ��Z��B=��<���;U?���	1cn�A�/�r����Sa+,I�:%  ���<�ca�)���ʂF���Ф��'W2#e/�2�?���7ғ8P�
U��!䒨�&�#a0���aւ�;"�νe����Q,G�̚,�O��'��I*A�Z�ٴ�?����M��!C< iH�ؑ�7H����t��O�I����hX�Iß'��n]91��1�)D�z��ȫe呟�dN��Y��sŭ���鉝mQ�4KQ�� )Ð�b��߯gǑ�`�r��O��$^K���\;��z�(���RשJȾ��I�?E���@5rD�A��$[���8I�V6���ذ�)§'Ǜּi������E0����ᑡA�&�p���<�㡓�e���'�ҟ���'ћ�&UZ��C��]Qv03SB�)Th��
�C���HWb�* 
C�ԗ68|p��O:�O������9Ct�%�K�o�A��Od}0A�I7:+�4�)V&t��I��aQ ت`3�e�����)��d�䝅Y�6y ��F��$�, �	#�M+�i������O����	�t��=�1m3�xu�W�i�N���O���)lO��֭ضw��Q#��������ɒ�M[��ir1��u��dE�u�LU�F@��iq?	���t;�+�7�r�"&�G�}�%�ȓ!��P�����K�.��ҫ]#PZ��a�lΖk���tS<��=!�eZ���ŮH`YP1�'�Gi�<	�홚K%��c�+�;	�h�[�EOa�<Q�ԭL���Iޮt)\�v�GK�<Y�.��Y�T�a�i(D��̸�&�F�<q��F�0D�t��e�*&?�HX2"|�<�����{��,9w� ?=ܑ�f�t�<1e���!���2��5V��x*��j�<�AH������9���\�<9rI��M��Y�n�5��Q� CX�<�$*�+1�x�ʓ�Xk�B���a@W�<GdX�<���c% ;1��I��O�<d���bļQPIY7���I�N�<�J��f�X���1Di�%�Sj�Q�<�"��b�Εa�Ŕ3�6H�̚S�<��]"���C��e�N�+��U�<�S��yRy��@W��qB!
[�<���ҳcm�` 7�
�4T����Iz�<��ꕚ/�|�!�8in2���R�<�æ�=~��j���\
���A+�q�<�S���LY�ћ�hZ75w\�B�#�@�<	tN!P�, (�'	�����H�x�<9D���"�@ 
e�i(�倳	�y�<yr]�co�E+У�.�qp`��q�<���-2H��`�;E�X��5St�<� �I�����rNf�]�P���QB"O�M���4P�>�@W�L���s"O��rB	�(8v���n^y�����"O�壠�}�ZP�Q�H-�B"O�E�`�D5�h�K�d%��"O���dHޞP|l��l��ZG�eJ6"O�6i�
a�@�1�$�E).D�� ㌊]7!���O8f<�%a D�hȧ�A9/��ʳ�=4���!D�XUϖ����а��:w$����(2D�p�"3Cf|�gO29��� ��,D���pd�f2�9��Ɍ2.��h+D�|��+ܠ^ܝ��HF�k��];�m)D�,��f� Ȍ9A&C[�d�ʅ�ǩ-D��(�F�~Gd�q�oL!22(8�	+D�Ĩ#O-os��iK��923�"D�\���Ͷk9Z�	 ��M��j2D�� 4��T(�c���$0}*İ�
3D�83�&@7
�TA��.��`S�գ��2D�@�+�[��(k�)l�h�3D��0��E�S�fp�	}Shp��);D��x�NWxW��b���*�J��l'D��@RAV�t���І��CIV 0�O8D��(S�@6x4����(ѥO]D<�W&4D��bO��]��P�/�N^����2D�,�L'T����)�%�\LH�%?D��L�7
P�K"�ěn#�Q�,/D��S4��#B���s̅��۶1D� ���-<�IQ!@3G頔�
.D��Ib��.�d\��^�w�@5 ��.D���B��KQ�=��G�A8�R�!D�����]�t�5&ɛ�D����%D�����׮�1V��N|NA#v�#D��bÇ,�:�ٖ/����=*� ?D�\��L�;q{��t�AF�M���=D��R�d$F�}##.Y���Y�@ :D�p��A� Aƴq�Ԯ'��hpL<$�h��	�'b&�QC��y)�h�I��y�Gͼ-�<rU/�O�������y�%�63��f��m6d�s����y�$��t�
�� #J�� ����yR�VN�481u�р{�����4�y��$f�RQ���s������ŉ��'������I8���f�#K�b�8����1���x3�*�OXyg�P7*I����'�ȱQ��94�`�E���?�v��YXftZ3c�39��� �`�'��8��ˍLon�j��|�)�Q��5��o�dsA��(�!���2dN�"�n^��`�!�<�R����<U�u�ʀd�T����wlRA
Bg� ܂��f̾b�=�<��&L�`���d�*>�A�$�ٌ;�V}�`�U�h|����'�ݘӬU�TM��W>c��	��dklqA�`ˡ��*A�Ivu�h��VW؞4��.N�����FU�Jd ����L$�����n�~Xa�/�S��$H==�xK׃�+~':�z7`����)�7�r� �T0#G#��g^���M{�'m�)A�$
�F ���%E�-��'L��q�B�r������>X̙Fl[�%�*d�pμQ���E�c���y���6�(�(�ѣ
�	u��XP��'{�tm��dx�������;$8�W�_)Y\F�Q�go�5� '�
B�m��Z?�N�pQ
#�4��A��	�?T^hh�闤2��1x�/�z�X��U?�%��_4W��8˰bÛ_H��85�F�][5�3/8����I�P��=��ԟ�7�C�[A��H���E�m�I&�n̓�'7^訫矇O�LZQ*�>}DPB��.�uv��/[E�|2�*��H_�l�1�I��f�����3S�*\|pºib֐34�U�{8XʒŊ�BL��W&:E�H!�ǂ�*��EI�J�9����v��(=jPH����Ũe2ʅ2>������)?i֝0kV���!�V�V��bمZ�ܜ�&�\�U���[ �u��i�iN�������T��:,8��3�h�!� 6	���C$����v(�W�WHY��J�>@E`x# +�2�f�A%���
�����9;@X9
$س���3:U�J3V�V����@�<N�r�#�ʠ7vj���">�I �$�U'A/\ݚW'�9+��12͒(Qt��E��[��Ti��APe�,N�·'K�*��A�2� ��6��f�jJ�d]�<3t��q��0hצm��Eϖ�G|Bd��d�h�l�@<ᳰ'©9�� 6�I#oo@�xT��}(����K�`֒,ʆ�ċG ������j�0��FċE.��a���q�t���dH$f�q0I\�'�蘥/�:j0B�9�Ă7�0�D^������VX�K���f ���l��$!E>oX	) �P} a0KF/KZ�����C H�?]ʂ�W,3����&��+��[����U؁`l"P$�#y�}[��K�]j�9h�a�#L���:.^r���L�P�Zq�+A�-�|��#�T4�j���7K��˲跟�Pv��?#<��䜔,9X�`���4T�=��G�I�M��c��q�tHs��,�r���rV��0!��+�Hi.OkL@*o� a��x<*���o�}���	n�ڶ>c�Z	&	�0/����@�5��F�U `��4��"�o3�K+O�M�rlG�B���(OP��$@�5_J��f��#6��hZ�I��D��ˉ�Y�j�q�F�O��!I�t#�\����hi2�Y���8���iR����&'I2��r"�	�[�fi�e�I�|u~�2!�%[��[N���U	�B�$L-X������>��)K�3�r�
Gm�;�����Q�N-sWcX�v�x=���	t|}��ȋoL8��P�7e�a�7GVhK�!��B}�-sp�'���8�D5"�F���]
<�A�%�?CVL���u��C�4:���"���*0�ԥ�5_��	�j̨!�%���|�w��/?�˓{��2��KA4�:jP�B�|��א���)=��S�)X��%��CRJ_�Z�����)uӶMbB�3{.v��P�kk�C��)tѲy1�+D�Z���`�j�c�`�)qR����b�$�3膆
�$2�Ѿ*V!�ĝ�#9n䀥�Ȥ+j��Ł=U{!��ˠA�&l�1d`�AB�	!�'괜{w;dfn�c�G�8R!�d��p���X�X��ꊛF��	>�<��b�}��ԫ�� 4`L���բ|�d��o:�Ox��m�>k���c[�?x&��Qe�s M���X��y�#�3@��P{�|��Y���'�O����	d���&(�S�o�����"_,|�!��	^�Su�B�	Y(� @�h^�G�b�r��ݢH�jر���m9T��ny��9O|��+4d��M3bܮߪH�"O� �ԍQ�>�e��	��|S�;ON� �m��W:���))<O~q����cF�5x�Ȑ'�^=q��'D� �7
�a���Z��	���pp�&y�Qx����#���Βw=(�㦃�W�^�ၮX(J?�#5��#�b  g�G��x7P��$g�6`��@2��sV|x��w�:M���&R�1Õ/P�/��`hӦ.%8Ir%�2���s�d!��˿xB�=��� t�ՙ�m!D�42�C0t0H��M�>���q��~�㇀�'I��ڳI	\x�����=�1��3x��s"�<�O��!&o�=q�����A8�����.Rn�:����w=��h�S��yRe�k��e�q+��/$�u��aQ��HO`ͺ�CL5s�0�|J�"��y�NM���ʦ�h|xҎ��<��O�%z^�h���1j��Y�G	�	�I����e���\�k�p�A�,�!�?i�Eѷ/m�p)(��D����X�<��	:$4uj��2����*c�?of��c�%3씢}dg�m�Uf��;�d���{�<QĂ�(?�� �O��HΦ��I�F&P��Ӂ���	��H���	3l���`�G{�q���'j_xC䉖m��x0' D�=��m��a�7����h'���=��jJ�w�LL���D�&�Lx�J\؞������D����'�-)Y�!�z���g��xh����'��x��ʮrB���D�I�I[h0:�}��R�\ Wc�R�O'�T�2�V)
grDx�E�qF�,��'�epR(ܠ.��c��K�Za�,�&@��$����>Q2�>!��.
\��$�*d�X���_�<1ƀG�f�����ϥeRB�zCo�� y��h�X��Ɉq�E�2bF�z]HQc%m�##j����+h�Y�';�H���Զy�Lx
a�@U��i+�'��(����H:A�AR��ၪOLR�I������ܽkrPTi�N��(�phH��0E�|�a�	�� 	7��#G. ��ꂙ%��uy4
	�u�<̈́�8��R�4.�$A��-�$'|EDx��Įw&|�ge"i]�<��w�E,6z�E+t�O�5��}��"O� a�`R"0����;�<��V��o	2�q2A���S��y��?H�0���E��Y}�AHw��y�!��1�Ys�*!X�r9��y2�Q4�� �EkFaC�y�	��E�����ɟ_�ȹ`q��0>�.��5�(̲$��#z��DH�GۋS�
�j!턪G~�Ѱ�'�
���I�7�S�O0ZM���D*
? %Xfi��� �?}�%�R �z=SХ��
��!��$D� $IΘQ�Aڰ�W�tm�g �"C���I����	�p핧�����2vxH�G.����0�ҹ*&!�䛎{�%��NG�)��۰.�/~,�ڢ[�z��2��;����D�?R"6Ih�&̀/�4��(��| ":~�:��Ԉs�Ւe��2<�d8���iɰ��ȓR�`t�G���Z�3�&�����鉲4������BY�O`�0˰$Z; �.��D��*?�0�
�'���C2�M�|66l�ӫ��?���
�'?�� ���Y��)��U���R��yB@�(_�I�F,�?������>�y2B>�2�E�R� �Z1�^��y�c@�2yJc�k��J��PC��y��̱O"��3���sۨ�� ����y�n�[���!`��0c$\�`���y�̌ޞ�;�n��`-p���'�y�.}�*I�p�*��@]�y¡��TH���ܩ�
�9�ʏ�y�Ģ`��u%!�l�~Ib����y���i�l��8~.a�q�͊�y2h��2 �Q���6m�� �q�ۧ�yb�TnX����ԚcJR��Ce\��y2c��*�$j7��!K�h
s����y2�L�d�P����Sl��r��
�yrʒ�^r�ai�"_4��I��yr��2`,0�*���W-n�!�W��y�M�=D`�ժƅ@>I�*Ԣ��ybϻcʦ�sr�_�F-�����#�y�Q8x\b@�6��c���4�y"�=^�eavb��S���s���yr�M�X%�P,�N� ��A���y��W<tO�u�7���2F	:�y��/qM��MQ:��&� �y�Z�L�T�R�O�VР�!ϕ�y"`A�W4l���'�ډP!`J�y�
�L�Ā�Q�cX�p^��ybGV��Y!���=B0��y�dI�0�x����߂�F÷
�""F��p�l�:���P�'[�;T��z��J�J\tR	�'����mW�T8�W�ɼ'�<��'�H�2[�4	ׁ�3 2<x	�'��1)%.Z	?�,���`\��y�'�\=�t�M�5����%JӿF���'Q�|��� 74d���9k��	�'c���ċA�%��s�N�4l �	�'y�P`0�P��	5�ݦ,�Bݣ�''p����7>��XRCcR�x"ld��'�z-b��TA���1%��'�b1p��F9�Q�flϬ)t����'6�L*��7,@�Rfa#Jz±��'"&��A�֙29������Y��'6tq��P�B�!s��Ї6h�		�'��0����d�G�
5��Љ�''<�@` �p�`��f�H�>_"-�
�'厤;s�����VnX�80d�P�'�h�����S�h�k6|S^4#�'�@�Ƥ��;½��/�&T>��'x`@c���5,(��[�1��@q��� ��yg�,$�@z���R�L �"O�-���<U�����MśPO�{�"O>T�Q.��v�|�(���8�1�"O��遬ن\���#�kP��`��"Ox4b7J�Y�4P3�k&�2�[�"OTA�1�<'�|��H�x��	�g"O��R#.[��y�ef%� (	�"O��"~v�y0�F~MF�"O�xGoۡA9��D�]?'����P"O��x�"��1��)0V�ǥ92�B�"O�,�1a$ c�I+�x��"O���e��<nϔ���"�
e���;�"O|ѐ2a]UU�,�9��t�"O>�фA��ꡢP���^�*p("O���g�(>y�g�0�j�:'"O��a�U�e8�$�ʬ{���b"OP=�-�

v]�ы��K[�	ca"Op�I���S��r!V�nA����"OfT��1f۔5Å`\�[5�5�U"O����-ͣY�� Bb��"#�l!�"O``Y����w_�, ē�`p$g"O����SET��:��T#�m��"O�d(���1#}�$��̸r�"Q��"O.]@�`�	e�����2r�@�=D�(����4�.�XФ�tҔ!�*'D��ۀ��"�xr�k@J�X�)&D��S����4�rH�� �*h����M$D�|�J�\�&x�nۯa�V=Pv�"D��B�6P*� `#���P�&F?D�4�aD�j�0�1rK�7K:�ɰ�8D��p��uA�I����32�Q +D�Xz��>"/N���NF4w�.Kd�.D�����"����+Z�.�ܥ��,D����4(����f���M��G,D�0K�fEb2ֵK�B�(ش����4�I�,Ф��˓VXt�b��q��X6��6db&̈́��RPd%�1+\�b�@"��ބ/ĨMq�ۑ��C�	#G$e�E�D,�TMz�DF0�z��$.~.r)P�{B�I�g����K9OTf�8��y��U�p�$aīJ:,!��� ��DÊS�dx�{��	6|����$�D�h� hU!�Dֿ`���`g"߀;خ��T   >TqO�Lj� ]8���P�q?�	�ӎ��rRPԨ��5D��Sb�
-8l}��G�69!�(p��%D����
$�"�"�w����n9D�D*%�32�B��"m�
�6��.9D�{���xSn	�v�[.Z���)�l,D��J��Ɨbt�ga�K��1�W�*D�xbe��w��D�u�;���S׋*D����*A/��A�B ��F]�@�#D����	�V���a��^p$K'D�j�/1�lx8Ĥ[:�1��#D����$�~�ђCؠ5� h�,D�|P��.�9#w�ֿ�C��<!J� ���H�S�$#�^��R�R�=+ZP�W�
��>�Q��>)rh�$VS���e�8*���Gˏ�"�6i ����O�9@���&5�B�c�ؼa�ؓ�鉌O:��Pvn�*?a`����8B�(��xeX+��V|�e�BݕEH�X�S���&Ӡ)c�oO�p=��Y7R��*�mˁg4BQ�mզ5�@��33�4l:��^����IO�(�eۡ'�R4De5H>���.lTI� �$�c�j��y�NL�Gh�3KZ"��|Ű�~����y���9T�(`��.�t��6GBrJ}	݀��T��.)�zt�2Mi� ؑ��D'�p>fKZ�s]�T:�G��]V�+�+�C���IϻS���y�aݜB<�	9��9�g��w����]1O��;wm���R��&��2�%i3�I�V.�8qa��c9��� ��<rj�$k7��3W� �У�a_�CŪ�0r�$W?r��2lZ��$9P��.c��Ap��'���d���j�^-A��
J�<@Ehƛ.v�8����"4 �͢���34Df��`���*^^,C��<J��=BA`n�>|H��֬m��Jc��x�[!"O LZR�P�5Ѡ�,�- ڔE���WnX-����FԒ1@ MXV�ʦi�M�[�؉X6x�a��$��U&e�!�qW��ˤg6�O.2�E�lE�2M��3�
ы���_~�ڗdO���|9Ѯ��?���Ǐ=��e�4AٷSm�Ј���{̓o�jܲ��G�	� ɶ�O�4�-Fz�`�1�����D�d�eX�]3ZK|Q�ƿ-���q�]0|�Â�ի0 �ن� Y���"�Gl�X���I;��"O2]�h���!�'���	�r%�ゞ9)ڒ�st ��z�vWW���pC˔M	l9;��~��Z�G n�fdh�́�+ P�q�
?D�`(�� pmΕQ�Z�x�a��K�j  ��T�1�,�J��(��`*���ON�W�B�d�(`��Gz�E�厏� ��5��ߠ@>��G�9�O>��A�A$9.x��V7]�f4:&�I�2�*|	�� ]>�uҟ'2�E)ǦҷP[� ��N=,f58�}2�;pA�)��ɟ�pK"[?��D|2��(��Ň��ΕA`��]#l�S%P
Zp��!`��?4���J	����9P���G�'p>=���P�2�$ �2��x�'l��֢�C���)�I�'�><��Lm�0�,��y�O,�m��d�-5\�؈�h�&[����'��yY�� i�����8~<;����� ��8O�s察�o2~��'BܵO���{썒EK^-j��f���2���&|�|�#�M�O� mۢ���.V�����d�f.v�ZQb���Hh� [Q��bq8o$�I"kG�>���zr,�(`�d��/��]1���B��p8�e� 9�
�%�>�|�����i�v��+߉0�R!���*%e�P;m�/@p|9�Y'[��˓A? ���L�$lp!�BY�c\�dYt��ʧf���H�?]�4��MW�o�޽�ȓF�5�$��oRQ&��$I$"�i��I3°�t.�3���I֡	HEȟ'�D��W�H�W������

���'uD��I� U��	Y��ۍ�(�8��>�D[�_��ppu�٠H�Q���⌇��q�@D!^�hr
7\O<�'�N���ԻA���"C�H�;/�`���=G�R Y@�rTa2�<� c(J=|�슔���O`l��+ q�����TN�-��	s)�{�Di�0��y$ބr�ҙ��B�P%!�B
��Č ?������+����*�"'��T�v�C;�B�	�iX,��^�(�xBs�L�k�B�I	]72aY�'�d�v@��._�ZC䉚����@�>�Z,�%eڍj�C�I#Ir�d��H �FH&�y֯�t{>����9
i���!Y�����%6_�i��Ꜣ">!�$ݖNMȴ���ӊ"���C��F�"2���R��yj#|֍�#Q
@@��i��/���x��J�<1PhZ�FY���g��-u�0a�����<)%ێy~���<E�$#VE�F 
�d��Me,]!�#к�y�h�"_���`\�@���&G�������H)�w�'z�HZ�i�"3Nd��ۯc%n���b���G�>�X@9r#��AΈ�YrBۖ%c�L�ȓC��8v�ՌH;ry� 
�S�2MD|��C���ډ��	g� K���?5v�U��!�@ Pԛg�[�|W�DsBÇ?�!�dE:0	�Y�R`N�%��,J��gN!�$�+"�UY�"�$5�^A���),>!��O�'$*���l��5�
�tH�%)-!�$Ѻt?Ji��C�9��D�&�P�0�!��<T��#���D"�q��hޯV!�d! �Jt!��#��'H�PQ!��P1f��������̔=����&D��j�ř2޴Y��D�W���"!�%D�T@�,	�)q-�z֐�X� 6D��bEǙn�xi '�L_�$���
3,O�ђ�N[̓a�&ɠ�hPp�6�O�f6�i�ȓ#a�lr�%�,U0���H[@ԕ'�@��)��ا�ONBe�"N��.-B`�?0���x�'����]�p��x�$�A�x��}�CF7���]���%��b�#`�t�2�Q]�!�Ģ;��Y&
^jܻ�fY��CK�\<� |Pq�[�:�F�����*p��%1!�'�V�ˎ{"�+<�(�&�B�iD�qPđ��y�HZ>?�Ё��&x2(��C�yR�FuHI��$ t�Hh����y�eɒJ��Ⱡ�#o��i#�R#�y���
X�ZesfKZ e��Ms���y"�B�n�2!�A�ψ�bՁ�+�y"M	w�P]����5	�Y�����>�G>>'�Iba�_�E�@�r�	6@��Ȇ+Y4!�6�t�T(�p.�ݱ���&(���`�G_2Xj����|��2E��{I�K�戃y�!�PSR�8a �P�H����Boy��JK#+���K��s� 0��&W�C\!�q��+E��'�B��"`��q���-؃i�T���O$���F�l�lSϓ<��]ȃ玫sDL�{eJX�~݇�I�n��C��G����M:k��(;�A"�@0�'�z��U�!��T &�Q��|�Y�'�$���˸g�����3�`b�'�.�k��G�T%�Y Iͮ%h��
�'�	��	^x�,ȓa��#/rY*
�'p���l��c ��L	�&� �'��u
C���hwL����=�@��	�'Z�t�v���~�%�/j@�};	�'(x�j��F��:i�bO�J��j�'�.lbu���;c�}j�Ë�r��
�'��EÇ �,gh����� �	�'%~��-�G�^\���3��H	�'������7H1��GMq,�{�'��lB�$Q�'��i"'���'���8�G>UvHyDO��
8vyQ�'��d$WaD�8��ً�����'��}j7��#x�>��*��tr�0��'֝�5�۪I�M�aꙚo�j�{�'�Y`A��� ����n�@ɇ�z���B�Q>k��p�+�1\��T��#J�U�1�A�;�FY�ǭJd����u\3[P2���0� 
��Єȓ\��ɓ="@08q�>w�F���h�l!�7adM�X钾r0���ȓH��`x��D�����jN91�f���H���Y C���!��;']��ȓ?�=��lɣ\��!) �9H!�x��6z[�Z�hN��F�ڼK1:4��p���T�P&i��!�Sj��M����ȓ.fŻ
5gٴq�t��p�P�ȓeY�!�T'|e�YUDě;>nX�ȓl������S ��d3"E1PE���[+�`��㌬0�H�`�M��1�1�ȓ[���Yӣ[�{Z6��0�;?���ȓ:b|��䈑&d܀aDŜ,�*U�ȓyؔ�����'>�"�;$�]1����ȓi26�A���> ��K�!M�{��ԇȓz�����\�g2�	cc��E���H�VЩ�̨�,0b�j���ȓn�#Ɣ�`��=���E�����t}k"A/�� �ˈ�-{����j,�Yw	 4�u��!D�GL�`��Ӿd���h��$���REB�m�!��?qw j�B��,~Dd�7k�B�!�Ǐ\��}A%�@�Z �)�ȅfj!�$H)yp4�q,� P�:�BGJ:�!�$"w	t��爒�b��m1e�X�!�P�,�FUXsn��h[aKG[�,I!��9q�l�b�3Fp�[�e�4�!�� Hl*�=R1b�т�f�<�C�"O�;E/Oo |��C,	z�,��"O6Xs�j�jc��Bf�Ši���"O���jTq�"x#���/t9�|0�"O�tӖ�|�����;��
�"O��Q�@�$v����f�v�c6"O�Á�Ө<�i�¤�!N,��"O��B�F-	)�=;%��EG6A¦"O��5+�A0Р��э,;��*�"Ot�VZ�6�C��.u[S"O$u�@�������Dn���F"O��j#e�+&L�6�O"T�踪"O�Qf���Cm�=�!۷_�ѹ"OpU�D*^s�� �T��-Ht�R�"O	�g]�T�bH��ơ77�[�"OX��G����s��`) �²"OpY�dES�l(�b�?."�0U"O�h�wd��N��7�*u`:�"O�1[��('J5s��Bpn���"O:s%h�c�D$�d��{P���r"O,<{�EO$@ Mz����=��b "O�Q���Y�u�\C�2x:nx��"O89�Rʜ3&�5Ue��.M�"O4�[��6pr*�T�	�(t!�"O@@"gN8��y�5�T�HB"O�]0 �H�W�С:����a�����"O�X�%`f���=\�(���"O�X0�$څ[�R�:�G\>H�vLq�"O栣�G�41�2�&�4:�\�"O�����څ
9DT�0����!�Ě�X��T[�0aWvU�f�
�!��7~LZ	��+�,W%��J8<[!�SL��AN�VU@�K</P!�?J��h��MލKĤ��rJ��!�B$m�  ,�L��@�`照q�!�P0#�:a�-�>~��r�E0 !��
h�ʈ�T�~����G�l!�S	�4REZ�Y!��Mg!�DI�@̼䡶舤|�^��E%�$Ik!��~��Q� AC&	Ӥ�]!�#��\���M1
 �fC�	L!�D��$�j��]XĲ��%�\�6-!�$�B�\5)AB9�~�"��ʇH!�Ӎm�n��͜JH�q҄ޟ@+!�G�+����)Ý3`�d�,!�dݠbށ�(�E8�CBCE�#Z!��زIT�AegS�J�&I���0P��NU(�%�oD6�Kb�G.ij0����� �s��$SG���$�E�ȓ�r� a (p	�5���NY�ȓ�J��	Q�m}���M�7�4U�ȓuuF �FIO�\G\)
�o\�'��a��n_���	b�L�MY�i��܅�'n<S�υ*��k��S�u$����l�Z����K% #�1�� �;% HІȓmV�Pt�P�@a����I�ȓK�	J��_+E���aKЖg'�0��Vb��G!>1T���>0Nh �ȓ~��9�ҋ�,@��!I��E�ȓ" R!J�ʌ%L��"��� ɇ�m2�( A,<4��\,��T^���FN�f̂`"�e�E��ȓ��5R6���ы�E�z �ń�����y��&�P|6%��S�? $4������)v���];��bG"Oz8@F�)J�h�Dͨ:}�!��"O�sĊ�mҰd2�2v`1�"O�S�j�Y���h����Ҏ���'���3R'Ӿ�uS��/̨ɪ0M9D��jA-R���Q�Q���P���!�b3D��xtAј1��{@+ƼR����A�2D��d��5�=��"Ȱx�^5Jgn-D��0�"ݙ'���ʷƨI�Hi*�*D�@����p���qe�"\�.�)D�lS��%䤙ʁ�b�ʷJ%D�dۂf�(�
�@�OZ*'rؚc�&D��+�B�9��K��9XW�P s�.D�,s��=8ݲA��R�z���j%B7D���M_1k��B3bV&^tb�4D���w�б)I>��qc2(o1D��lD'�J`��? I�%��_�<Ys�'0
f�J􀅾&) $�b��ȓyD�d��?�T�1�	�D�ҕ�ȓ<T�3�֋UZPYb�!R<�
}�ȓu�L����Z`��"Ԅ��$\��ȓV���Hp(B/�q�3��=\4v���24I�q�IlM��/�X�ȓA��b!�
'U4�1�AET=��Cbe	'a�L�� -nV]�ȓ�za�%f�� ڵK�)��|��8��e�\d��On�:D���T�ލ�ȓC�����������S�Q>|�X��+p*\BկB���X"��>}�R\��c�,Hw�L�t"Y`ň�`�@�ʓ}evm�f@^D�@��#���:C�I  ����S&Jv>��%$I�C�	�p�lT����@��-�WA�,��C�	`�q�-��E���vf�>x&B�ɖm)nMp5HΜP~��ұ*ӿt�C��3��)�*t�NIS/���B䉭8�0\i��]�(�
U���-� B�	!>����.�z� ��ID�>�
B䉪'���#�ԡm�����ˁ� %�B�I-/z����	�:6�I���8e��B䉱"��ͩ1�X��m��&ǔ��B�I����:��U+e�M�#�� Q��B�ɽ�R�o�V��t2��N�~K�C�����▫�	R�ܴ��/��*�C�.� ��%,	�^�t!%B�RC�	%Z�: S�3�n(���"4UxC�I�w�K�/�5H�8��-�� ��B�	�i��p���\;8L���6	Y+\�C�	G�(KP甑4.�Aa≃+��C䉺C/�y��ŏ�Da|C�f��}<vB�ɐj��)�1K�5k<1@�/��-B�B�"n�	�f��/����	�0|B�;-�(�%��32�C�ņ�0��B�	�;>�"��ŉW��Y��$��B��, �)�홛E����V�)Y�B䉭?Y��	P瑜-��hQ�ݙw��C�ɔ/��I"c���#��f`݌L��B�I7�2�`��] �9ae,)G�*C�I8<��v� 
!�m;'Z�:B����}����N���`Ù��C�I#qyS`�j�Ы�bZ�ZU�C�ɯXT�Wm�~��Ybv�� C�ɘ;]�r�G�6Nֈ1s!H�3��B䉥ZM@A��+���c"��0�B�)� �vQ0>�3��^�G�>��f"Oԋ���"�9���șK�6�Z�"O����mԖw�D���
o~�U@�"O�аq��!"1sv�<f^�5��"OL�+GËA��Ke,�O�W"O:Pzu����p3,�-���"OҘ��퓾|1@Aa�
ӹm��ś�"OL3�'�Y~�`��_�yz��{Q"O��H�`�1z歑$�g��!"O쵢�@+du��*M�U�q��"O�%�#�Ֆ`dF%�O����"O쐁���I���q� �4o���p�"O~l��Ŕ�8�p��nO�>L�x"O,���K̻e4��rnD*V��Q"Ol,�a&ʗeP�L)�l^��>�!"O���5��lj|,S�K�q���"O��Q�!I��е��"�"ORUÖ��(n�2Ɂa�C
*�:�C"O�=�T�H�x�F��Dd=�$t��"O:�� �R�o�����	B�Ne�t"O~�S��
,/�&	�3ⅵ����w"O���V�A�4|EA޻d����f"O&%A&lA~w^,��O]��t ��"O֠�� W�`L�M ���*J<*��2"O����&� .�q �%#&�]�"O�!��M�#T8~)aD���,��Ա""OP���uv źF��&,Jr"O�%[�y��&V�b�"O�iAk?J̜��^q5��aƞQ�<�6�۠S����aMF��ye�B��/gˆm��*�i�d�"��*K�DB�I�rrDܳP�X�'6Y�G��!F��C�I/�|�`��O�pN*!)&�B C0�C�	�dt|��!$�H#e�ц��"{�C��,EQ|RRLʦa-Jh��"R;{sTB�ɮ`*<Qy���/�HP h�!"��B�I�@�
̻�/8=�T	�b͜~�BB�I�m�Q�T!^+D�IPi
P :B�E��9��j%v���_�\7hB�I�=4�C''��j4��9���0:B�I�C89఍�Li���5LZ�vjjC�I�vT^�Т�W��ܥb��V�� B�	C��e�aR3��љ�MV���C䉶>�|�y�o$j��@�O$C�I�i��e5K�(Eh�O�;��B�	y��싷"Β)p���M��7��B��1b2t�2��*lL�����M|B��< �r�;�m��vp9d.�bVB�I�I�A@c�f��;�̒-ĔC�	8y=0� Bb�&������
}&B䉚k��$HZ�y$��
���?�`B��I�>���J	?����'�@�%��C�I=!�,�
�!P����#��`��C�ɦ+�#ҥ	G8�ȴ-�ʹC�	�>%����N�H�X%���N���C�	�m�� ��2��&PCI�C䉳s����!i-,��`X��+�(C�ɷ;���3h�Z����ڰvN`C�I,�61ԏ��4���X��p;>C�ɖxt��J�)J�k'���X �>B�	�R0�,`�O�F
�$�N՝e�C䉢Bt�Sq��(�p[��GG��C�I1C6���i�_�\ k�>dvC� ¬EXu�8T�`�u脰�C�)� l]�T�� HjU��ᓋK��9�"O
M83f�5D`� S��٥(���T"O�%A��W�`=�X`�݁v�Z�"O
�K�E�k�,@�
L��BY "O�LC�Cӝg��!�L°τ���"O�$��똏pjae�],���R"Ox8�I��2�V��tע}J+�@r�<+�+LvTIrP$�>���7��r�<9⃔�c���ؔ �zl����B�<!�o
��|	ئ��_�`��X�<��B���e#�$��t�D��x�<�c�Hp�|劶[�4�y�Q�Cr�<��fY��&8z�h�Z�f Ѳ��m�<At�8JP� �W����&?T��b��B+v��Be���h�T�3D������S�91�J5[�ʼ�!�1D�0C�M�����Ɲ$L�T`�*.D�� ���;� ���*V>WєpE�+D���MߣRk ���G�.�|���O4D�� 1�7
�P�J��޸d�
y�=D� �b̂)l|%:�꘿Dh�� �I<D�D����	f8!�� 4�V�9D� �f�#N�l��1A�
n� 4�@e%D�1��ުg�2={vHT�m� \�C D��!�P1V�zia��7��平�?D� ���W�/Q�$���6Q��Ѓ��=D���ů�*���3@��W|���n:D��+t���U�B��/D!�֌9D�xH�*ڕPH1u�[�����-D�ZwD2=,��f�ʯ/R��'& D����m%W�:�c�I ,,���4L0D�(*�텥?�򽠲��U����0D�!F�-��J��EKt�z1�+D��s��B�C2��Sk���`�k��*D��6
C�ri�}6�S>T)r�`�%D���DΛQ��E#��о  ��g�'D�p����\g�y	�.�l�W�#D� f]
�j�m}Єٶ'!D�D��#�M���s�'	�,�Ve�%�$D�x3��ȰH�H�1@I ��! �"D��JgB�Q0�0'��p
(��a,?D�\#@H _�"��E�̭	��Rb D�[��/��- �]8��u�7J"��<�w!�x;r��փ_�=�b��c+�B�<���<^�(+LT�o�4�)�j�s�<نmU	H"i����#x��91��o�<)T,��p,�i6,�*4�l����g�<id_#`�)��� @���HHD{�<�,O�s\$��1��I���� ��P�<iD�D�>v�0��狛A�V@#�n�N�<����0���I�O����9s	H�<	�AǫL��X�2f�)2nM
t`�G�<��AA�3�q��E�L�lhc�\�<�!V2P�d�F���)�L��a��V�<��H�K�P󵩛f�z�"�W�<�#G�6AiX9	С��de�"eTV�<)����j�Vn�G}�X�S��N�<��gN�	�4 E�s؎���eI�<qTGd�V��c�XݐQ�ƌ}�<�4�uj����b߆� A�Cw�<�#^�Sޥ�q�ЦaJ��ԤOX�<A�b��f�"�VND7_~]R*M[�<��JN�2���r��!O�1xT-�P�<�0�]B��Q��)9�ڬ"�'P�<� ̱���
�+S ���,]#y��,�3"O>0�dLсG;@3�O�^� �A"O`�d��,���D��ܸy "O-�6)�F�(؁���$���U"O=��.{W2� Vʆ���,�w"O�$�pl�&ϔ�TdP�r��,�v"OHar򌒢����F6�<�"Ot�k�H����y�+D5��l�g"O,�(�HЮ�F(S�M�a�Ѕ��"O.�x����"��<m
&D��"O¤څ�ѽ��AH�L	�S����"O"���P�C� d`#I�D�ȥ�0"Ov�C؂!}B� D�Ѭ@u�$"OhhY&��?�(x�`��3�<z�"Oj  S&��6��a�׋2���
1"O�h(Cʺ*��Ő���,at�Y�"O���RL�"EO�L���50T����"O(M���:����P�ͪgO0�@�"Obb��C�qw��� M�Wk�$y�"O��Xg!Gp�|�9#��>K,�1A"O*�����C�:���J�1m;��"O���4��I������#���W"OF0�g/΀�$�dO:+�x�q�"O���b���3bh�I�+o�|0%"O����?���a�`�!��)�V"Oly懽x�`P9��Z9��ҵ"O��saG���.�+l��`"O��`��ϲ4�l,9����[��	H�"O��p� �jB@����BK�"m�!�Dگ||d�����Т L�!���n�Ǣ�T�����kM)a�!�
7�Q�rCF�jg��0�A�a!�ļf`:�;Q!�YZb��C̝B5!�T )⍣w�R7^���(X'!��@8ֲ<�d�U�$?��a�N۽!��V!�8��Ņ�4>9�9)0+	�"!��U�4��P��#����#Z��!��!#������<ePv��P�$j}!�d�q�¹�)rN�\V��"@y!��,d����%SM��a�螴 y!�$��t���0q�NL����fV�o\!�$M9FbI�F��]�Y���S�<AfRE��5��"��6�ԥ���LJ�<1Ҡ��5�vm�	%Hh|�� E�<�0 �/\����Q�ًl�r8�d�A�<IäHǶ�[�Fؾx�䛦+W�<�$OD�'E�]*7��5�h�ӲF�l�<i�(��>ܒ ��� �9'
��w#e�<Qn^�*� �X�څ ���:T���g�M��b!��߁Q���%l)D�D���2H̘D\%/Q��(D���[���͓O�>E��B3D�x�G��⠬��I<��B�+6D�0r�F�8n�>(��Ŧm����D�3D���&�U�bG 5�v�G���p��1D��1ͳf�&(�u���,��|�H0D�t�!��(A꒤�9"F���$.D�营!?{\�Á@F26�l��*D�����^��	��b�P�����X�<��̩flXcpZ��l*r
�X�<�BO�M|4x���3�1"��GW�<��e�!�ޤˁ���,,DT��FQ�<	�"�&��dP�@�:lb�x��,�L�<�g�=O�Isg��;B�<��C��m�<� �Xb��G�8� ���.\�r(��xr�'���U3[B`4�#�g��x�'&,x�S�V.Ԩ���9	��8ڮO����`\� �AlH�~Kj��2�H>��6�>�M�"~n?N��邬�.0n<�{'�+�.C�Ɍ1/
�uL�-&�r�@���C��=0#6�Išò6���@��@"O�����-*������'�H�R"O��hTb�p~蘂%щN�ܸ�"O����L��fF���ĕ8 ۴���"Oek�.<`Gt����~�:Xq%"O^�ˇ�לT�x5�۠YXp� 7"O�ɓ�덝R��L���\�1OP��"O��FX/+&L"�X0ZX��"O�3�e7����� ��D�(��6"O��Qt%\�zO�š��B�Pй�"O�8c�a*&:��R��HH����0"O>��s�M3
@)�e�f4d!��"OZ �`kA<nT���,|��"O�R�l�aNy��!ӂ0x��ڳ"Oj%�Zh�r�V82e��F�Qb!�ۢi����# Q:��@��f�k�!�$�(k�6��稛9i�<��tO"C!��#;�v4�Sb�/e����O~I��'n�"� � ��x &@�$l2��'�X�`��(	���%L
3- i�	�'z$@�$.|�`� �� �(���	�'W.H����,0疥h�k�&r0$)�'@f���X :0�P� ?L��a	�'˜q�#�3
�
��2��u�|R�'ުI��AтFʦ��b��>pTΉ�
�'�\�P��%dUb+Q!���I	�'	��y�C]�Z�LX�Q��X�X���'�ٚ�Q�H:�1�K5L~R�B�'��,����:4���DMD��X��'�V�zgg��"����r��&0\L5�
�'
�%��ㄲ]�Ps�!�$^{N-�
�'�9I�8�R�x!RWQ��1
�'|~��<u<��9�hXO�
�)
�'�8��7H�-#����oǾM���2	�'�:e,`|$�Z!.ԭG��z�'��Y��\�m8t�×���:U*�0�'Ƽ!�3%��)sPݩ�Mט{���R�'A�w R�EqP�	�Ʈr�n
�'�P��G�.:^({ӊ��n�Z� �'�Șs$�.l�0�2�ȸR��u��'霨0�7��0.�;� ��'���s�Ͷ�t��J���9A�';:x�5���
$�ŬҩD8V]�'2�Ч�]�|,�/��B�~0��'~`E˴f $�������'���kԍ���LB�ƕr�6E��'��SF��o�L��U͐^N��[�'��D�Ш�-�I�a��VFޝ��'tvX�W'W:G*]P!�{�Xp�'�5.U'BA�УX�>��=��.�c�<���1ly��r2�O�u�P�15_�<!��B"��S�܋��\1I�o�<a�"x*u݆!.�s�/R�<Q&`�-�0������h�*}k��c�<��$�	C.�A����4(�\ġ�ND�<9���'L9� Y Ƴ=(�	RC�u�<Y��V/#� �Bɑ-"�ʙ��}�<�7�n������e����a�<� ���ɵRh^t8È	�>n��w"OB�8������	�<���c"O�5�c�;C��H�CЀ�C6"O
ݒ�Ոx�r��g&8���v"O�`邃~X�Ks�Kg��a:�"O*��֠"j���:$(�"O�!ᑋϤn}
�fLZ�G
ʘh�"O:�1�A@�N)��j�	F�M��: "O*y@�X�԰略�l��@"O؈��R�����_���e"O
h1�
�<U�F�s!��;Q"y��"O���ǒ_��kť܊SJ����*O����h�*eDD����<��
�'}6��𧟼�~9��. t��	�'^����43�t���^��bղ�'�a �c�zW8��C�̦��'�
�;ì�	��$	t�M6���R�'R�� ��A�5��!�NL?Pb*�'�J	�GJsv�0� ��KZ�a*
�'��Z�M'o��Q ��4=�^��	�'K<�J�m�� �8X��!�:8*f�C�'~ݐL����9��م7�؁��'�Y�C�ɏW�`��F
*&4A�'�B��e��%�rm��h�(����'�x��>_��A�ٽj6��'���
PM�0d`�e�x��x�'|���0g�>h�5k���$U��'>ą�7d4�ԭ�ħ9/����'�Xi�CB�I7�k!��&���*�'�J�;�ƍ:^�TU�q �� ����g�~(�r��"J��9�aɗ
fH�ȓh�f��whХ1��@�&d�rA���ȓ��!&���v/��l�+F��̅�V��H����� ^*'@��7`�Z����� �*�-�7��M�ȓ�ֹ��/Y�r��P�3�ɞ?^�E��i�6|H���q]�hY�*@�Tݞ��aM4�rr��L�T!鄨�!y�نȓ�2LpW�H+*�z���B��
��ȓE�H����!!�ҁ��C8N��ȓ�<IR� 2H0�,h�h���"O(�b�F�3P����ʅ���"A"O�Er"�Y!D}�)P�K$|����`"O�x���_��J� 
#w�`4�b"O�A�&�8y�̙�W�M:)��u�"O�`)��/R�0��ꎔn�Ґ�1"O�����$�J��zѰ�J�"O�"�f���q(ȾZ���"O����e�� �%Ɏ�v���"O$Mۃ���R�N;��C���"OD��N]	]@�гh�.	��9x�"Odع��5^�p#IȻK~z�+E"O�Ւgꋙ"�UcG	�CM�p��"OFH�ъ�V� I�/�EQ�<H�"O`�H��\�:v}�.�]bD�Ѕ"O�xC* �5AV��ä ��s7"O:I���:N�t��4�2<GЄ�g"O���1Oߓs���veؿs(�! "O�a�eE!\yH�#'(ޡA�"O褒�ʂF�
9@� �N�<�q"O~���,O��D�ҏ�d�Y6"O��&"�!*x �e��W���"O�\b��З$4��.H�P1!"O�����Ș{�Tm���M�V�x�"O� L�0��;S��ݑ��֍-�z��E"O2Ԫ��� �t��sO�*Ǹ��"O�,�c�wD�ha3��I�"Of���B��p�`��#���x%""ON�x��+h ,��W�N9n�0�R"O^t"�� �S�.����'0��a�7"O^Ԃ�l��ZD��f&ϱ^�0 #"O��HL]+t��`2Dԧf���J�"Oؙu�Y�b�VE�T��""O  �	sޚ�ۑo�9�Q�5"O���/��CB~��G�X��x�"O��`u)�*x�|p�,�Zǂ1�"OZ��*z�*()`K�(#��(Y�"O�)�K�W� pDQ+C��j�"O� Y�o��]\��
��,A�`���"OJ�	�����`b܉#��р�"O��ӱ�[����oK&>��y�4"O������Q�4��{���"Od���͒=XHɢ"$AFt��"O�����,R��q��"�a)�"O�b�I�X��t���Ќ���"O��B �>(>�#-��8�z�"O�А�ƥK*�Q��� �2�B"O|����+P����,��'���ʢ"O¸�e�S��{B�2N�v�I�"OTAPr�L�truH ��AY�"O&$�s��00�!�e5}�m`C"O�p����>c%��AjжoA���"O��+���2\�u�5J�"�m��"O�=�f���JXp
�>jْ�)"O�=� $p�T��B�J�M�"O*���ԲU�X���a�H�ٓ"O���p��gjl��f�P%l֤�`"OJ�y��	3�A�v�.P�D�9#"O^5P��U�%Bq�waƠ@�\�H2"O�`S��J�-�.L�C��P�X���"O��0d�7���*�/�35Z��g"O���ׅa@�KN.H�xw"O��0���a� yd�A�"O$0����&�UFݾW�&��"O�Tc�lE t���e�P�65c�"Ob�2�C/�a�NǚC��Q�"Ol1з��$���$K�-e�t�8 "On4)TW�9�����.4�,�"OZ�����d�N(�Pd**6���"O. ����=e���C@�L�x'�H�R"O�ҥ�"`�RQ���4C^�@"O�dh�IľU
Y2%��'�x "O̩�wa�Q?�y�n�#G\�ڰ"O���N,T?a���.QZ)t����	@��<[�%T�9��ʟ��P-���:D�p�S+�`X�#�@[�LAKW�:D���R�C7n�1(�Q=92�"D��ʶោ}��mB����V��2է%D��A0$��f}p�x�GK!���TO>D��h4�T�Z�,�Rb�Rkr%j��:D�Ġ�M�)n��kӎ�vmX��=D���# �/Nl�7��=�0e��&�Iz���x���9���E�&����G�?D����d�� Qd�@��vT��Ao3D�������6��2�(�<,�;`4D� q@J<Q���iF���>G�)9�'���D�|c�-r��KB����
�'s`���Ȅ,AB\ё��!9Gδ���� ı���Z�¢�+v4U���<a��4�p��2�Շx�v�Q�`��Smf#ǘ�8���JN�b���?J�*�cD�� '�B�S��]Y���KB`�P�)2pC�	�d���9$����|�b�i�sOhC�	.?��q��-a��@���;@BC�ɀ@=�a��|5H�iRjX�fY�C�	{��]"D �
s�����?�,O:�=�L�pxe�X:4�b��e�rR�͓��?�%���[�Ni����;7�2Y�6"�T�<Qa!��\G��B�K�5#���-LS�<��!�������= }#YI�<�2͜)u���bG��fB�qC|�<a�%�L�<�C$�1l�^�B�p�<�ǥ_Q�ə���.��=�`�';�yd�oX�	1
֮j�Y�dKgt��Slt A�pe�-.!�aZ3�!�$�����c S�^�ʍs�R2�Py�Ȏv�>t3rAI�M��4��:�0?�)O~���A��Vp^T��6=L.���(�S��y�%6aY�����5,
Ή-W�֍�ȓy��E�8~����P`K n�ȓ��lI�I!Z�� ����\pD��ȓ �Z����K�y5Z�o2
�� �ȓ"��d:�j���U"B�\.Du�ȓl��ȗ��*{��p�`ʕ���}��D�t`���,"��S�/�&&$B��cH��g�[�.��"�;(�C�Ɂ5d���-�>��!��B�-�B�I���5�� �	 NC��hO>�*�%�"�4�`b�N�\�i�N'D��&�ײo��y�- �D��#e$D��C�O�d.X8V���C�\��� (D��@���5�z�Z�Λ�c�Py5�>��T�j��A.ç(��� �aI4,G$M��S4̼XۂQ2p�pR)�.>f���hO?�a�Q���1[���if�6?9��������EL	(5�9Җ�^��@!�"O6�k �\'bfD�X5O��4��"O��@�a�3T�91�͉#{��#"OZ�AEB0�*�#�A0 ���1"O�01�	�Pn�P���wLy04"O"X�3$	�ZXv�9 c·T<-�eN/�S��y����/@��e9�p�V����'�ўb>ѫ��/]T��R&-tI" M;D�8���,f��7'�>���DLx�<��� 2��7�:(���g�I�<�fZ[	>�b�,��� I�J�C�<	(ۚdv���vlX�9�G�A�<�уY�p�=h��;ԁSQ����'F�𙟌�r+�>zO�yI�#T�ՓA�1D�Pq��t�ق'���tҜ�j��2D��{��Wj!�1�PEb=FK1/D�0�$H
o����+���0��,D� ���s0�8�R�fE$�<D�8��!;�$đ��[$D!���:D�\�⦆�k�BS��.{/���`�:D� ��oK�P6@m��2@��1�7LOl�H�E�+� �P����^�yB�s�Dx��mL�'�� ���y�V
T!��c ,H�P�U��y�L@2Kд$���8�d�y��)�'x ���TTH�c�"w��A�����m��QP���8��Ї<tܕ�P"O� ��;V�ɢS�l0�Ԁ�r����"O�`��!�>O���-˖$?2��1"O��V/��f.0�g�M���u"O~��(i�N���k�n�P�Cs"Or���VuD$�!Lڏ^��yI��<�I>E��'Ī�q����r�"��e1X��O���;�)§#���Ȥk< �&m����Td�}��Zz욤I�/J��
���n�J�ȓ<� �cK\��Ij���/V���Q��H��*TD��!���"2=��/,@�sRaQS�e�1�XNK ��ȓ3,><3�O�D�iY����jH��z�^8
7h��+(��1�߄<ܪ܄ȓ9&���%E�!�F�G� ������?ɡE�{�����J[<{Ƶ����L�<!sbߔw6Y���ґ}D��Yfg^�<i3�֊mx@���(R���'n�X�<!���JhI0ύ'�hݩAfZY�<ɐ�G?Qvn���#��:O���wc�Q�<)UA�l#�̣�bƙL�\���K�<�q�Ñ�#�mH�#�h�:A��A<�#TPR�@�N�pȐ��P"T���a��E;֧C�*��İt���^��Q�ȓ\5(�3oҼX[�@(j_�+k���ȓ�
\����.��ˀ���-�~��ȓ.�Zc!�]-�j�%���jU��-.�)�$"�:TvjQ�q�>
��Dx��'��p�e�̘�af��l��	9�Or1QA�ֿs��!tiϥj) ��"O���'P D�vp�`(r�9A"OU��[�R0��N�bE��n��yr�H���<�H�'4Vl��!Y��y�B܄w�ܔ3���1��]� ,��y�gZ�j�Jy���-rs1钧�'��{��_�����H;��@�֩�ykJ�Qٶ���J(2�H���ψ�y�"�b�d��"��,'�B-���ד�yb ̳z|�S�"0!J�*U���yb���$�q[pFX^Sb�
D�"�y�*�:"b�23�)P*�T�����yR���
��ȫ�k؂�F�@S�+�ybh�n��Ʉ�Z�8 
\��yrH�R̐D���|DK����x��'�Z�&̞� 3X؛�Bܳ/���k�'�t�[�o�W�
yx�@Ι,3LtC�'q���o�a��fhL;6��|��'6�LP ��G=Ȱ�7�Q�_�����'��Z�_�+^��N@�l��,��'��cDG�)~0X��̫x�*�B�'��x��) Ii:����o3�5�㓙�D�OdM��L,h����o�#I� �(�"O6��B?玘KWnS%H��Y&"O��f'A w�U��=J	$1��"O��ddH�#��M f���P��Q�D:�S�'qۂ��g�Yj"��Z�ߣvv��(����ێ@鴄�צ�!�4��(>8�ᖩ^�/=4b����
XD��d����օ�W.��y�l� ��%�ȓM�qz�+C&s(&�1C
��Ț��hZ�8'	7ib����4���Y�I5���X��V�&kf�pmi��B�5���Eb�qVfX{�@��..B�I%�X������U�4䂤�S�T�B�ɀU�%��&�4_E<M���
B�)� �lb6����&=��)��|�VU`�"O�UI�O�3�1S�g��X�j�q"Oj@+5��n�f(#A,;W���'e�'�h��fաUU��ۆÅ �ȅ��y��'��y!T?U}����a�v��-3�yR%�`U�#�I�jR���yb�Ɛ:F�墴��
3<`T$F�.��'U�{2�ea��CFB%c^�(BL��y2�ثN�@*w-�.N.E�&A	�yb)@�wՒ���DoG�2�d�7�0<���$ڼ3P��t`X�Fh|��ef�
��X��	#:���a��I��P�	��C�	n�r��̉�-�h����T48ϸC��/����`O+6 ���$_���t��`Tˏ�5!�	�kN�p���c�6D�l�AΟ���=C���ht+ֆ4D��[�'��9���1�L�a���#4D��RǬþ_�ȡ�RN�sS��邤>D�TxB�S���Q,UeX���6�!D���b-ϭ{�r��-
o�ԅ���,D��gd�9Q��`��(�1ҙ�G+?�	�c}��QFG[�U��)fڵx���ȓ.[�xR��Z�#��I;0��2\�ل�$�~�Ȏ�j���o�kM� �ȓ��e�#�D;bS����`=��@�}0c��*!v��*� J�h��ȓt��p	��̑I��l�F*S�%�x�ȓDF"��E�ŚV$b�����1o�����V�9��ū	����f�-f��e�ȓfL!��*�*lb�C�'�&x�(H��PE�� �X%iFY�7J�()���ȓ]�ء�q��>)^��n۫t�1�ȓ#�@]BWc�S��|p�X$J+�Y��P!��c�B�4�� h�B�����g��ܐF/�S38@cb�U<���.��)�?�=�!G�(g�]�ȓK� QD�"J��)���$B:���ȓR�±S��(w�Q�w��"�����z���`��/0uQ���ܗN����ȓ/w� 	@�ɮ_�x�hu r���ȓ\\) rkN�7�@�yЭ� D��a��+�4�,JV�ɰ�N1xP]���!u�߿n`�\�2��de$p�ȓ�n�# �����,��ȓ?�l�BmD�G:N��4���N��ȓH�J�sPM
>TEBSE�'�L�ȓ8�6d{�jS�B���&���-0���E����%�2WVDaG�C32̆ȓM��Q�q�Ӆ:�0Q��2K;�\��m�(�	��\*y�l;$@-s(����[
�4j�*f��c���c/���{FŚ�'`��g'ی/�̈́���P;�F�#�Y���_1��1��_�����	�kBj�z��Ϊ`Յ�j�����5)X���n�k[��ȓ?�:h
�mR�&�:�J��W)u޾$Γ�hO?5�N�D��xh��ъs
�W�<D�h����$ȵ΃� ۶�"P�-D�8 g'L=<���9��#��Q1�,D����Z�m+�)��˫� �1
*D� ˓g��~"����*J���ɥL$D���T�[VPs��05�|��S�.D��`s�N�l�����͐I�E���^�����D�5���b�Wk�( vl�S�!�� �\�d��#(.T�f;�n1Z�"O:��A$�z���#�����1�����i��+��ȁ�+r
 Y��:,!�d���${e� rD��)��Í
!�Ă;2��ӵΗ&_b~apN�!�Ç�<a�0��Mi�|�4��6v���:�S�O&�+��Pdt��tIH<0OFLi�'�TsՋY�b�*��S�C�zt�0[�'��M�#�3&N ��u[ab�y�)�S2:��jP�@(|=���"iqnB䉶PgEX���B/@�s �V8u4B�	0�2U�2�4�lř�(��M��C������S��aȎQ��A�-nx�B!D�pG✃�0u��K���0` ��?D�dIC��,aJ��5Ɩ�H�:�x�+ D��R�ϑl+V�;em�{D�@2�=�hO�� ������-R��ԦͿw��C�ɑI����E+(ČM	�Ÿ�nC�I0BĒ� � l9�U��"f� C��d�,a�Q��B�!P	ґp��C�I~��0YS�Z�
�p:���*+&�B��^-���㝉e�r�h��[YnC�	�y����5�"��e��c[�C�	?H~8�p�O��V-�I�B�WE�C��.n� %�ׇ 9�6$�$³PЬC��)QF,H����3������x�RC䉀�Х�&�� �5yӰ�hC�	�f8lD���C�v��4���Pj�6C�	�`�|� �(�6$Dp2M�,xyC�	'�.��܂E��y㵏L�XS�B�Ʌv}�Ȋ�G1�9J�h޼E6�B�	[���@��6rua2�	
DJ�B�ɲ=N�A@)P��TM�p�/}xTC�ɧ���X"/�m+\���h�C�	�F�l(�ʔW���N T��C�	�N������"iL}�'���"O��@��[��ؗ�E�e�V82B"O�A�2H�Д�2hQ�kz���"O�y���σN��]{�'��X�ۂ"Op�Tb�/M�(��Egޖ��0"OL����ШY���x3�0���4"O䬉b�'6�b��Y \X�i�"O��� �G�%��!��c�.S�D"O4�q��A�z�mA�a�S�<�y��	K�O�����&�hh�7�O!?���x�<��o�&"�Ȩ�ӆ����d�"
l�<������2�-P:��3�L�<I&�ҫ��0ذ�n��1��KN�<�2�ގ	5�<�Q�Չ\A%ӷ�M�<���	�%��hH�&�Sx��b)�t�<�qJ�9Zθ`�2���J��@��Rv�<s�H<���K�O+���lh�<A��K?�y���>xu��3���`�<qp&�}� p��'�(��-D��pr	��^XXb�B�z ��ǧ �hO���Y1�W2a�ҼW@��C�I,;�n�����(�){�$R�C�3`���`�9�x3AŶJ̐C�Q_
9��/�"l�d`�J�G8~C�	����$��{z%�Zhq�a4D��p��9܍!d@�2�����@$D����+�ISR���#S�}i�Up��"D�4;0����qvmO�U�Q�G�3D���C[�?���aSd�9?V:��2D�� ���P4A�hԒ@R�>��y��"O��S�Q��`�ϗ�r4i1"O�i� �˿b v��1��R�t1@�"O��%IH(pR�@�)�<j~�P"O�kc�E�J��@��CI\̰!"O�h���yEr8�Vg؏ g!!�"OzͰ���)��|S�/_�}e@�@�"O� !&�A ̒��F�0�'�'x�Br��*l N�j�+��"�J	�'�䢵��fp+5���^�c�'q�l�� ��k��z�n���(;�'����&�ɿ)i8p��-� �n�I�'g�d��5&R�J$�@�@�$a	�'[,e	� G-\Δ�bS��3�xIX	�'&���J�6�B�[�)�%x/�-:	��?�*OƵ��f�>4?t ƃ�ێ�p�"O�ӵۜn�0�#š��V,�f"O h��JI�N$݋¡�!M�8���"O��x󤆥�z��b	4M�A	"O���*A�X(:��� 1
��g"O��C@^e��8�"��*(B5�`"OLH���'p��d� �2�*=�S�'!�O4H�t�m
`�8Яx��M� �!�Ą�G#F� ���	B�ءRub;|�!�$A0����L91��H��j '�!�I��I��dʼg��(
�jV�Uc!��3�^9���@�0�gQ[O!�DBG�V��s'�a9��P���pK!���]Z�d��� @3Z���Mx!�dG4�l��&��a0А!�l��&�!�$Vv�:��@�
��x��#{�!��ɾ=P�pr��U%��1��+t{!��
p���S0%�-v�VU�(�wd!�D�9*2�� #�4����^51u!��0`�����3�2�z�%�:i�!��ٓ+�pU��E-��#2E�/a|B�|2A��q��Y�.\���(R��T �y�̓0>Fb���Y�MUP-�T��yRo�+n!r�%ƽt�l�b��-�y��T*.�a�Z�:�(�CU,�y���:�f�y���3J��zR ו�y2���rv�"2N�����L��yB��TAܼJS� �}��-��� ��0?�.O"�a &��^R�AP��C�1��Y1"OR��ꙣ_-���"���ꩰU"OĐ��MC�1�d�Shښt�za��"O�Ȓ�� -��*�F��u��Dє"O8������\������1��H��"O,E١n���$@�I�1��q0�"O�@�ЭW9 �@��&���rV�'l�'�D-B��Dk&��0�&_1
 �'��H �<R��P�%�5+(�Y�'����3ʈW��rE%�(s�1�'dS��N\�If��) $x��
�'��t�ǝ �r���ƹt϶�`
�'�L�J6._�^�^�BO�=}}�|3
�'�JM0�V�x���jBGB�_��	���D͂3̺m��RMB���3!�d؂,�����C�M�����)�"A!�d݄J�ȱ�P���0~HA�H³=<!�1�����$$�98��^)-)!�$ܭ��p���z�C��̙X�!�O�|^���l܅_�2t����2$�!�Č=I#أXh)9 �q"i�O6�� *!�1kښ'b�`G�JE8¨�6"O0���I��H� �o zJp� "O��)2NC��bM�, 0��[�"Of�rK	K9��,�.9�M1��'��	`y��O�H��j�l����{ �!�y��iV�\(�?
��kE��5�y�,ʧ:Kr�JJH9ze�p����ybM�""B�Є�1~���3iѝ�yN=h���ON�i�t����_�y��	�R�6��tk��Z�4 @3i��y��&X(�pF�*� =s�%S��y��_F�Ru�d�\62؅���y2K�nԊ��5.A#�7�߹
_!�$��<���7�G7(Bp��K؇\!򤗳m��I�&̅4$�aj�=\M�C��@h��0���}�h����5��B�	<C�H�z����/,�S%�IX <C�ɳJ�h20��}���R�ݒ1�*C�I�x�^ċAE�+v��&��U�LB�	�J��D��曙!5d��U�E�h�B�ɖD	�XA��cN]�ª��(U�B��\Q�1Qsj��@>��yA!ڎG��D���{�	Oe��+;��n7D�Hw����c5���'�T� 3
6D����D�B�P9@qi\��͐2o0D�|
C#@GH�����,�I E0D�D!���L�h�A�(^4��Z��.D���� �#e�6�)cn�<ޠh���'D�P�e��Q���8r.��G��	7�0��<I�V�F�}�j��$i{���]�<�p��.S���Ch�S�$1�T��@�<y���(?�$9��
` ���@C�Q�<�0�SQM��9�P�y�LH�G�N�<���ƍ��G�=�����d�r�<����*2���� �))��Tz5�Ip�<��*�l��T�ī\)��X�ǌSm̓��=��j#]����VX�$���Mf�<	^��Ts0/�8R��� �U�I:b���ɂi��H�֋�3Y"�`��@�B�	�(��]ATM^ �D��ȓ5<�B�	1}� 㐀X�m�Xʂc^�3R^C�I %YJ��T�!�����-u��B�	�͸�˜aC>�͕�~�c����	�vAْ'*1zt��ţӔH������?E�d�'rb�`Eh�'/�A����Dﴉ��'�Z|4���$cnX�D�8;\X���O�u��
�+4�Ĩ�*�+~u��B%"O������xhLI�)v�4��t"O����G��i֠,*$(�cj���"O������"`r��Ǩ��V^&�k�"O4�(VE�`"�Lʥ���f�騀��TE{����i�.`���\>��a׫�$S��2��hO\���E� jB���Z�V��T;C"O�9��ND�&$���i��m��{""O�h2���W`s�\�9q,<*U"O�1��ȑ�bk���� �A���0w"Oڌ��H^�2�"Ȥ�؏~�1G"OX��㒁d$����I �:O��%A�
�C�Qt�TT�&/�!2���%���IM��:.�h�e�Ŏ%%P���W3reC�ɔj8��s��˖K(�hG�T�9x�B�	�c9�Y���^���L{Q�ǖǢC�I%p)�0���ʑk��A����Pg�C�ɬa7<�
��]B�U��"�=�!�� �Q(�d��U?���Xg��D��"O|�ؔ@E��� ���S��&�Xr�'��'�t�:&LmS,�*v%� p����'،���¾ @1�¡�d�pɛ�'`���ǀ��3�лr͜	d��'c 8B�/��V�ⱂ���P�[�'d��1*z�ʊ>,����'��p�A-L[	@pC�2�Υ�'l	� Q(:H�GÃ?o��Q���%�'03�=Ss��}� ҧåVPF`*O��O?�	�U
b0@��8q�2�� `�0B䉾n��\z$��Rݨ%
�yI�B��u�#tA��
�z}+F�޸NM�B�I�	
��5�P�4J�0��I��B�	�"+l�@��_�.�#h��?�B�I/�t�QǍP{IB!��	�B��䓎hO�D�7�N�0�(^���
S4]�!�DJ�}ʵ򱢝qג〉�<,�!�޼ba ���J���iQ3Ԁo$!�$�����Q-��!��{���2!�ĝ�}�z=��C�?H�ޘ#V�l�!�֛:6&Yq�fS�@�BŘb��2D1O��=�|j5烩d����(ΞE�P;'�[O���=y�'_���\gK�7O��0<���DU/�4X`V,��HE �p2k;}�!�d%oJ|Kr�N>��P
�?U!�Ѥ]v��b�!G� �U�D�A�!�d'$��:G*L�������ے�!����,�c�0{c@�q�Æ
5!��I%�u�#V5NQę ��/	a~�S�|@��X9<�C���>kS�����>D���]�P���)$2ٲT{��9D���A�̳b|��S&���l�jt�+D�pss`@2�FZC�z����o�o�����䉉�>���D+JҝA'��]@a~�V���1 �<���%�ma���do$D��Ȕ�Y�w�ba��œ �ƽ�c #D�l�E�/�T���6`�1��6����8z�����ـmv�y�#$�soNC�	��|���LL(�]����1�B䉪c�0�'L�7�z���1\����hO>�r��Y͐��Ǘ�hlR4�EF&D�|��ʜ"h�1�c�@,'�ԒW�)D�|�1�[�o�aS�l�t��貵�,D�H	1cP�M=��c��LH���My��'��D �	��Lx�k�""��'��u�R%��4��;�n�	..�[�'u�y�ܽc8�,ʡ�@�"��D��'����T~��x�! $Jf����9� ��D(�	���eP�����-:˘A��"<D�� "e�#y�p���B/o2����;�d���5O4�3WL��.� &�ԅrTx���>	U{�̤�f-w?
�JG��j�<Y�-�$��D��t��T�U��i�<��ह��������V-�I�<vm�1w��$C%��.��@�}~��)�')4<��q��D刧��hk2��<���ap�,4j�BE\=SD�ȅ�X�II�F��bj�K�e"ǴO=�B䉴%�x��	*3�@p	�톀ZbB�I[�69@1c+\�:��L%F�vB�Ɍ²TS��E�b4d�ޒ.�VB䉣E>�ؓ3�J�Xd�@ڹs�@�q������s�끝X���KA�
ΈI�++���<E���� �T¤i��L�$kw�	%$�Jt� "Ovͪ��6DD���9A����"O�	�t(�O���V ��T[j��"O��$V$U�2�AB�2I�2�"Oj�ё8�x���;6v	G"O�i3I�y��B�n	:h'^��Ā<�S��yR�N
If~8b���3hJ���$	�0=	����/ h�挍�X��p��}��'C�e�'�2���w����
C�?�� �S��y�C� �	2-��9G0�3P�.�y"�2V�&,q�Q�[��dH����y��VF��!뙴^H8��F�	3�y�(�*L�p��u(Z/mg$Ɋ6���y�e_q8)Za )g����ֆW�y��C�U�D���m�]��\��fҍ�Oz��DU��^�B�ً8d���2�!�DO�Y��U�=���技�'4!�Y�4���a�/�j.�$�EDP5(!��ֹ�B��mM~�\����Q d!���*]�V����_.}���ɱi^�!�EOa^����S-c�.]�B\>X�!�" 
����&RI���s�v�!�$ʚ/��� �40.p�oՉB�!� 7"�������C��:N�7iZ!�8L5��Q�AO}� 9Wl�5}�!���	Ipr=x*�$I�4�[/!�ŻF�XhӇJϕk��y�`�s�!�,��͛|WV��A��%Y!�D^G�]ˆ`�q>���.J.<S!�$J7Z��m�t�K�IBX�k�+�D!򄉪m�z1p �\�),�+љ !��枈CBa�8 ���ēoy!�$�� <���
�.D��,��s!�J$1�\����(PQ�7r!�SJf8��܀p��C� �!�d��!i����͜<x�𑓢�Z�K!�$G)Vڐ��s�V���r+\r�!�dI<%;����B�$r�����T��!�d�2J.U�$H@�ffl3���M�!�d��8�&x����/tN ) p.Ðj�a|2�|r�� +�Fљ�m�:#��T�v�T�y�-U*��TJ�%#	N11���0>	���ф8҆H�ק��q����B�ƕJ:�=E��' �Q��*L�\>�����#���"	�'n"�� �\�7,ư��CX*G�
�'�b�j�ǝ�@�&�
�h0v��	�'^����A3�h-�t��!n~D`	�'7��CF�?z)��
�aG�f��tH	�'��"�cΎ%
� ��׾4 �	���h�(��W��zm�!��#7�!�$��S-��
UΨI���YH!�(A���s���L|�*�Z;&!�� 5h��!�%ddE�%:.z�!���(SU��a �2]�04��pp!�D �o�e:,@
fJN$��7qX!�D�`Ӛ���ʅ�A5Tq�0�K<P�!���OFX3@Ą.o]e�Q�;N+h���5��Nx�$;b+�+pR@�`a)�(|2`�%D�`�Í*�6� w���,r"�0D��y�ĳS�f-C6��=��@�ģ-D�d�q�G�Oj����@�j�lp��,D��qc��N�v����o�n��q()D���OW#;π�Rw�<yd���(%D�Dѷ���-���P_� �k�A6D�� �|¦)��'@fYy���+���Z�"On�B�ݨE �а&ŏ�Te���"O(��6
�6��5��xP�!B�"O~p�VgU=M{�՚A-�B!	�"O�83uf��$�4t)�o(�-s�"OH�;!�C�I��q�ɉ�}�|t��"O�A�,JP|�j��l�i2"Oʍ�r 3}��2�\?m���06"ODxrpL�:p)����OX;��L*�"O�Ѐ̆;"�^�T/��$�er�"OZ�eoW�J o5<��"O�ݣ��7�$Q��N��,Ш��"Oh�i�Z�(�KE���_�h�`U"OƝ����A�p�� c�-z��93�"O
m�tE[�%�vD�TO���j,��"O�%kЎ�5'�N�07oֲT��"O	��B�`Ii�$� ?�	��"O�Hj�h�����x�B���z���"O(�P��*o<����PoPd"O�i#�D�i=�6��>9ի�"O�����O�~��`)v�Y�^�\�V"O�(�G3#��q��G c�ii�"O���)�<A���ćM&'�,m �"O��pl�r��qK�%���@P�"O���lR��V)�G$��.s�X�"O��)b�l" ԩs%P!)W(ՉP"O�t��>%F��R%܎��4R�"O���I�xdb'T��p1v"O��0���.�f�hT��8�h�"ODi ��3m����ǰG���"O�8�CD�v���c6�ؘ8Ժtڲ"OF5�$��)��A�oP�/��X��"O����I )	���퓼Z�x�@"O��'�M;���!����%_�A�P"O�q䨍�_�|�(#�d@L���"OV��B^B!R�xS,��NzR"O��k�ʒ�H �U��<Zm�� �"Ob��F������&�k�!Ӆ"Ox�#�ϋ�N���#��S�@�|�RE"O��!#�3j�+ץ]�c�|x�t"Ob��/	�0ƌ��7�S�&-c0*O�P'��($�#&�9N4���'�,T�S���Dp�FF�rb�
�'v��ph�R)VI�զ�m��M��'�1���#6���ի:T�,��'0^]��
�nbX4��BK�t �'yb�5(Ib6��t�Al�'a|0&�� ']>�Q��?��@�'�|�:���A�0Q'���I�N�B�'\|.��=z��@]̒pce��y���1�r��`b��@���d��)�y£��=%�L�'�ζ2�pّ��Ǆ�y2$�5l�0�2�OWq|d��R��y�mә!�<�۶�]�K�R���!G��y��/8�A8�KOGx�4⇠S�yBC�z�4Ц�R�=����b��y��4g��ܲD�ު8&��Ä�Ǝ�y��z�L��`! �6P���Ѧ�yb,'�|R�k�A�|���V��ybl�gǆ�J�j���nX���˱�y�+ƾHʜ;&�U-���S����y"&F�熸�W�
�j�90�L���y��P�+��|����5N, ��
]7�yr�;~�j��4"R�0&}y����y
� �:q�O�h�%��׾|�z�c�"O�D���
:�Hs �I�B��"O��C�ã+OD��v��k��p#�"OT��S���7�VБr�:[���Z�"O$�+���}|p���۹1���S"Oj�n��h�Ћ �)�"�*"O�u)�L�?/n��!A��|��0{�"OҀ�dY���UA��\�)��K�<��MX@����!�́Ɔ[D�<�a��5��N�D�i1/PG�<A��I :5� �a+�J��B��B�<��)P#(P���)�;<|F< �b�z�<i�	��:��y5Hմ#&8зH�y�<ɱgч!P����O�w=�K7\p�<�,�0@�K bͶT }+1��a�<�f�Q�B��e�/���C�_�<)� 0j����]��Rԛ���t�<����u�ƥu��B焐C�hSp�<�r�@3�hɃGH�<(S���d�g�<YÇ �$�ґ�Fȟ'�`�����a�<��az�� ���^�:��T�<�R�Uu�t}h!��1"�B�� O{�<)QjKr=,xh�������Dz�<�QF�R�8�a]w���ը�v�<q���{O�|2�-X�P�4%FW�<I�&�]Ɯ�D!өav:�j��V�<I2,�!Z25���>�vl��(�J�<ɖ�ͳ��ɺ&�����qY�<�
�n��]!#�[郎	vo�b�<!�n�>8�r0��X
����Q�Z�<���p��0ء��|Z� ����U�<)��� �B��FC� �~)�V�R�<��K�5[O�5��iR�kr�͠s��M�<�D��)��Iɇ�2nVYh���N�<�������U�V��/`2��g�_M�<!2N�}�ܡ���GL:�
��P�<�+�<�.8�ЌC!j�� EgEt�<Q�� �?�6Qs�fM�	�c@�K�<Q��]yAQ �!BP��E�<��O}xqx���B��Y� ,~�<��FW>v�4��V,�T�nQ*�
|�<�����nO��0GC�6�����#Is�<)�iP�hM��x�4"L<@BWn�<q�Y	���á�&B�R�`eO^i�<��C��LX0�C��r�%��a�<�S� =^��! '3pGt(D�S�<Y`杠 w6�� �;V�*u1 �j�<��aψ^�@M���̴Uܔju�k�<�p���/f���\�1z����P�<�Ӎ�[lQ�D�<1�� �O�<I@Ň �����%�a�'\H�<I��Ս �ɡ��9P�T��A�<Q�B©2�$�ڷ�,�j�I�@{�<a��9_��p�D,I��U�!�x�<� kʾL���r!F����iV'�|�<a�Aƒ<?�i�E�p~�@���N|�<�ph���T�����MU�4��O|�<!�@Bq���AnƀX�-�6��w�<�vN�m��u���M?u�Ep�/�s�<9B�
+��q�!�I�%H��p�X�<�4'Բ+� �c*�'��<�F��^�<��ԕ	���3W#^)�e�v�F�<�W�˙�|8����a�c�UD�<iP�/2��9r��� !d���K�<� ���h[,b��va[���4"O���ᇖH� �hB �?u�f�"O��JbNԶg����ԎN�mn�"Op�*F���!����m��񢤚�"O��"�]���pB�S�H8��"O��#qJ�^��5� aВ�l���"O@�!
^� �``
7oҘ��� C"O+ nܽc\�H�B���3"OH�a�I� d��m��&���"O�t� `'n�nY@+��hn"P��"O<�H��� z��t'��<a��D"O�a�f��'d�#7�/9T��"O�R�t��� rK� NDQJ�"O  �BE��{���>J���1"O�(�[|fm�B,<.H|�B"OB�z-A�}�reԏ$\�9+�"O�=�@�/):(uۗ�ɅFA�	�F"Op��R��"1�ڡA@�/΁Y�"OP0��A�H����@�܆>!4�Ɂ"Op@�p��	Y��7O@7<��u"O�����ϭm��Xr��4�d��"O�]����(<�C�C� l�|��"O-)�KD;L����#Λ5����"O�tCŬ5�Xhq�6���"O�#U%F�r�Ip�'�8�2�s�"O0�$�
P0`∏����	�"O�i�E�<0�^ɵgB�\٘,y1"O,����-�^�8�N�B��!�"O��s����}҅�-_�<�۷"O�����_�-̚�#���V�l���"O��#�Bct���&�}\b�+"O�%ZB	|H���D��@s&"OXɐ��֯.-�1aj�8�5"OX�R1�.y"T�2�MR����"OxI���ݟrr�!C���X��́e"O�`�#]�f��zӃQ�C9F��6"O68ADٞ>�ܒt��
�l��f"On�	GiR��&w�Pc"O���������tۑ��I<P�ȓ;��d��Ov��Uӎ��cb�ȓ	@⽱���9J�V�jʁ'"a�ȓe�Jꂡ�%k��T2"O
�B^��ȓ-�T�h�!���A�b�6U�Ї�B���t+X�:lT���ӵ{QH���1R t�3l�Gܰ�𪁮2l�=��Uq,)��M�}�jJa�J'�� ��UK���2#�C�`��� t���NX�V��Bp���'Q	V��ȓUD(سp�'�e�6|bf}�ȓt�X�4lA3m� ��HF����ȓh��4�T��=��4�P	[�~r���ȓT���&�n3"��֣*�)�ȓ25��Q�������B�N��RŅ�$E�� G	H�4���1N˗J�T��F>yڇ,F�*ϸq�0��':���CV$:!�UB�褫4�֥ �i��S�lq �%C8(d�
ş2�8��ȓ����K��Xw�?`��]2�k5D� 8C�Q�u����o�F1���/D��`6�0WF�=��R;.:w"+D�d�eFʝ
ʄ����*H(����d'D��K鉙r0h�+�7����#D�,�'H�m`�Iդ� ��I�cn7D�d��'I��mܛ'i"Q���4D�� \K`L�'�BqaBM�
�r�rt"O~����+�Rq�P?p[>�X7"O��娎��"��J�nq�	��"ON$b�@\���fj��BU( �Q"O@�������͐`��	 =���"O8��3_&s�:1�P�C�;*v���"O��"�n�?F�`�;`ϕTl���"O��7���=r�ER��
g�Tt��"O����ؤ!�BP�SOύ��;�"O�E��o�g����OӇ���B3"O�Sūד-��a��̒���u"OP�rC��?R�x)!���*$4$@"O���A!��|���#! ��n�-ڣ"O�P��C�t�b�ˀY�m�b�*�"O�a�쀌�b��2e�?)X%"O��1bٿi�b�C���w3��a$"O�'��Q{��!�e!���"O���֩ûrJ�IQ�(��S�"O\���n\�1�D�h����B�@@(�"O��95��(6�X(��8G��"O���@��ܮl �k�6e:0V"O���i�#2�
� �K�~7f�P�"O@01S�ҝA���ڕ/�,fͲS�,�S�����m,C��9G%x�\C�	)7㠨F'	�z0L2 �:	d�<�	˓mc�a��"6L�-�6'�6`����3����kT3($A����,��P�ȓ
oڰ8�G�/T��!�`۬I�|�ȓs�҅�M�J��đ@�
�H���#�������cnl�P�j��m�<�U�/�S�'nQ  ��ןd��0��O�KJR@�ȓ\���G�;he�E�"pEy��'0
ec��ښx�P���H�*��x
�'�&��`�d���`M8*'P�Z	�'m<��D;����G^�8�T���'>���aKɛx�&4�u��/��D�'�N����<
��a5�P.v��:�'�@�'N�+x�� P�ÉiiH���'���hVeC/�(
Q��"��Q�'ڴ���(8h����l�8	�'�0���� 
��:dǍy�T����D)<O�)rvG��Zv�6ȁ˂k�,n!�$��}kE�6C_����6e!��?J�U��C�2�j��C��SY!򄃦z�`�HDV�n�6��D�*E!���B�@�/�2U�n|�0.ȑ 
!�D�	Q�0�2��B�������,.�!�DD�~����N���O_2�!�dǃ[�T���KL�I��8�S���t&!�$�<&��ks܋%C�u�u.܇M�!�dB7r�Q�d��+Y^T� �O�Eh!�DI����@�+ة<h�)�W�֚QQ!�dZ8sy�(�*3]Mµg��X6!��T��PXi �Ae���U@$��ȓ���T+W�NǂD� �[k}�q��|��Yh! ��F&&}3��ڱx�X��VN� �Ն 5<��h���{�"u��'d�Pg@E/~r�� ��17�M	�'D���'�-C�b�0�"��}% 5��'��]Ӧ��;f�0�ҏ5o�d���'G�Ļ�C�{0�)iG!�
�4y�'~ၠd*@����V����6u��'��<s��R�:V�t
��1y�z���'h�UI��߆D����%D�(9��� � �T��r'��9��[G#h<y�"O�� Pi�u�##L+�}c"O.<�E��#0@����!	(����"O����(͠K��QIB��93����"O���w��m᠅��6��`J�*O��� �K�6 ��MP5]�ڔ��'�m�0oP2��y����X�0�
�'@v��P%�M�Õ�P@!�
�'
�H���[�D�R|���:w�|�;	�'0�q���B�2X���#�v�h��'����t�(=6�B�����`1�
�'04��BO
�t�#D.J�o�.e�'�(�@uc�:l0�����6m�΄1�'�T���Y9 �p#c���n��p�
�'>j%�
ĝS�ܓ��F�c��
�'hĄ�1��(@k�=;��_�^�x�'�j}�S��n�=��Z���'�r�����_<0B0��{��(�'c�4��݃[j��B�R�b�d8��'�pt����7N���6!�Z�r�H�'`�85�zl��f�Y�B�[
�'�^�u�͠-q�p�YC�D��	�'%(���C�<c�~�{R���L����'(6�
A�[������0�X��'[�Ғ��S�\��gX&j���'�"��	C��Q`#Ƅj��#�'�bL�lЌ~�����%ex����'�
A�����,�C�NX�8 	�'��<���X2w��Yӳ�R�V�"Dz�'��	�+�}n>A3Vl�GpL4h�'�.�ig�A�V ���U-��<.����'è�QG_�8_���f :ˬ�
�'Ԝ=i��X,%b虊���wa�M�'Ȏ��a.�?� ��V�l�r��'ؒ�ȅ��v��AJC'�#i,>i0�'ª�1�`H�Un<P�[�N��'�4qȶ�{�@3v+�C�\�
�'������\Xc5l�:
�'�l�hq��Mqp\�e&[3��iY	�'�N�cW�ٺ6���;U�V�-r�ġ	�'�Ld2 '׊QS�)�QcW�=DD$��'J8x�1��o�yPJ����HG�<�A�_�c�,�e��`����7 �Y�<���I�C@)yU'	�h8�SA�M�<�����`�	 %%��!P�hEF�<ar�_�1�r$��nB*AG"�9�F�<����.����MD��q��[i�<��BA�8IP��V͘���0��h�a�<Id��v��At�L���8��]�<�2� D@ϖ5n�T0��H�U�<�U+�u̞0�FĖ쮀����h�<it
,l���0o�r�n�b�/AZ�<i�g_3�J�2 ��7ᖀZ"J�X�<�G(A�l����-Y>dRz��+�{�<�ˌ!&La�g�:=�`:0(�K�<�� �C�D�t,K�6Ț�)u��G�<Q��C2;��qI@�0�j@��J�<!�E��3�-��:�jVD�<�a�׈Y�� �@�����I�ah�<��F�lY��A�l�{���e�<�7���@X��FO�$�Zei�{�<�mp&MbF��Ym�m����L�<��m�9Ԭӧl��V�f!�&A�~�<�B�P��t�dK���@$�e�<� l����J�4z`к�\+�����"O��ԭ���	��	)���p�"OV�	�c�'F �W��h�h�"O�=q���?��`�y�F���"O�Q$��:,lHė�;�����"O�|X����a"!�aT++��-�g"OX�bDʄ87݀�(�"Y
�Ԁ"Oty�o�P��Dܙ�p�R"O��P�	Ү�C� ��N�~MX�"O�TP: _�J�ZM�K�bv!��On�2|3�$�o�X�����bh!�$B�0@B�%��~��!�6ğ�kV!��ϗ/���C�#�C�Dq01`4!�DK�{�TA���E��J���AY�"!��u�$daˈ;Ĉy�qjԻV!�d\�t��3�o��?Ӗѹt(Է�!�Dϱ]P~mڥ��*����#��
'!��&[R�z�J؆`!DU�!K�1!�,C�t]q��^
B�w�O�H�!�I�h��M�꒯5�l�q�ճ�!�$�:y��d�X�wʮ�Y�`û|�!���)�����!:� =PD/ӯo�!�d�� ⒜*!�@���I�	�M!��.�Z4���͓Dd�܂p���'�!�d�&L3�E�
���>	2��΂g�!��W����a�	�9��d�c��I�!򤊧pE
Ic�iñe��%�w��6�!�R�Xmf�hQ�@�'I���#Ȯ2U!��AD�q�k�W(p����A!��9�F\)��hK���!�"P'!�dH-8P4���fi`���7!��YR5�v�T�;Sʰ�S�^�!�d
�E������0s>�y�/
�!򄇟O���� �Lɮ��Q�]e�!��$i�lM�!B����m+�l�I�!�䄦�� $+�5c��ݠtb�8ag!�dπK�(��k�H,Fd����~]!�F�E'rep㉩;�8���`��\!����\�1T慴�4� ⯞�I�!�$I@�|��0��W���"R��,!��*���q��ݠt����ia!�Dؙ<cD!QQ�ֵWf��MV�jL!�$C�"��)BTe�(4PqyC5M-!�D�o^����
4f4 P8aAҎsvў��;�ʈ�EA"4[Z������C�I�J�����5��ٙ�'�)2���+�I�p|�H˖E��}�s�G�fKB�	�x��xI�Q$Va��#�҈��b�E{J|2����'��`���_�L�&DO�<���]�A�y��+�d��Y���L�<9Q(� y�zQ��2��	q�^�<q�ŦQ.�]K`�>/�]q@"OW�<��#rD]C#�%)5jx���V�<���]������'%ͺ1�Ii�<!� Y����˗�؟P�����@���<%>y��ۓ-J�P�f�L�۲�9�-#D��a!�v~|
C��n2�إ�9ړ�0<�QG�0=}X� #�t$�䀥�U~�'�?a��[�N\�$�gU�LKo<D�����{	nq�F풿 H�D��$��@��ڸ'��aҴk�.XfI3G��>!l�q	�'.Α8Wb
�u��WK�|J�'*f(�P`��#?���!L�'\�,����)�d)�f�������N�	RbS��y
� �)��P"#`���%��)6#����x��)�S�Bm,�І�<�0�t�܃S7�B�	/Q�伺�+�;Oq�a"n_3]� B�IEsvp:��^��>9J�B�X�C�ɟR�ޭɅ�ʥc70� �g^�,<B�ɗX%�|9`�@YJuY���*CJB�I4q`:�
�҇7.�Ȕ�5l�TC�	<r���FF�� A�88�<���y��)�&�A̽�f�	�V�L�vF3D�`B�Gf���UE���5D��b�
�&��-�3��<��*5D�|k�cǙv��9b�8E>�!�M2}b�)�> ��4�����Sx�r��t�N�;����Oְ�6�˻R||��V���Fl�%���$7lO�� Ao�5�r4�JڈoUB�q6�O���I�/	~�yJ�	_*�!�&�,!��mt\���j�?��蛳Gۀe!�Ą;4�"9�4ț.���$�*	 !�ą�-�⩣b�ˍo�h��iB'�!�O���a)Di��&(��o�!�䂿a썢�`F�]am��W�&�!��p�Fh�(O3$��ʆ��>,@!�d��yo~S�LM��ԁ��	&�U�ȓ�`���̉M��1���hq�ȓz��PЪ4��(��m�%vɇ�\��l�lپo��hb	H(�(�� �h:���[,�[�� $�Y��kI���`mܐQ�9K��ۤlR���Pֺ8�̅!D|b!�gE�L@��Ɠ_*t�.V�6���j�͟9$6�J
�'~I���=�H�g�!'�
�'}4��F$Wl"@C��!��l�	�'�:q��I�p�r��Q �4=�l�1�}Ӓ7�1���<E��N��p��|+�aKC�� j�Q�<��_�ȱ�P�P1$��f-�S�<�C%X�"�ry&X�O�����Lċ!�$�2���#���<iJ��	�wu(����'k�����ָ.q|�+rڜ;�`��'��E(�*vֺY񁆏64���C�}"�*�
��ѱ��� i�Fԋ�<dPB�I�6����EфK.2�A*!�"b�F{��d��7z�뇁C$R�I�SH�~��'��L�q+�(ò	��N�6.�p��M����i>�&�@�c�X����{�bӫ&Ѐ��E7D��	O�wc�Q��ăh�t�0�I}��3��=K^��U��g���a"��0| ��00T^��耿s��P���AܓE���D^�O8�SulݧM�n�R�	2#�B�>IO���'%�$$LM�n�;6Ks	x%���xR��:�c�m��UJb��f��$�yri�,W��Ь~xv�1�Q!�y"
�f�t�1eB� t+� ��i���y�����>���`�p�� ����y�AϚ}�:��a��:�F�B�Eڑ�y�B��ly�i�"^�h�H�ْ��y2Ƌ�t��e`$�Sh��Tqeh�y�^V����#
�̕f	�y��E Zve���w�8�b����p<���D.~�@ ؄	Љ�����Ư����Ps.|�`�ťq�L��S	R�q6�d��&f]['�Z*	+F�BH�+B�,qD|b��rw��S�"��
��I��C�I
zX�|Y�O9K&��7��0�C�I7ph@��P�Z�5�e��2��C�)� NYPc�Rf��t��A�f8�S"O��0b(:G�\	d�Y�
|��kq"OXsĥ�;w�a�f$�[y"= �"O �`ņ!����%�� 4���"OH��G^(NA�� U�.y�$�'ֲ��I����'K9b�ZH�F�&���A-8Q�#�Ϥx�h�b#�*)BJ����k?Q���Iv*�w�H�^ܼ�ғ��l�<�f+�3&԰�$�,k8�S��_�'DQ?��6e�'w	\�2���4� z��)D���gHJ@~Tv��4��$£f'D���1ɞ(��i2*P�+c��r�O&����>�C���O(��+�3�$���"D����*�:bƂ�x�AV/��� "D�d�'�Q�uȢ}-���P��}���p?	b� [� Z#�MK�|a���Pa�<�e+B����q��O%T��䲆��[�<ҡ�$?'���G���$;j�R��~�<A�i�* bT1tǝf���j�Je�'��'�>��4kH�uHP%a���\t��`+,D�[LKe���C6�Sh�j|�Fd����z~B�xJ?牮wХ��)
%W
I�#.�%V�>���Or�>��}2�\� ��R�ܣD��{�aX�hO6��dL/�����A-I|4����6
�!�䐈nXy��V3c�����B�?����>�n
�8�F�ڥ��%i��hr�+D�H��([�Y�Jջ�`�nҠ���*�P��$pN�>�ࡘ׀��v�X%�E6�	U��ϓ7��7��X�|�3�VK�Z}��l�"��QR��H6��Q"0���'�ў��.��)�x���=_�Np��e/D�8q�,Ah�{� d�>����?D����ަE�"�Cdk(�!��!D��Zu�8im<�H�lRE��	K5!2D����`�<\&2MȒ,P�gr��b�.u����I,Hp�����31��ؒ�Q->C���M*B@�U�I��ɒ��C�I��r]�g�\��*y�Tf^�#FC�	%z;x����� � fn8~<���>�E�E4k�rQ�֎�48�@��G�
I����p6O���$�Y�Q\*����3�b�I'"O`Z�#R���+�%�8��]r"O&��4�T��P;e�\6i��0"O�L!�݋T�%
�!�"M�=�f"O�ܘc��H|:�!��	�I �"OX`��!�qMr��&� DuZaX�"O�$�����ydc^#	�qx�"OF���)[zN����#�ƠR�"O��q��H19�t�A�G�w�Vy'"Or�J��(�@���JӾx�Tв�"Ol�a㭆0n�L��d��])Hy�d"OBpx`o@��\��Ӆ�:t ZI�p"O�qeJߛ=�(�C�#B;Y��ӓ"O8�H��ԡ2N�1�-�����"O0}6%�C�lq%��	�!��"O����ᐭbW&H�k�r�乲"O,� �X�BDU3��E�ӠP��"O����75�\	�@�
�p�d"O4�Y4���+�V�B�mZnHXX��"OФ;�����88��+P+���"O��5��<�tMba,��`��"OlZR甉^Rp��*o�pAb�"O�����7ה����Y
u�2��"O�������\�~��v�?c�Z���"O� p1@��P�P�.YB�X�p!R6"O�鸡c��QTqI ���v� ,Å"O�h�ANM�(�*F�O�F�^�"O�E����h��  C��|a\!�"O0�����]����B��c��;�"O��JF�W�q����@�����	S"O\X �Hx�)�!S|m�"O�}ӷ�)'"v8��;,�AB6"O���Ӛ_�F�`�L	()��\��"O�Td\�}����� QК%%"O���-א>��r�KY�.�pa��"O�t#��;4��B�
0�N��"O�D2֣F�~��]�'(��0"OH%�u�����e�J�y�H=�6"O�:�E�6'<���,99p؋�"OحQRQ�b4�� ��-)�a0Ff�"�P�#�
/n��DԞv��)2� �|Jy	a#Ծ@n!�	(�z��4�z�Ic��Q!����0-Ќ6�ڌ���B�
M!�H _�|E�ס�AĆE��a>>5!���
�ܒ�*�P�*��fA�Q!��.�V���
��pʡ,�!��X�����C'��$��Ab�K<+3!�W!,��\��*������D6�!�� b��,bQ&�?N��h�$�2z!�@� h���8s�x<s�M�*Oh!�P�*���"��=Ǽ�r���m�!�dZ�
���K*�d�b�lV�!򄃞3���b��N�zFơ��E�8�!򤝔r� "�B�Q0�ň�C�!���O(�`'d�(R?�q�A�FZ!�dŞb�2�Z %0R;*e*��]�X!��
Ҋ��F�7.2�I%�[!�!hiBҁM,_����GR�/4!�䕤{Ur!"k��{��y�ǅ �!�D�e6�KP�8s���F�>�!�D�8-,�"�Jie����%)�!�ʿi�J`P���5ZJ�З���p�!�d�;k=���W66zL���]M�!�F!Z.U!q�O�8k��3��S�l�!���/_dMcu��(!H2��'(�6E<!���)Mi
U)W�Q0��@��B�!�Q�d�d\�g���p9x�c@܆�!�DC�3��ٓ3�3!�P�"���w�!�d@�TR�(fB��� c4�� c!��&!;�*aK�I���s��O��!��&�&q �Хv|ғ��q�!�Gv���{��_'nR���K�'�!�	u�,�e�,�X|P�i�$3!򤈟��M2�O�I�8��Ǖ�:!�Q9����e��>�ޔs�Y�!�DB$FqBQX��L)�nɘ�ʏ!{�!�DQ�xA�E�d\�K�T��U�̒:�!��:2��eqѣGQ���!B�)H�!�$�3P"F|��RC�^�����!��&MBP�����G� �3��V�!��էU������2�@H���%�!��\�ؓ�M�^@�m����S�!�$O&b���B����n!�)�^U�F��'ҠM�!�Q."i!�gL�0���2m�	ʮ+H!���0�!��쌽s�|("��Q;!����$���p%�=7��;V$�35!�Ĕ�+�.����H.�\�&�E�*!�� �<��Ń�`j��:���4/XP��"O� ��"�� �F�U&h:c"Or�Z��U�#�� ��
���@"O���g]%`�pɐ���DLS�"O�|
uIN�Kྵ��뛺(��H2�"Op���>{6����0�&��"O���0X�
����8Qr���"O��D��3f�뤁ͬ1n�yp`"O�|:l�?K̈ ���o#.-�"Ov�Ҁ�)uo�4`��I!��j�"O"�b�*'N+ ��l_�>L� !"O�бWㅧ@��`J�*K�Q�"O�h0�锵L�v�hAJXn~� �O`�^��I�d$�5� 'J�>���ӂ=�'ð}/X9�w�ƹEKJ���w��0��3`��P"�	��^)��uJ���mS�Z���Q�&E�P��bJ�*��N�W��P`�W���p��{�}�����pRE���]�؆�<���'ل���8 ��4��ܔ�Z<�&(��!�a"�)pFA�򫝵a�~�a��W��l+��Ҕ+��]���!�Aש�6=r�{MʧN�<#>�b�i�2e��ǀ�q��O������)E�� �	�0'�8��'_�<
6H�?S܀+����X��`����`M9 �����5�蟂yRƢ	�U^����	o��єA+�	n�����'��	cpkФ9���w.M4E�����X��?�kN�|��X�!������>c�4BS��7��e����D����"6����dU�Bw	yD�׹i2��[#�Ɯ]��xS�&��v��Ц��97vh���'�H���6�ȭ�3�N/ft��h#�O�xl��/_�6���M�b������5�B"=�$b�.M����uf	3R�H�eB}>���	@�7k4#�"cJ�0�E��U"
�Q�FS� �b�X �Lxu 4n0G��U6n�ѱٽ=�9BnF:,/Pac�A֚���`C�p�h���B�����G�g�,��(�~��	MҪ�r/H�"">4�ҋ[f���TM��"�DR�"+��51V,�~�7*���#�4A���l�&����:A֙�`B�4)r�ضI��*L��kd@�?�mZ�o�4 �B��@Б��"H�{x���㇂Y�l	��5D��%K�'��k0j �u`JV�'��M����8a%���ÃBC�`��J���p�䋗�95:�p��1_���A�+�dɊ6GǄ�J�B&kP< -��	׭hv`|؁J,˚�˔�Z!DO2��!lB��(O$�k֪)����t(�#AG<��Lbݩ:2GJ>M�hk�n�$̶��B�P64DիtA�6�H|Ba,�(-�y��U�O�|C���0�Vc����Th^��jBztX�	Ӻ�i0�LO�°�ߜyĴR��$�J��dު���w��8Ã�+p���%7�=����50��a�h]�\IS��2���U���'D��
Y�c�<�f�ν3��x���L��lZ�¬؉7F��)��a�0�PƅO�7��`�D�9L��T�ȗ}ը��[!J �BL���T	q�ЌX��x�d[�����Z3sj�Ye.E0@�������uղs�A�W�Tk@d[=�Pk-[0t�t���V�O6��E�v�݆h��p���jOv16�.}^�GzҊ_��]�q��7#3� ��g��<��H�k��|������!z覹�V�׵{R �G�K�}�2��n;o�tA�W�A|�����O��K�<(��Ct��QKLV���՚e闦Y��ΐ7h�ժ��ڽ^� ����E�V`Y-\!���'Y:lx7�2V�2����!t�F��b��� �1[H	\^,R+D��~��Y�A����䔼.�j��@ۑvA���Gi~�7ʞ�V�LP�I9'���B�&G�u��,^L[��x��i��R�_�xS�T����DA�
;�O�LY���/*@����3_�$YAG<4�DQ�p�V�}D)��|�s�U�U�I�4K\L�я6TS��	P\��)g���l�г��"�j#>1��?�D�3`A{T�R�������><�C��@�R�h��*_u˓�p`R�F)�x�?٦�߀f��X�A�E�|�T���g}b���s.��s�J�ΟhC���2Yp��0�R>����B0J��Y#J9�":q`e�6�'�xh��H�8N�B�B5(��Cl���'c�a�G*+@�(r��O��z��%|�d7"?��	���#��3=4~��Γ�P��&!2� ��i�X�"h�M�^��'��\s�b�CLɧ�Ԃ@Izl�'���j���3jԃ�����'� �0
A56��5�"�Z�A��Q�O>�oC��Y�Ó@�b�9����G�,��eeN�X`D}��@�f��o"J�J@*��a�0M�Ro��/�TB�I�F��Y0N�j	�`ybh� �B��vc���J�!q���8;�B�ɵe���U)S
 ���Љ�?L3DB�I�PZXX��H^+Z�@F�r�<B�)� ���G�0XT��A�8]s�up�P�<Ђj\S���ɣ������4x�(]*�nO�X������?�<t���3���(�@�0��)7gÎ0!�`��'�j�@��8��".ҩ����X�[@� �a7r"�?�z��X�g*p�j2+T�D� 4!Ũ,D�DIb�(Q�P�W��U�4EC�`ה&0p��-h<���<E��'v��t*�w(J(�GF�W���y�'2�yJ�E�<;�ja�`�\�E*j��'X���3)�z��q��'6�=�7�ˈY�҅p�b�5	�Yy�F�)�O(��/�i	do.DN��q��]�D��W�T�r1g�8)��"�,i41Gx��M'c���
%"sP>!�A�;,��P�E��[��P�"OJ�=�(H"*.�=e'ԓt�����ӂ!8`���W�"~�3t� g��5%�
���D��u��$�&U���#Q�4x��Mj���L�z%*aE��l��n�<�g��*�k���)����G&�\bf$�/�.��ʟ_w�y��R ���(Q�B�H����{��9O4x�ׄސ#wh�0�,R�c`�IJ��{b/�Q�OgQ�6�أ�,� ����J��k�)��.K�0>1�L���p �r@��BQg؞0n���T<�t�'�IY(�w�Z�ȑ�C�sjx<��'�� �S���J�>1[��ĵu�Vt �}R�ݣ��R� �q�O�4���/k�l�a l5�����'
��3E�X4�*��7+�e�����X=U؞Y[��>���>	V�B�e3��)��3V]�l8���c�<i�DŌ	��;e�E�z쾅	�,�ᦡ�A�~����v�'ۨ-ysŇ\�����y+4i��1T����Nu���@)*���Ң���ř�N�Mq!��PD�{��#���
­Y�c{�O�`[֡YRP��I.ff��m��52`lF?Cz!��T������؄w�2I�K�mz*XpU�8n.��'��"}�'��X�1��w���4̖�&�8���'r���kF�2)��l�	��	�n ا���0>1�e��L9�x�[Q M�G̋u���")�>c_���!tf�+�jH�e&�!!B��@�!�$�L�Τqv��cr*�*e�ӭ;��ɳ��s�i�����Έ�;�(�MN9C���b�.7�O���+;^%|�;���]���5.�*.y3�a?�y��Ҋ0�,m�t�V,!�5C3)�/�O$��%
Q$f�A��4�S
R���ÆN	x��ĩ�E�6m��B�	1���UG�;yq��c�.��~t�1A�_@��w�y��9O�3f��	O>�Lb��S�l�l"O��c�C�|�xH�!##Iz��w:O8�����8j
��7<O�9B
,&�L�R�aO	6N$p��'y@�!�a��Sx� ����#CȰh�GKs�2��a��%H:��2a�.�8aN�Vռ��q!T���"�!.c��m�bv�' -ړ�Z&0���c"�DE���ȓN�AI�h<)�y���_$���D�A���������s��4KE\�*\������!�t*8D�0ʣ.M�g�!8Pi@%�I�B�x� kƁ� ��`�`�Tx���� L�B���s�L��V	@���#7�OX- �F�^�z8 s��`�^@ץ��k� 8�Ї�"�yC~����=e���)���HO�'͂� �ң|ڲbO��4��۟	���r@�s�<��(В�lU�	�T�5�GT`�<	������8t0���f�\�<1��a��pɋ5N6K��T�<��nG&��Ma�3DQ�z��WS�<�t [0�� i`�ê(�|i¤��`�<��ؾQ��d�G*��!��Âa�<6dE�i~
���e�pt�(Rrf�b�<����x�^([�ǜ(~ʜQe"^�<�.X�N�9�A�� u�c��_�<��⑮Dp´�� {��ݬ�S!�� ��&#I�G�Tx0�C�`$��X�"OB�q��\���0	�H�h�(�"O�q#G%{ߨDX���%<ľl�D"O
٩�N�c��@���U��C�"O����h[�]vb���@F58��8z�"O�����NG�Ժ�hڅ@�*4�6"O����H%C\ g�G�Jqq�"O�Qr%�t{r�Vi�rV��ӄ"O�ɚ���ku@M�VH�3sE�qU"O�����.WB ��U�FUf�p�"O�Y���B�!m,�!r�W  ^zh�"O4)i�I�@�Ly�bA,5�{�"O��F�TY���+�%O���!"O ���Qax�k�KQ����"O:��1�%:�]����|��s#"Ohٺ�J�"@[�2�"O�1���ֵY.��#I��a��"O���G��w=@EH���ν�f"O�T0@��E���(3J���>I�`"O|,҂lZ�x0��AȆ)2ݔ��"O\p`(؀ %��1P%�� � "O>���iD�_`�0B���FG��"O�U�����l����j	�1���yb(�
	�H¶�P�+F�mc�-ݧ�y�W?���P.Ph$�+��y�&�V�}�d״_Z��ٲ�Մ�y���xڒe��܃S�2�a"��y�G_�7'����8\�^�����y�J	dv�a��
�z�"Ux��G�ybF(�z���U�IK2���y���(v�Pd��nѺ��^��y��DL5���e�jT��E�y2�!m��*2I�x�h��ѫկ�y� L	\`���~�N�;��@��y"$��D��ys҂K:p���I +�:�y�@4 lZ�w�Խut}��H
�y2�Qc�:a�*B�p���M�y��"\�yA	�(���A�$���y��V�!:���vHIңS�y��JO�D�;6�-V���Ĥ�yB�.7�z웳�� �`�5���y©V�W��1�NO����D N�yR+�!8�a{�'��t�Y��X��y"F6D��z���2���eAҨ�y�W�`�<0HR�^9|.���
̿�yB�7f�Td��:li%_�y�)];�4�6j���|g	� �y��As��S� �
+Mԕ�Vl1�y2j�	i�����O�$�� 	���y���9/���E�+��qx�y2��G �	`��;,�<��*�y�Eϫ�2�X���..��b`���y2��`�n�9�K�*7O��r _��y2`P�$a{$�]s_U�w�G��y���`8�x:�웳s��=sG ��y�iY�e�0]c��C�:V���aT��y�J�%�2 �a�?��1�4��y���_��d"��޸+�D�tʁ�y��ߕ�&�
T%$-�.�tŗ��yBA�J��|�á�VH� �Å��y��H�Y�z�x �T z��3��
�yR����"y�7���>EƜ(RC��y2`C�i�n�c�S6&��A	��y��� o��H.o�W(U��y
� ��Qh�4a�!	G��u� i�D"O\U���]K���C��&rf�1�"O��2��L+
L蘒�a��k��x"O�!sj2:8�	[ª+}�h�"O���֍��.w���\i�у$"ODٻ3K�>y��j�E*� |��"OXPHD/ў:��@��S��I�"O@E�G˃& �"dA �y�r��7"O���oӪ@�(4��
m���"Oδ�V!á	�`0{q��!OY�H0�"O�l�d��1�`�0aW=18���"O��iZm�Xl[�Ϟ>D�BUS�"OjX��C�7l�7D[�ṷY��4D�p�*�>S�dܛ��+����5D�89ǏJr��$O�.-��Qئ3D� KЂZ%��Z�_,Y�T��u�7D��ZF� �D���Kԥ[7�l!�0�7D�t���X l�z"�WM�>���5D�4#�N�<��-17*U�.�AKF &D����iL4p F�1D�du��&D�xy���pG���6A�l�V���#$D��[`fB9c9܁�u��:v ����&D��0�&��y�^��,���,��T'D����޳*�	�C�e��iv�8D��B��ƺ��a6cܼ!�7D�����!]f�1��)Iw����8D��z�@иzlx3�)A:_����=D�DIb��g��C���u�htP�*9D�pȵ�В~tN�#m��C����!4�ɀB�����'"Bq"-�g��6.�����bA�'�@��d$X*V�R���c�*Lp� ���T��reOF�3p�T�q�(�Xbd�	3�n�)RO$��R���'"�
�ޑ�7��"H�����y�bȼ�b�bu�B=�qHrh��Px"$^�-ǈ��gm�d�|y�[�Zz��",ة|��txƉ�EF������-Ɔ��w�)]N%2#b�Y�`�F��x'�������ڐƋ4����M��_;j� �ć$�t����\���c���Nv� bJf���]C�� 5[���&z����
�^�D�'N��y�-�h�ʁ�O��n�ҡp!'a�꼃Diͩ%26 ���-H$h����J�ƴ
�c�J��{���!��)P�dV��EO �D��O̸b�.��-T���31	���")p��Q���Tj_�{<�Ybf��
��p�O��;�Y'B
P��ubK�,�p)�G<��IRT ũ^(�,��@��t��p��GZ������):�bl�F
_9uJPI;U� e��#?�5#��Q�ҙ3"������0}�4E��K�#�X�����ڰ���R�_�4ui��).����~���+�I<RB��	�;(0RH�OܶK�B�	0Y��U��=x�MZ�	��n���Ǌ:��C�!�05�:��3'�;@��q�3�Q='&$�j����=q��M�!����Ӭ]�9�A��U~�ʓM�|���ƈ�V�I#���d�Ƽ�t+W?B�d�h ���Ll���)'X�9�J�'�:��' ��"�t���
�a]�J�:���{���r�-�A�T����j� D3�HZf���d�'� 1���O%�`k�k˵*6��P!��$��Y˖�ɐn�j]ٖ�G(�E�lk�xS�KS2nx��&��;E�����͊T�85ۆg��hr8�Ck�,�~��Y6=����$�)T��B�D]9�f�3�hv���ͯE�9�c��8��D��5�D�����'y���pE�2n�����FE�=��v��e��G�`N���� =>��'`Z8xê�'M����Q��]�2�bL���_Iy�hɉ"��4�@�Y�iH�X�G���0?�c�K@AZ4	WJ�"f�1��kA48��JEG��r� ʓ�VȨ2���rΣ?���+M4�<���G�}�@��G~�'�^HB�iƜd3���'=�a;�I�G�NUy7��zl��pweDl��)$M�U��\;�2�8�ѥJ�-\��A3Aʳ�����̯W�j��'��9S���Y��N~*���I����Ĝ/�\ Ð)�c�<��] o�2�Gɶuh���S}R�Ј?L��3�|�OK���c#�@yҭ  Ԍ�o˺nI��a�!��y�
\٦mr���[��uȲ��;��[��a��ET��0<�P�����D����e�[P<�pH�2�9�d��}�`�[5(�r�8��1�� �£��'�<xQr'��[fB��"O�)��ߥc��1�f�sn�5*e"O2̳��Z�\P6�J��:k��5��"O��Wʗ
.(H�B�7<�"a�"O�������@�k���x�H�.O���
'���d^�`�EK�D��!h*j��|�!;����WkXWbB��P;#����
�8T�ȓTX,��/�SB
�k�*�!��Fx�`]��D2�	"��N@P���(j���+q'�*1� b"O����*+�<YԧU�h�H���f� <�l���̑Fy^�S��y�M��y1�43P41�5�3���yob����蘈4���S`�	�y�_l���(3�O�<�y�I+lB����?!���b&�7�0>I7�5��]cD�6�|Q&.�9�X԰� K�v ��C	�'���R��>�16gҷ	�%c��d�?g�(%Yv%˳A�"�?�b(�]� ��u�5?�x܈�2D��$K݅>��dCWgR,$�&�N��B��u�S��4ps.͖�����i溰:w����"��G��wj!���>n�� �A�H�(�GO�nA��F�6貔�
�~�f���T���ŧ(:���*׭�:8�|��\6\��|�@`��#q���V�Y%?�����,��02gJ�ow��"~Γ̾���a�<?ϒE+���B�0Dz�!�g�FP� 哺p�p�#BƏ)H��`��S���$G >'n踢�;�OV���*�)�p�[�^x�!���'jm����;g��ɯ>�y���'r�n�0 �M*�8C�	�n(Cp��#(��p��뉒{d8c��Z��K<���ө^��,�"ܭ?\~�B&k^�C�I�	>�c@�j���� �d.��� #O;���OX0G��Oj��C��#iuE�N�2�Q�"O|L{�+�<i|��jtcS�=���)G�imvy��mν_�dd�j�x�[�#�q$<x�7 �o�J���Ć��U�(�?�QIĬ�0����VR��N�<�F��c��x��#�y����!�s�?�2DXQ��]&��}�FDOV^HȫV�Ə*��e`q�Lh�<��"�(�"����?sࠥ"$](=+|�
@����	��H��IF�w�_L<�`	��Y�EVC䉐,0=�S)$�rl�c�T�2\$�$S�:��UB�'�O ��&� r�� ;E"W/"1V���'�~���N?�A�	;R]X���/T�L�W�J�<9Pjޭ�t��'�'Y��[TUx}"���<�:��%�'"-�H ���VJJc�qR�)O�!B�靃JI�%̚y�@��։�s_PE�:D�<�0cbm)�'�4U��)#��G�����v���fr��l|�P�`�lx�;���/X�b���B�8M�@I�@��SF1�2�L�	��qQdA[9���s���򇊄P#�2�A��\hz$�?D��p㘣E�F�A5MC*������f�0r4.R�,d�"_nx�xp�k�"}ْ�B���% MέQ"�O*P�D$��e��te��b�a|���A�r�B�I;�f���˻l?h��4|��#<�֯W�z2�z�����O��p����Ey�` �pp4��'���h��[Dr�T�G��k3�Zm��r����4}��)��<y�X!K�Q��B�9ot�y"e�Z�<	�_3p9Z���Y�cl
���U�<	�Ejޞ���.��<�Ť�50^|�4j�+u�f ��l�H8���A�_2['l!yЈS0SY�Pj�(Vr�ڨK��,!��*6jdjf�|x@u�҉'
��8A��401G�4�ʶ}$D�BdL�r�qʞ��y�)i�	a��B�1��!�y�BM�`�zC����� ���yR���L��qL��U��7�O8�y�m�5z4	n�\�{�nd�lF�yB	Z�M�@�f+�3 �~H��G%�y2Ș n��5˲H�KiҤ3֭Ā�y
� v1�!%1*�>Qv���a���(1"O �! ,�6	
<�Dg�|E�-�a"O��`D��V	��b%d�,59r�+q"Ox�"Fϒ�6��VdK� Z�+&"OڵR$��y�^�q�DO/��'"O���b��j��U�b�D�H0��"O�i���ĝrBzXr�Y,��q&"O��J��M��NYH$��4��"O*D�����Q	��3�H��1"Ov�#Ì12��x�W�F����"O��Aǈ4@�Z���,�@`�"O��
H�1a�H<j#G�,
Ɋ�D"O���D� >&�hH�/9H�ͳ�"O����D�B��0K�+7�!s�"O41I@�ߙ!$�
�+ �hH��"Oz�f�O�R%�+��l���"Oz���-Ә]�&�W
5w���"O㖤׆g	n�+��T�P�=��"OC�@T�9q��TC\��"ONU�a� C��uk���=6\I�"O�@Q�S�`,:�(��68E����"O,��֯΁����`\�d;���"ON)��#��U���e��E��e�c"O2}�酜͂�z��Էx�:L���i�@�1!̉.p�V���	`�`r�H �4q��	!��m䝡`�=v�4��W�X?'!���0�� %h�M�t����ȭ,:!�$��h��ٹ��)!5ģ��\�!�d�^�����Z1jQ�b�!�D�)c7(8�u�4|Gdc��E�uW!�$��Kj��%�#M+L2F 4SS!�D��j4��`ݻFdtd�ȧ->d(��XޭK���O�l���fݹ�T�'�|,�PEt3胢E)Z�l��gⰈ�yX��`�CJ�����O�$4��BB	\���L��C?
8h��B-,4��E��š(��iIa���שG�.MT��1a��e�cʞ�j�t�Zm҅CQ"	3��];�䉋ç'�pXA�ʕ�Li ��ߚ � }[R��V�TI�� ����)���v>��WB�.lt�u�Â?��D���Y{!��nڹLtP�b��є*�X,�'�h�RI
A��9:�1�62;��f9O��s�;��p�8��퓚/�"EH,V�N�R0�Z�[���q� ١�����S�O�y��%�F�81bٛm�J$�e�'X �	��y<�-�uN_>���MUa�00�ȓ1E���Q�G�F�
lZ@�q�ɅȓsU�d�u�Ȓ,Vx|;��/�"��� �Д��
J�v#KU�.z����W  y�(�T֮9�$�x�t��0D֠8�+E5[8r�2��ɂ,#0���nV��Zw�ѓq�n��ܼal\E�ȓ=���D�>'P��%�Rh�R�ȓ��z��^�o���jCI94Hd$����H��BC�r���@ֵW&��ȓ=(�@��F=U|pr��E16��ȓ|τ��咖_�ܐ��n�y0�=�ȓ5�nJc$˸2��-�5I�12��l��x�����^<R����lֵi�(�ȓ+"X�X�.F��
4'k�}r��ȓOj���K�#F)��/��]��o���� �QY��j���DJ����m�(���%D�j�T��2� ��@�h���dO
%Fn^��XG�E�adB.|*�1�A�}BT��F74�صD�,#�hq�5�C:��,��8��fa�8��06m�=w�B䉐c�9s%$è���Y֯
.j�C�	� �� �U�>˲,�'�ȤC�)� (��b��+q�� %���S "O�x�p�d�|i#5��"2��@�"O4�)V�S(+���*�.��"Op��� ��PN²o���f"OJ�Y0��]�T(q,ñ"�$!r�"O>�` +Ř|CP;4�ƣc�T�Ȃ"On��Gh�`�諢`ȗ�H;�"O���K�*�~%�↊0�B�8`"O�|SA"'.�Ah��В�ΈP"O(�:B�^��� ���8�z��"Ot���<Y��@���*5���"O2,Y��4P�[e��B�UY�"Od�&g¬s�Vl�Q`ϒf0�]j�"O�b�F*{���zW���,�T��"O�Re��b���^�V�UC"O���A��$��,�7Z�c�ЀI�"O�����בB�t YQl��֮�W"O��@�a�s��-��J�?)��A&"O��դ�<�Ѕ���Γ �p��"O���Z�z��TY�f��O�TpH"O����\4X��8���K�x|�]�"O#��>?�� ʔUf٣�"OB��'˔�0P��/7S&,�#"O`\Yt��F$A !ĢP[���E"O����nf����1eO�і"O�Q�ѫ�n%z�!�RZ�Ժ!"O���glU�LWԁ�F ��o:��"O<����<���I��ZN �;�"O�-�2�XTf1�"	�Q@���"OB�RhÍ7Q谀3%��p�Ʃ F"Ojd��&�<Eh���`8s+��it"O���r�͝)P4� �@}�p"O�qpVǋ�Z� ��WB�>@	�M�"O&p��x�QckR�#��<�"O<-���ZA1�tZ
�;+����"Oά�A!��)��y�Ƀ>�~)�"O P��?oOv�aIC2l�J�"OrI�P�ƑYH*EHW-�T�"1"Or�P�� j�L�A�B�_��B�'[�ݠ�kո.@r$�"��N���
�'\V�X0�3�Bu�E��NT�{	�'0f��既r�~j%��w�^�z	�'eH07�K���[� 8h!�M��'yd�2)<�����=[JNU��'D01@iA7�p�7��b��8�'�ʄ3�&�����Ĝo'2��'��@[�ǛN�x�A�I�k����'�]a���N��p�Ŗg���Q�'f�(e$R1�����d��JئY
�'�reI�,��QڀY��J=E��A
�'ˬQ�sk��{�4�1W��@�'�<�%�'��@H�*NlR h��'"� b�X�Ԛ��T�2kܵ�
�'��)j#m�-84 �(N���-��'q&U�G��5>@H vk�B!rYQ�'�tU�$F�,XR�b�h�N��$:�'��m��� S����턣T��	�'߾�j A��y��SJ��s9Z��'��j󣒐4��\��!�/x�N@��'/���T$  r�ݨr��<b�	�'�2=����#��x��ϼ?z���'~Z�Z!#�4Z&��1�F9B(�"�'���֦�ˤŁ�倍]��  �'��<�`$��t���)S��H���� :��aA��k8�@5�]�>�r�C�"Ox��BL`<xtbvg�S�j@:d"Ohٱ3��yG�
cvp%"O�i�Q2|#�앇v��M��"O<���mR+i
��`ܺ3vQ�"O�Y��MQC���(JYCT<J"OV8 �h "		U�;(W�Ex"O�6�V>gJ���v�Oؑz�"O.��3m��Dؚ����$2�0e"O���F��ͤ�	��í��Qل"O��ұ"V5S�@d�gI�O�
q[w"O��C�j֓t�`e��t�P�A�"O�D�� �o#^A���N�,��!��"O:a�
5[;x�I��V�.z�w"O@��%a[aq�0أaɕBUt�Z�"OƩ�b�
4�Ru5��s> ���"Ov�A�W�"ɼ���&ԥp��ѣ"OrM��M8�p�hS̙�y��HJv"O���k�H��H�0��w"Oh�IaG�᜼"���h�U*O��S�O�2^��y&�H�c(��' ���Mr�&u��Ӷ\���'e6a���+�R���J]T�l}I�'��	�-ݨF��!�J�b�T0K�'uRXx���Z�.��,�^�TC�'giR3�#1d@y�.��!�H���'�v-��MY��D�D�Þ�jd��'$D�"���&5-��j�!$b����'�2��'�ӜTt�"��V�"@���
�'��!qr̉�5���X��9d�d��'&4�a���uOtT;C�I& �x�'�b�!�d����b�9/J���'m��h�N�/Yg���ď{J���'��(AI��m.-�,��"OΑ�bo؋$e���˘o����t"O�=q�JB!���C�/�"Y�n4�"OF!aʛ
]j���K�����"O��Bm!dD���M
�8���"Oz	�eh�t"h�p��<�6ey�"OJy��Ϙ!j�.0c ^�mr�&"Òb $Q��0�@ ���X�p"O��AЁ�w�����B"��9�"O�����8�� ��Nԯ@�\9"Ox9j7�چK���#[7�D2q"O��(�Y{b�+BG�U$a "OjQ�Bd�"�(Yw ��3���T"O�4�`�,xs� "���
)�H��"OX-s��)9�p��τ?��-�'"O�Ԓ&LWPfN� ?�"O�Q���(r�x+�,U�K+�Z"O��I��J3u*nI��ׯiT9��"O����H�e
�IA��Z#���"Ozi� Du�ܢ�闱?�T�`"Of�@ ��"�n�Cq�<o�q;�"O�j���P��!8���=V�%�u"O,b�O|/������H�q#c"O����	���KvL�%^J�Q�e"Oi�gC�#R�#���7-�C�"O��Q&E]9lU� 1cȶ�Z5"O��0��-(�b��&�ۊ�1�"O*�	0�(C��M[V�X�{���W"Ol�"&$NW:���F�/vs|̓�"OL	c�]���`�>m,au"O��j�M�%q�J�s��:S��j "O� \l(��=���׋/H��cg"O��R�"���IF�C�0��Q�q"O.(���G*.9��@��Y�n�S�"O�|P��I�a䪑{T	 w���PG"O������(E�ڬ.B�c$"OJ� �o�t�a�lQ8 9��"O���CĀb�VY@��N����"Ov���[Dg ��&	%D�f���"O8-R�B٨hI��0��9�`1!"O0Y!"���v��b6�R'n�R��"O�-[vC�4#�Є��%	{��"�"O��#Κ]%&\�3�ƀ���k"O���a�q����J� .�����"O*l@�ą��Aϒi���1#"O�,��'F�-<hm��#׫9�켲�"O~A(�ҝ$c�{1X�p����"Ov��� J7����=-�P��d"O�(9UG^�DR��#��M
���"O��f �11�����6M��,�yR���ߊ����xH���J�1�y�%��;�Qۂ*�[zm��T>�yR�FU3�ڱ�˕x��2W�΋�y���BkD�(^���V�۶B�p8��rKx�.%��y#v3��a�<�$d�����g�O|ABqk�\�<���>0��Ҁ�2Y�P�d�m�<yp"ą'P����T1`�N$��#@g�<Q䎊�2	J��f(0y<�Q
�c�<	���de�hӵ�V-{�ƍ!��ZI�<1��@�Z�����,N���n�H�<�3�7�d� �_̼`!�D�D�<	��mxU���,#6D���K�<����cB"���ӳ�ҵ���^r�<I�ᐴB��e����+_b�5�j�m�<�T�L�%V�ȣ���l����l�<Q��A2_htq� E�D�X�����h�<y5&N�������].Z�����LI�<��f�B�:��[�9S�9��`@�<Q�f��.%��C$����r��}�<YQN��'��DC���q��x���D�<A��"�f�� �?A��꒩C�<If��s��9{v�Y0��H{�<)��]�/���$HǗ
fq�mEv�<)I��_>Yp�`P�/
���h�o�<a" ]:��|�2�F/>}1��[i�<)�ˇ {���k ��	dpa$��d�<����_X웱'�o�<�h��^�<y���a��H L@t���Z�<٠)Cr����!�ds���U�<)F�8P�����?�Ev �P�<��.�M�0h%%��T}Px�v��F�<	$C�8�\�y�+N<*�&���E�k�<��2N<�`N�L�c��S�P�tyw�r����?�}j��?y�46�2a ���搉t��+;�4Z�_M���O
y3��L>)�f�3 xE����O��V��!u��#��=}Z�l���U�U��Ybw�;�ө�y�/�"�lTP�� Ѥ�bd`�=�d�D�O�|m���\��>���cj^����������+ׂ!��W�����1.i�!'e�!T��e[�θmq*�'���^�m�ן0�ڴ��I��|6�ؾ����Ê�Zt� �+){����0)t�<l�Ο����%������C�P:1����!ݦa/d��֮�
?W�e:��<Xj�@Ō��z����$�Z�nڼ&�h)!�v8�\�l	�����Œ ��B��^rb����d'�����T'��P�Q�h��Pb�#8<�"ƌ�
ېx"FעY��5b����#��b��$=�DS����Iwy��) ���)� p��Oφ�j�j��bf�j�������o�i>i���da�՗��2�� �L���(v�v��Z�G4lO����A@�<�6��	ĶL
T%j7��J�N�T2tj"j�8t0�p��e6�Y�ҥ�	ڟ��3��f��`�"|����2�*faJ�	wyB�'��w�O&�
ҏK�̉se�D�v�%�
�'�FlR�Re�c�S�O�bmR� ږ�M�۴�?���,��&&?U��6��O:˓���Td|��4�[�w 4i�lݹ��O`����W��Ob��+�	_I�P����)���[ܱO������,O5���'3�'�+�,Ob�y�b�%���)&��.{�2�'��O|��LZ�h;�&�+B�$���i�1ڼ����'�ў�NR�M��<��ɰK��
��؟`N�z�Cp�����>���/P��0���(m����I��@��2�MaӜ��<�O�b�'���i�<�A�BI�8� ��}�kbj/��O�b��L>i�nR`v��
��W t���Rɂ�n�fy0e�ĴV���i�'U#}�'U��
��[5*�r�L��1�,-�S��O���W`y�����R�r�3掀�U~q�� 0N��`��c�"�'����"`��ICx�9$��6WH���{|�8�oZU���
�4�J�``�1C�����;v�<��0�X��i���'��|�O��vgG"(�������u$�mq��Rwwt(��J2�O�1J!+H	U�"Vˈ �pH�`�ij�� "CǌP���X��'X�80a��/Q�́�@:&"(��4&X��ٟ8�J<���?H<9��@�n.� �f�XF���B�X��-�O杓p<dqC�G�EQN���dޱ�M�O>��i��d�|��c�6 :  �