MPQ    ��    h�  h                                                                                 �kI=:�	��iX�D�l�t,��,�r�%��,}�"�&�/L��B#�*~�}tU:�X�k��1D`}���\�*�oh�Ry	�j����Wߞ�K���Q��&���wR�wv�1<�A���n������Y����+Q[���QU�?�9[��p��"Y���t���w-OL/a�A��J�� ��#d�m����t�g�����#����^��W����}�z ����\�w��GW�����M�A��V���7+��W��t`�O�O��l��|�uF��J礳zE��Z���_�q^����/��s���N��k[U��BhYOjd�]�����J!	�E�g˴�՞5�eZ"��k�'C���L,���aT���I�ӿJp,<%D�d&7��኿}���X1uM{A��������-@F�@-�<�x� 'a����Eb@��V�v�5f2
$a�U���^��Pp�_�,:�K��u���1����m�
��=b�����>M�-�k@����%>	��I�ȃ2�a6�YMS�{�h3N�u
0�9���טA8�X�zq$EN����hao��s�RoEt��h�:{��v��u%�#C�E�{ ^#������짬�[lJ�9�C}1]`S���&O�%�P��4'e�O��g�<EI�f�MXZ�Gl$��]"i���5/e��N$A�t�F�.�S^ϵ��4��h���3���s�	u.�+Ш����O�yf@�w>2��?�4�!�pմq�X0�b2��}���w����Vw
&Q�P�<8F�p�+4���s����|��}93�q�\��H�@�2������Ô_��b&M����{��Z�8�F��JU�Vz�G��o��i�P�q��͜���;Z�eTL�x��)t��\�I��������H�Y᮰��j�	��7������ч��di>��.���-)t@��R�G"]-�R
���wf��x�A�ۇ��==��P�){Ls�׻�]�������t�87��6'dB$1�qs^�{��ǁA�tX<��0�5�B��ez��P}��Q��r\M��6]ĥ�{�	=���.d�(��G$�p=���qQemi$iT�k9[^�o�m�|I���Y�ܟ;M��i�����������H�b��Uco'���JnE�TR�5��KS�J��9��&%� ����SqkòI�&$Ad_�c���6Z����R!CD��@x"w�٫YfŠ�{�hSUW�4ڵq�-'�2��
"��"^��q��+�ϸcA �'�*�bZ�ƝC�;!��7�He;�	��O^�r����/ �O��1k$\ĸ��@�4d/}�ύ��T�'.��l���6�V�~��o;�멝0	a�+8W��`5[���WX ���e4��M�w.��2�o&x|'��E	xUz�`����{weu�ƺ�\�Y�ӳfkQ4����ۤ%��3�uA\��W�=�e����0/����ST�놊<�K�z�������G%��rv����t'�;��߀��=6\4��<�W�|�� �׿����7����B�0MZe�`�\n��f9˩�����x��(�N�RQ1�Bd,�C�T�𹩍�L�K���琷���kz��E/�Ă?�-�L��m����ˁè��%{�"8�TO4�1��28��=�yL
�D{�n��Q*ʧ�Y֩@�:�߯>����$�gQ��{u���	����ermhy��Z������lE�4�c�x��������7q�;�{��[Y{\Q��s��F�XFK�1r��Q�l�0�9i�-��O�-xl��g�YEŨ=z=fL����2�*�nN�a�{;��xs���Դ��VXk�P��S4Yc1X+X)�K"�S)���v�	ZH�pH�_*��A0aP��1P7�Z?視��/�bzշ^r�
ǡF����
���K
�V�����Pm��+޵�	=���#����(���d�����c�8l7,�-m�[��̯(
��y�urG�e�S��'?�v,�p��:���-#�g2�N�����ۼ�c=�)�s�
 ��W�Z"���d�u��W� �6sV񱅞��DD ���Kh)Mc��q#gd=\����qΥr���`�>��O]���pj&�l���I�ҹﻱ�,tӪks���b�Jj�1��/�87�G�X����\����Ǫǉv%\I����$?�J8�B�α�}��L��rӳK�5�msH�3�D��s�ӑ���2<٫=nz~�>�:G=<i��<yP�a���S�R4�E���F�����\cXu�(����j���^|�U�\s��g�Q��A�� JxS�����B�i I�a�ƨ��L;V��y�-�A��y߂YB����y��=��҈��)w�M�e�M���(�B.|�~%1-J�:K)����)塮��ŋ��'�c�$�A-e_9zd�[{��.Η5갴��S���q�o��QgR�Rt`���Os'��v��%�I5��3X��3VЯ����#|��[�[��
|��I�̠��;�O�B�e*�]3&�����qi2�p�d�(Z�G��)������m8�2 'я��5�$A(�~��9J�.����P����03[Њ�{�^������c[��^s���8b� #��$X�:�S�Tt�g���U�����+��g�6�E]����`G=w5�_���0b�A�i@`�9��zkm�hT�i��|���L�\Ƀ������?}��:�r�8�@g5?��k�Z�%�s�Ul������פ�5ٟ%���O�4�e�g�6�Z�����B>���@Eu��X��T��U�>v���鱙iy)�VRҎ��J�y4�]�Ϥ����hED�����Ұ�7�
�@����'���z���eQz��p|���D�X0��.,�� �8��y��q9^��!Ѡf;��"��Q0
I�����ϭ��z����z����k�Br]D������R��*��k�=��r[�[�������U<<�s:5�Q"�-I�k�S�>i�n��kA)4�S�R�ZP��av��MB�p)�e_� ���5�֕�`V�*c+�f�&Y �3��k`&�'+b��|�A�KD��)gC!��C�r��oҞ�a@I|���W��9���̅s�H\B7��g���O�?��M�>���藟�@CF�ޥ�".�ĄǴx@�#VX|����>����܄���CD�S��whUs/\\�����# ��B��m+��o��&�����?�5ŀ��2��4|}q�w���<�����o+��E0��?s��T�"�Ƃ�ȍ�o�+O�2�7���0| �ك'���Ev�'���W_�в�����C� ȓ��w��)˟U"�hTiCd���ӑ���e=���C�ˏgŞpbGZ��*��Pj'�>�<:��h�T]�=�$�必��A̕_֎7N�z"��J\uȰʓpu��'}3-��@(��<M����Ly�ʏ,�������v��@2��Oa��4�D�Q��ęz޽,��N�w��3ȗ�?zm��D�bTΞ���oMxDLk^�-�h��������ʟa7�"Yȴ�{��'N$4�
��y9�]����o� �q?΀�o�ҤZo�G�Ͱ�Eo`��%:6e�v/A%0LC�,Y{; ��d�V��H���['�|9���1�QkS�8O&�T��m//���g�/uIД�|�X5MvG��$�)=N<P� h� u�N?<9���E��SQA�5(�� �i�3i��)�	�Q�+�;���G�6�r�އiA=??�!�{��� �0�A�m~;}��4��F�7�P��>&l{շ���K�$+o���Q���{ɜ�����=e�MGƚ��m�ҒE�)��^D_0�Y����iZ�d�|	�:eU3���B�oV̕�`$������!}����Ee�bx�?ztO[�����::��7�n���î�j~T��S7�:[���Ѣ1d�n���n��I(-����HXG}ۚk���V�_���+���b=�P��qL�f��^IX�� �g����5�qx�B��Jqn����<�b��k3<l�u��)���I]�}�p��0�rOޮ"U�]?o{��س�2ɲ�(�X$U�Q��%qql�i�K�F�&^���E�I���t���d���m�������g����U^'��⾸J)���oLQ5'�_S���6�����0 �U��5�k*�IIA��c��6����X�!>�����Mw��8Y����N,h.D�W��:���-"4�!U."C�^�m�/+���c|���¤��F��z)�C�a`!�@�'��;Ģ�3rʱ����lė���O�ً1����3ol@�x�/���W�B�Чh�^�d6!Q��~��;ʵܝ��&}e�E�y�r�A�v������W��L�-�o��3'T��	��2�ۢ\l!��W�e��������Ҏ9@��>�h��, �uܮ��R�1�� [�A��/ �����a%����Wz{NJ��&yG��'�-W��t������߻��=фM��x8W8���B���\��ٳ�ӓ�}�HM���`� j\oT��!�4���[�.�ü�E�<e�R�/7�=6����4b��a"LC�C��.���z��E���:/m�����gw/m&m������Ȍ%��8¼f4&x5���Ɂ��y�9;�n�$t*e��Y�����"���ε��Y�$�頄���<��j�cemkԄUZ<(ۖ�R7E>�c�kg�Q9��>� ��#�{M�GY�~�Q��s��_F��+��1m��Ϭ���zOi�����xG,Wg��!�C)�=a���B�Q2�4_ni�<^��;�u(sǆq�o�Q�r��S���1sW)~��K�:w��3�n8�	Ok���^_��tAKx�Ԛ�lP�?#,z�$\I]:���1
�q�F��P���O�s�KEI������ۘ�zs�+���	X
f��a#x:�c�����J|�M�7�e��Ι�r��(�ٴQ5u�b�`��8h��1x%���͵�$��I#�ą�������QG�K:k�D/\مq��M$�A���ݹp=bW!�3�����u�R� �N��/4M��C�l��g��e�����'�M����;���X��]2�Jpes|l0�r'�9^���Ӆ�'ǥb9�U�,��/XP����\:- آ�����%�8I����?N�z��?���b�}-ű�vt��>15���H�� D?��*��6/0��op��~=�:��i�gS�J��ơn4*�j��l��
����u�lD�Kjo1��y�SUuڨs��M���B�" E���V���i;:WaM�x���V��4�A�����r)�>(�y��P"^A��EdwX��� u�M�nD��KB�K�~.�-�zbK;�2���<��������Scb�AH�9�Y�[VDG.	��K����[�,Woh�rQ0J�!�_`{IO�rQ�t	%�Or�*�5k'�V�7>�#W��[�3���#�D�k����;<K]^���x3�-,���k<���u�G��)��)��8~��'���*)���ݟ�W��[l.����|������3�G���Шб¤���y�_�\���������խ��Oqg�F��|��{�9.����q2�]K,��[�w��ʆ�#}Պ������T�m���d#1|�L��ɞ�U�8A�n��2��r��f�;�$?IG�{dَ�mlQ���qc�߭�5t��OO}� 0��QWr�TJ��@u��WE��X �nT(g>��T�˟����R�1�*�Pj_J�Cy/У����_ұ
�DqU$��&��UP�|څ�jd'tkz����.�ẻ.��n�����/�0�+{,G�כ�4�y �q��ϓ�z@fv�$"`u�Q+*��.����X�����y~���D��������]?���"�Rl�&���=L�[m������)d<P�n_Ss�U�Q=��I�!k���>����H9�)/k�ǭ|�l�a5�����mp_Y�ý%�5�"b׻! *b�f ���3�ׂk�/��Η��fܜ�3K�O�)���!lŠC�3��k�9��;+�4>�Wm^�9��� ۥH7^X7�-I�g����E��w�$->����cJ�{B�C���c������ӷC#���� �S<t�ru����2�	�N!w���/�Idw0g�@H" rsb}�m����j����o�ڙh�����L��fol}�搃p�����*//�#���C��w�N�]���3Y��j��OZA�IƗ�#;
|��&�����|3E�,��f�_p��c�5���坛<}��{��dJ�U�B;hO�xdY0��LDﱀya�;��j����Z<����U�'�����k��؏wTؓ>��1��z�r~�Z��7g�5�}�]/uC �Kz��b-vu@#-<����v�Չ��;�}�e��vlo2MTa����䤷D�{���o,0�=�R�n~����hm�L�f��b*���M�z�k��Y�h}�7����]��	���aR��YC6�{h��N_ 7
f/9�$��Nng�Α�qZw��k?�� $o$��K�6Ej�F�l�:�aQv5�t%�2�C�3�{vC����⥑�]��[�9S9�!D1S�Ss��&�A↝�*W��Qg`B�I':k����X��G��i��<2�.��{��� NZ���j�d�S�DQ�Ё����8�āH3$�=D�	k��+����2ȳ���#�m0�����?�{!��W�g�!0{�J���}E8��������n���&����2���&�b+��������"�3mn����>�q��N�֨+d������H�_�1�֌��U�����x��u�U�9��=�no� ���?���[:��j��P�_�e�qx��ft��5�8��U�&���@�â֮&�j�w�8R7Z�"�E�ѽ�pd_�a�hΐ�K��-_���^G���������/�ڏ��6A��h�=s4iP��dL)g��U������z���s���BZB�qi�Z17��NS���6<���7��)>����}���er�p�=�P]�~K{�E�3�d!�(�V�$�SF�{��q��9iح�!��^:t�I����! ���^��ޫw���vM��ݘR�UY�h�=�J�f*��fn5�@ S� ��qj,�\d3 ��t�>8k�HWI,�AZ�Fc\G�6�;���خ!9 o����wsk)Y����B�h	�uW���A\�->1�|��"�e�^�H��m�+m�&c��:�]���I��լnCWP)!���;�;�[9n�9�L	l��;җ�\�O=SI1�f�ĮCo@��N/�y��c��;ϧ�d0�6<�I剝l`��;��fL�!��tI�р1��F���q��[���v��GJ�(Fxoܶ
'�	���VX�G�-�W�e��ݼ��T��I�]����h�Z%
[*�uw!(�MY��#�Rr}�Jh��I˜�<௾���z,����@G�X����F��6�t���;p���\=l�~��ԒWig�{���救f��]���M��'`�G�\�Z2�ܼb�D����×�T�w��R�N�8(S��A�ʐ���U#L�cȤ���SU5_��|��/�:]���پ�Vm�/t�hσ�8%���8�D4��Y�n�~�ܱ�yG��Ԛn5}�* GY�/��Ԏ��̣��$~�M�_+��n�O�eh��/bZ��\����E�[c{~B������D��@,-{��Y�	9Q���seu�F�*���A1hf\��r��	i1���EI:x"�zg8B���4�=\*Eߝ!d2A^�n�I`قN;���s��
���L���y�S��:1��)�ngK����=��	�	d
�&��_�-Af�H��3P�j�?^�q���5X%�B
�<YF�w� =[��LK���CՐ������}�+TA}	s�y_�#S����M沚$���pM�7�F��ƿ��(�D9��Fu�B��[񏏓���������0"���#�酄֠������ҝ1=�_�l� G����|�3e��kW|M��V/��ד���� ��V��M����gG-g�O�N� �B�5�h������c]�Mp`��l�yۿ	��T�
����`�z�bĩb�sّ'��/���� �4{�\���}dN����%�H��{��?������o���d}���Q.��)R�5C
H̯'Dr���c��Q��(�����~P[u:}�i� ���ÿ�aw��H�4�b[�hھ�E0����u��@�9j*�@���GU��!s������wޔ @�a���K�iVK1a������VFO�.[A�ɭ�8����@y������[��w�HJ՛M�3���VxB�;X~I�V-@EKߘh�m��ׇ������W&�c��Ac�9po*[1	�.D8��c�鷷��>o#�QQK�	��`V��O��b��FH%�u�ǅ�s&��V�R��#2Ț[(.�@�l�?���V�l;�f�x� z�3�iJ��§�7�f��ް�GU&�)�����<P8Y�N'G���<��/ϟ4�.��.�fD��H���	3��e��d���ݤ]�tٴ���-���'�n��WI��p�]�J��g=1�ċ-~��Pd�t����]���V�w���AT:��{�_�������m*�Y�_�g|l�Y��{wɹ�����>�I���m�ArA�l�6C�?�U���c٩�ml����v�c�|�5����fO��T�ۣ��lB��Ϙ��Z^<�T�E���X��4T���ôS���u�_����3��N�JC�y*��@O��q�.�D�9����k����@S̅��'q]-z}��I�geG�E�͍��"��4q`0��C,�׮���ny�q/3p��D�f���"�!�Q&j��Z��l(��^�?Ø�D"��O�x�]:���?��R'>f�.&%=���[H9���8����K����Ks���QX,I}�k�ɒ>����&�)*��=��7�aP�P�CoAp�zf_����} 5��J�*ٸ�f�:O�~3���k�k��]������� K�1#)�!��C��)D<���6-��mW(�W9����{b�H�^7"��0x�����tC��>�a���Vd.C�H5��X���.�.O�#�=��X��Y�h?�R5i����IeLw�b/�W�������� M�y�]�mS���e$$��\"�TCO��v9���z���}��M�~i��m����Ra�>[Ѿ��R`�Ƙs���	߱eL�O���u#�>�|�X��Un�UE��i����_�\���u�-�Ѳ������UXɻhJ�	d��@�	?��թ����E�t���Zז���z�'TwA�}�����{TS���ګ:��/uۤ�U�z7�G������u�{�&��˝�(-=�@�Z<��1�u� ����CΣ@fv<7�2�A0a����)X�����	,���-�%��T��u��mٝ���bʥ��3��Mn�@kѪ䣣^��޹���Z$�c�CampDY��{C{!N��%
��9�ש4��#@qu@�X[��|�o_R��Ee�*����:�~�vPw%&jC�Z{��ݚF[��"�측�[��-9��s1�6&SN�f& O�!Rt%��`/�guAIB���rU�X�&�G�_\��AԿ�,���pNu���ݧ?F-S�g�k��ɢM��3�_3�	���+a���m���J�	�h�+��0?�O�!�$��=�0V���_}��������,�3�&���խ���Q+���Dȩ��ٷ��4�)����_��|"���zɒ{����R�_�T�WK-��aP�Z�1��]���Ui���8�`o��?���RU�}����1��e%x�_�tz��z��p�h�-�۞w�atj�#Ù�7��*�  ��ث�d�/��CN�φK-��8�䔊G3�V����@��UKݣ�a�8�V=��P��SL��ĻԀ:�G�]�׳�XA��zAB��gqdbL�Zbǲ��gb<bi��Ƹ�d���)}�~�b��r����X'J]5t{z-��n6����(ɸ�$��6�^q�1�i��|��]�^u&/>I�(S�j�A�l����-r�판Q�!J�@�3��UT�s���lJ�Iӆ��35��S]-���2���3� ݻ���Z�k���IG6IA�X�c7o6(�!!4�(�Q �w.d~Y����U,h�)�W8oX���-�*��%�"��^�C��R+H�5c�{/������m��0P�C_�!����;z4��̵��f��*�@++O���1�7��)8�@`|/.y퍍J&��)�^���*6W�_��9;)�;@���m�g���m��0�����l���5�N���H��#��o7'�&}	ɫ���-�"�,x�eF)�ݷ�!m������h�����5U8�U}u���H?��vKL�ú�eМ��6q����&z�)ک�hG6)�����݉�t�Ώ�����1~=6ȵ�P	W���6�#�(��h��8X���M+��`|��\%�˗�T�*-t�$,4�r\3���sR"��3: =,�ׅ��i�L9�����?�$�E�w| /#���p����Uamq�C�Y��%L�a8��i4ܦ��)�X����y�t��ձInp�T*���YǢ(�K�Ưo�Ց�$�p~�:�C�U#��9ec���_AZ�YB���E4 cV����5~�t����f�T<{��Y̴�Q��ds@SsF6Ĳn1c:5�b2f�a�fiL�����x�Ngs���y`]=W�C���62���n���T'*;q��s=�Jե�G6��a"3Sew|1��)t^qK����ڤ�	�%��eb_[o�A��Ԑ߆P��Y?��}�Z�S7�o�
N'�F,4G�{����K��ƭެ��Q$�0��+�?	�D��/#.����(�5go�VA���7]G���ͬh�^(��-���uC���VR(��H��o
��Oͫ�%�I`#Aۣ��ۋ�~��G��z��{������η�`���u�fW�#�g�A����H�% vF����M4��b	�gu��	+�]]������a�Α�]hw�p[m�l�;��z�ܹo�����;�����bo8��"O�/�4�x�O�\0ȿ�X��:%�%-x��v��?r��s���M�}#�ߛ,fh�d��5��Hǝ*D�yu�<�	�l�ʉ�6c�ζC~���:�yi湜M����E�����4 !X�ChS��y��-U�u�T����j���cUk��so&*�N��L ;���Ћ��iq|SaCd��i�#V��kɡ�A���ߓ����y��}b�6C�wβ��6�M�(�9ۤB_K~dڵ-�/VK�ҥ�����r�d��;���ՌcؔA~�(9�~[��.�?��-�dз�fo�uQf���t�`1�O$iȭG9_%⻀����h#V!���a#"[V����4��:�I̱#|;�����#���3�O��O=�Bc��aԏ�9G��)�:G��84�n'�4$�`p4�����D�j�.����r��gO-3��L���uS��Q�����od�R�,jU>ޒޚ���E�Og���J,iHa�/��?��[]��Z�Q��wF����Fu�I�ڈ���O�ʢ�mŧp�Z�Z|����}�j���S���$������r�<K�1�?����l�ĩUlG���Qw��UjH5�`߭��On9��7<އM��J�5���|AEF��X�Tޭ��orʡl���E*����RWJ��8y%�7n���EձI��Dg>��l.���I���'�f�z8I��d��e�Ƀ��s�]�'�Ҙ0�5�,���i�,y6�Hq�͜��.�f��"���Q!�F�乩�'P�� ��$����/�I�I�]5�_���R��I�#=B%[#y�3���_�/F��$��sk�Qs��I���k���>N�~4)%�$�cH�#�ak?���5!p�?_�0�T�U5�O�q�*�/f6E���3�9�k���u���=��R �Ku3w)�M�!b^C`��P���o8�1Oy���,W�W9 ���	�H�kU7]�畝�o�v��PN4�>+��Y�1��C�����0Q��LL���#��R�8�I��C,��h���D�3wy�:/M����R�69� (�����m�^�`rp�7j����()��2��V���}BQ��y�,��������Y��9;Q�-N����i�+�`0�O��CS�Yg5|~[��j��ļEG߽Ԥ�_&맲�Xz�,�����4�^�N�ڨeU�o�hEw�d�����r��QZ�1��� �4�!a�Zr�'���'�[��8+i�>T��еE}�6�W��P��7������9��u9o����ؽq-�$#@�\<^I��}Z��3�1$�V�vw"�2���a�-\�U�k�������,&�ߨ!җ�J��S�m����b�Av�N�5M�G�k�����_8m���S��ʃ�a�nY9�y{l&N���
�6�9�����Dմq�)��dÀc'o�-�́�^E`vj�"�2:g�evkK%���C_�d{�&3�5��ؿ�ޫ[X�9�+1I��S)�
&;|5�&� F����g���I]n��B�X��RGXE����"�t��1�8Q�%N����`��S�#���Ġ>�z�	3�t*z�	a|�+<�|��D�����c�̇z��?pCx!2]��]01�s*�}{_���|�H���B��&�!�(�)��N�+ ��߳���8���r���z���_��W����QW��|&_A����g��X.�����s�U���3��og)�<_U��i�����˧{�FJTe�>Wx�t`9��5n[���R��K��yl����jO�ƙ.�7�r�5 ��dU�h��w���Z-��;����G��$�>M��.���&��z�O�s�=���P��>L�����q� 
5�ا��N��",^B��q_NZ��-�m� ���<��M��Y ����.�}�5j��*rHR�s��]���{Uy����v�^�(�:�$f�ϓ�q���iǷ��T*^��I�1�I�uk���c�'l�՜�m@��,q������;�UO���JZL�����5�[�S8zڋ�d�#a ؞Z����k[D>Ib{�APA�c�6F��)nk!/<���mw�|7Y�Š���h��VWsm�w�L- �2��"t��^_��J+#G�c-��œ�B��rԋ�C͍�!�"���;U-����ʂ ���9���sO��1�(�ĤLY@Zz/i���(Q���ywt��o�6r���<sxd;{�-��b�y�*��G ��ô�����/V�,�����o�u'���	�]L�L#���Hg�Ce�pDݲ��h#ҿ�e��ɳ���Ѡ�u�f�CE5�����3\рXl�?�1���7}/zLG��9�G���^������t��u�g!�le3=��)���W*���v��Cxs���ǳfB�.��M�ss`w��\�ǌ�R�
�Ev졟���MX��jR��F�.l	����@���]L�i��Zê�z7�k�x�ry�/~S��+̕��tFm���S�Ô�%�Φ8��U47n��=V���y�֛��(n��*6f|Y�5����>�*(L�:�J$t	{�[ӏ��#�;D&e^%)�|�Zm"��5�E��c1I���������{~D$Y�6Qw�@sQ�Fq}T�N�1^.*Ͻ����higF��;�x���g�����n=R�~�S>�2��n�k��Q;Lsx�u�@ϡ�B����S l�1ěy)�m�K��N?���?=�	�Y�_�A�}a�:fP��$?�{�����N:��/
	2�FG����gvo�K����y�Z��<����+�LF	���o #	�C�$������N97h��Ĭ��(vz���u޽*�QӼ�I���b�ܪ�&�뙟C#|��'���'��bI�|~������ �����
ފi���a"MW2{"�������� Q�)�7EMMϗ�]�g�ĺ�e�xA=�^y���P��	�G]�pV�lA�g�5�=��kz��6��¦��b
��Ǳ/iVt�3}9�j��\���3�A�umZ%��1�q�?_.����}�>���Zӟ��5T�H«	D(G6��4䑇�ʾ���~��:��i�;��7�MIe���4��`�x���_����u������j�}���T�U���sJ �=�j��< 6t�����Vi�ͽa�ر�D�fV�-d�A�R��~�o�Iy0��<��w	=�щ�M����B{�~�-6:"K�,�����o��A��Yc�OsA��f9f�~[���.�X�������=��o�\�Q�����`�#O_���KN%�!R�;	�9�V<����#�][�t�v���5
��t;m�^�w��3�U��$��K��\�+���/G��Z)��.���86>'� ��ó��f����%Q.�������B�!3Gm����8��&�#�O������֝E\������G�@(&g��t�Jc����K���"��]�}�L'iw��ʷY�γV�U6ӥ���rm`�?�U�	|"J4�8����)����������rw��,�?Z0�F�y���%l�.��,*�אx?5E6���X�O`��Q�5ޢx�ŕ��z�ʕE�� X�_T9���*�����UػµU�w�JPzy ����ϐ��d�D�b�G�f�4(v`�����''�Qz�X�ce=x���+Q����jTI0��H,X`]�$t�yQ�Fq%�U��8�f'S\"1��QJ~�?9ѧ�2���
*Q�j�m��d宠]0����DR�	��d`�=�u[���nR���KmA��]s&x�Q�(�I��jk`�6>U���bQ) �bǾB</�a��?�9p�Ƨ_
�����5��o��C�*O��fQ��E&�3���kLD'͓y�����ܭv;K0U�)Ӧ!�ڲC;��2Y�
�v,�0�Eb�W��9#Dm�q��H�"<7����8��������	lG>F,��!��C2cܥ4u⸰$����#B�� �����9���e�B��?��wԞR/����t���� ;�.��m����[�����.�ʒ�C��l �㞹� GB}���t�t�#M�[�Q�t�Ѵy��\�����ː�[4�Okk�z2'�t-�|��A�E�u�˘E�]���sR_�����B�GH��Z�9G����U�6�h@Adj\Z�}���r������\KVZ��$�'
`E��+�)�TIs�А�Ͽq��C�ݕK��7xK+�f�i�TS�u�ƨ��HK���-G,@@�<��i��#��6Dq��$ԣ�e�v�-�2qa��v��߷u���>�,�$�����a���0%mϟwE3b@�p�iȇMd�ek�V���PP��Y����%xa��Y�z{�|�N% 
7�9�9~�_!Ϗ���q�2�w�>�`o�d`���E[h�}M:"�v�?�%9mC:�{'i���9@��|�n:�[��9_k1ěS��&v�k�W��D�`g�:�Ix8��hP�X���G��q���.��H��q��N�P���n:��S=����fȿ��չz3U���S 	�e+ǂ�㲰��2��^�i�բ$?+W�!M�״���0y�Y��}����V���ӈ��Px&ؓyգ��=+[/�z�������D�d��������2*v�Yy�������_�G�͔�)��P(�Us�&�U�~��.��o��G�����#�s�|˂����e[�.x���t�l��8����#���T�/�״�j�r���ص7k���v����4d�p����c��u�-0���`-G�'S��-��I*�K"Q�U�ۮ[=D}!P�.&L:(�J8-�;�]�S�U�d��]�B+��qZZ�BQ��(�����1<XlC�|���r��y(}�rJ-r����y]+��{0�i����5-w(��1$��d����q�Y�i��^��k�^��XtkmI���� 慟�}��+��Q�3��J�i�'UJG^�NܠJo���t�5jS�6�"#N�-3� ӡ��O��k�I}��A�I�c�.6����!*
0���w��TY�e���h��oW��F���-�ύv�"/Q�^0�%�+��ch���.'�����XC��\!*���;0Fl�����hd��'{On�1�9���@@5�G/��%��wj���԰��Pԑ6��������;�1�7�ΰ�w��i�p�ޛ�bqf{I��āL�~����4o�Q'@��	�/���8 �t��e|؞ݭA�##��z�O��8��)6���buH9�>k��,����aћ $ɺm����%�r�z�J��*�G�)��.���tw�g��-Rߧ�|==g����JWze���^�u�������i�Ma�m`r|�\�-Z��`߬�%��(ta�(eRXj��)�n�.���f�0�L/AJ�5����ٟ�$�m��/�C��z�ӳ�m7����Ͻ�%�#�8���4�U���x�-�y�/����7n�E*�%�Y��o������U�P$��C��"��ˉ���neY�?@��Z(:�P�rE*�cwt�=�=���m�c�Q�{9� Yk�Q�$)s�n�F�V�RO�1YB;�9-�׵i�_���x��g鎜ů�=Mg�߮�2r�pn�,{J��;'�	s��t�ۥ~�=j(��,Sۀ�1�G�)j��Ki�vz�*��~{	�bЧ7nf_юnA��Ԇ��P~h�?�ѝ�N�Iz/�%o�
�\{Fb��q-�J��K1����S��G���\�+��	��:�0�#����O?i�kL���v^��7Ө��n��^V�(QEg=�4uy�]�LtM���u������͡�V�t�#�ԅU�ј�֔�4�7Ջ�'��qw��f8�-G�P�\Y�W�0ݛ��8à�>3� ,�K�r��Mj�C�X��g+DN�����E]�� �ç���D�]��$pQ�l����𐢹�Z~�	����~�|.b�!��_~/�������Ʌ��\&��kǰ�U%c7��l}?����t�8�}�>��5���K~5�r�H���D�4W���"��/��}���O~v :NY&i܋��1�m��ڹi4�u���,��k��c�u���Q��j[,���Ua@�s%�ƫxV�H�d 1�r�K�|#�i�>pa9m���yV�̆��WA�w.�I��*{�y7��4����wD�k�l{rM�B���C�B�ʛ~�H-�dzKp�P�Ο�=���O�h�FcN*�A�M9�o+[�.�K�Z�|�5���voTQ�����`癷O�ߏ�}~%ا�ǖNnW*VW��	��#�؀[�JֽP�0[�g�;(z\�ju�]3m{z���xTt�W���"�G�ډ)	�>���8��'��c��7k���E�����.b��h���'�3�d啂����T�n�
�*��	�H{ �V����Aq�;�xgN��[0~��%x:����]�y]�>8�Gozw�B�r�W�=@��-Ӏ)W@�vm��ƀP�t|}���T�
�r�� ��ƕ��#r2��'}{?��t��H��I�l=�|���˦�5�+����O�ނ���޽�"�@D`��w���{E|[oX��/T�t!��5�7�`������n�<�J�Ey�$;��K��΁D]���"���A������?'�ٳz����}e��^���O.�q0���,��4��s�yl��q�b��hb`fb�A"��oQ�Q����En����O��Ecۇ��,�IQ]+{��P��RX��-y=8�[�X������.�<
��tvs�*Q���IxOk;�0>�:#����)���>��Z~a�e���"pp��_E3���GI5����'��*
}�flA��w33\,k����.����Kh��hK�k)�h!Xw�C��٥ҥ5X'�C��LWY�9>�Z�츄H��7�6W�Ӽ����z��í>a_]�OT��BCm Υ����\�?��#���;���?rI�e��.�P�:N7w/��/�@=�_�,� ��iw�m$A�Vn�����څ�6^�����y<T[%}x|T�o��~���~ُ��/�!����I�|����VX�O�5A��|t��� ���E}�q��b�_�gM�Ol��b���N��/�P�cU)Nh;��d�U��8����'A������U�Z�+~�z�('e��߮j��Dl�T����k�2��sް^�F&o7Ӛ͊!�U�o�u/�������Nޟ-�S@ٔ<'�b��Q�v�'E��ѕ+v�Xs2���a��m����0UD��H,�2���{�Z���F.Tm�P�b���Mߔ
kb��T�����պk�����a��#Y/|�{ԭ@NKq+
ҽ�9ڀ�׺GǏ���q�[�|�w��jo��ͷ��EVz���pG:ݔ
v�ST%���C��{b���k����Y��ɶ�[Θ�93^31?~�S��&�6���/t7߯q�OgL͂I�"V��}�X|]�G���0{��:���C���[N�%��V�5�}|Sx�F�<l�Ⱥ���0�K3���&	W�"+����A����Y��0��?��!h���S	E0�V��<m}�z���*���&'��&�)��q$�@<+�����M��V���O�ZL�4���vC�^�֔(�L^.��0�_��N�ig�DFΌ�lZ4��aȑU:�T�)�o�t²���'�֭���]o���me���x��1ti�#q��D��6B�/���.j�J�����7����1W�)ӰdKA��ԍ��7Qv-�#ʥ��HGD}ᚴ.��d(���=�0���A-=�*OP��	L��2��l�V����T��Z����SB���qU��������~���<�e�W���o�d��}��s �r�7ɮ�R�]���{q���v(��$�ٓg��q��i6r���2^&�[��I�o�{�������cE���F�����.UE�=��3kJб���t5���S�sË]Kl��bo ��0���@kѿ5I�ewAFr�c�f�6�H��_��!%�}�b��w_�Y���Ohur�W��뵭��-	b���Ne"�4�^K�a~��+�B�c����ɗ��陧�A��CCK�!E_	��o;�Zibʸ�����b�QVCO)z�1kqĚ�s@��/�6��^���b�/
9�Y/6���u[*�u�;�(��R������@��8������[qV�������1�FVoH��'���	"��Bn?�Y$ݘ�e`�ݨ�~���5�}�+�u���Ƥ�G�Ru�+�9�ل���>u�Ѷ���59w�ؾ���z��v��;8GGZ����.�.C�t�e�]��Z=�/5���W��?�g��y���},���g'뤺NM���`m#l\6����Cé{h���ќ����c��R�
�$00N�׶C��Kf8L�8�qX��K��H�hӛ/4쏂�{b���m�y���VI�
��%��8��4�\-�Z��Hy��E�fwn!-*l�Y����\��p#$j�ؠ�
�m)�q��eTA2��Z�L�k��E�)ac�	�x�K�E[9��9��j{�K�YvTQm�sѬIF�OT�o�1Tvh�s� ���Xi���1odx�x�g$���J�9=Hf��	�.2-E�n���ԅ;�s�G�v���84��r�yS���1�{)��KD5���J�u��	��_����_�N7A�˚�O�PYR�?J��+�D����J
�yF}����B%Kl������rx�A�}+@�	ߋ�eap#�9���z����������7�	.�h���Z(,0�x>u���G5ڏ�������Q��|�O��#�nJ�����&�@��K���uA�숪�ARu�h��3��W�kW�fk���S�߄��� �=���M`�S�g����:_���i�T�wÂ^����]9DpL��l��V۫���i
�|����K�N��b@Fّ�/�S穢ɠ��\� ���W���]�%�ƺ�g N?�����S�S��}�/����/��c5�mYH�'\D�Aسm�ő����Q:�_�~<�:�piפm^뫿ðc��tS4�����q�1���f=u��$�\2j�R� ��Uܩ�s ���

�� ,�;���7}�i��ja�!���]V2���5A��fߤ�Η�_�yR����ǯ�w�����M����J(+B�:e~��-,�^KK@��Y���C�N����ãSc	%�A�q�9\�[�\~.0��RB�w�����^oHwQ���䈵�`�O���Ѵ%�M���,;�Vr����S#�sX[A���C�+�y��t�;���}*��3H��6��}c�R(��J�FGA])$�v���&8���'3���1�Z���9�A.7Kk�㺹���z3�{��6���ߤ�%���� �x��e�����C���}�6BGg�4�{#�>ؔ��БO���&]R��B�'wWk��-���ѵK���[��{�m��K�|�N�2��%4.��/���Y��r����"{�?�0��F|��~l�-�������5{AR����O��ǲ���.c�������@(wE��X�gfT�*à�`�R��K2��x'8�wJ�1Myk�yo����3D�j�����|��������'�B�zi������e3�ۃ9Iܻʟ��0��>,i���~y���q]k�C�Pf�=;"g�Q�������X�͉'� ��� Xy��d���?]&p��v�RU���=�v�[��P��h��01q7`l5��s���Qĸ
I�*�k5�>����O�)���t~����a�(O�/I	pK�)_��@�% �5�~ׂ�.*�S�f��D;��37�Nk`�������c�VK��)	�!�3�C�Y&���@�"u���īW�^9Y,��g��H~��7	��n�'��\�afv;>|��ʦ��+C��ӥj^͸�4N���#��nVK���-ԲH�>4�9��51Sw�C/~���I��� �
��j�m�jv�Q~�HR��@��yOF�bG��T�'�#^}B��j����]"��!S٪AѪV��נƄؐ�:��Q��O!Ҧ�o���|�W���x=�A��Eu���q�_7V@�
& �}
�c���nX󋦠U�#/h6��d o���[g��ܩ���˱`���ZC�]�uN�'��I�i:��_3�T?�y�Fӥ��DEy�w�A��7.
���XfƊ�(u�� ��r�ˉ�-}��@
�<o�$�Ϡ�l^D���
����v(�F2TLa��@�f����/�,�����x���s��K{m�!-}b��򞟎DMZk�k=����#=>A[�q��ѝ�O=a�(iY���{��UN���
m�=9������u��qᤚ�IĀ��DoK3��RH/EQ�R�3�!:�13v���%��C�5�{�MB����V��$S�[���9N}�1��-S�CW&���d���̌_g��I�,u�^��XWZ�G	�Х�p�ͭ�B6���N�u����%7S�4V��v�ȵZ:ċ�|3�n���	���+�L��Y��R�T����?��u!�^���7�0�Tj���}L[b���Y�e�s��&�ՙ���m��+�p���6J��f�����O$�����<����������E_R��C^��_��F'�53I���TUաr�$6ox���m~��Bo�i`E�8{��e���x�+tq7��f.2�ܦ��p�
�Mu�j B"��O7!���h�D �d�1n்+�rL�-f�U�Ь@G��ϚoO��`�Ayu�M��$H�=z�tP��L�H��o0�qȑI��5����,Ba�qP�,��PǞ ��1�<Nﲸ2��P����}�6�sry����K]!�{���Z1k*�(��G$w�.�"�q�i���h��^a/S�>�I����^ʟX�P�&����F��6��ݟ��U@���UJ�����5	��S� ������c�
 �6�$�k���I�
A��2c��6��P��=[! ���u2w��Y#��u�=hPu�W$(�H�3-;��CG�"�8�^fp���Y+��c�`��d(���=�ԜkC�ٳ!`Ÿ	�;����ݮ�S����&�����O�z1(�F�J�@�S/����$�.���k����6�������$5;,�m$���;?x/��4�Xf1ݎ�:�?��6(�o�� '�Qk	54O���
�^Z9�e�|ݣW7�������(���J�ۡT�B�u~>��4��� ���E��ѰKɰ$��f���?z`���l�G����X��I�tm�o�8d�I�=sߵ��W0<�"ˢ�R���B��"�߆�M�
`h� \�Z5˃�ũ�����Ж���R��o��M����q@��f�AL%PV��w�+~�<��c0�/��܂\O�	�&m�݋�#�Ex�%�,8���4H��(�c��yxj�Ae�n\�*�Y�����0'�[�G��x�$�9��c�Ap��$�eO� ���Z�<�� E mc¼������0��Ux6z{���Y8��Q�!s�
\F"i����1Oʱ�οt�MGi�(���H�xi�}g_���N�=C���d�2�nK@��;��Zs)����@�3,���SQ
m1 �)`\�K��� _�b:	�k���j_G.A��|	MP4\�?��u���?Z���M
:�F�|�g� �vK�J��JKn�������+���	�8���#��G��������nD7I�*�Tm�(;a��mu���Bc�Z�?��-Ը͗b��*aN#-�T���j��ˑ�sk��������g����bΣ��:7I�R'UWC��S�5�nUg�4' ����z�M����NQ�g�&��=�ɭե�op�]��E]�bpG�zlR-��f�x�ۘ��,ӧx'����bۊU���/z|��de�ɻ��\~��d�&�%�v��b�<?p�J�_2w�n�T}�͛���P��5%��H���D9o��(_̑��቏DZ�:�~wҁ:�D�i�� �C��~��PE4[İ��F�l���W�u~�r�@j��1�GfUW3s�I$����~h] '��(�Ƌ���i݀�a/����gVmk�5�6A���������dym�L;����tw���բ��M����,XBK�2~�6�-��K&�;������V"��;B�Ӏc�?�A��9׺�[x�.k�&��I�r���NJ�o��Q�R����`���O֧��C,%���L9K�k�V�l�"�#y.�[BW�G�d�&]��%�;�������*3#'�qQ®�j�M�����BG�G�)?�ּd�8��'n%t��~�������Vf�.RT)�^�8��~�3��	������}Ƥ$W��D��O�>�y�0/�~T�w,�1��g�[6���ݻ��.��!�]�v�=_qw����Q�����f�6���Cm1f��F5|3]�i0��@���j)�vж�Q�rH�5���?khL�w��0jl3�����Ac�5w����Oq�̢��;�󹫍6��ӑ�{�E�|TX��TJ���[-0�m����k�S������J!=�y�0�����,��p,DS���ؽx���uGd���F�'8�z$\���e�����Id;�+0��s,i�U�Ly��pq�wȓQf��H"a\Q���Pw��Q�B�{�0��lG�5�g�]!����RΪ���'�=.'�[��g�$���S72�����sW��Q߰In&k�u>�����)���0m�a�����p&�B_��|���5}�z�݅E*�J�f��+�z�3}!k�x��dDt����ܾ9Kazp)$r	!NrC��-<���۲#�V��W�ʚ9t�m����HY�7I���	 �j<��rC:ӆ>�]X�EI���C���'��lܴ�#a#s�jq�I�5ͼ���y�����04+w�e/9|����"�� �"��}�mZ��L�:������"��u�ݚ�/�k�A}�'ܐe&6�4������B��%�"�E�ƿ9��\P�L AO|����{��?m|jA��֑)�|�@E�0����_�d���4�̝}�4��2Q���U_Jhh1�Fd{�Ӯ�+�"�-� ˌϕ��$Z�.��p@'-��$*��z�T�r��!�(�"�+�(�<&t7��r��Ӛƥi�u%�^�m7���~�-�@o�<�rb��ԕ��ځ�W��U�vcn2�'a����dz��V�7ץ,�5�t���c��|��m�&�bbq�y��!�M�axkH�ʤ���-�!σ
��a���Y%��{�oN�i^
�"9�n`�p���0�0q��r�\����o�ʬ����EL��s�:S�?v��4%�_�C���{��ݡ����s��[D�9i�[15�S��;&'q��(�l��'t�g�R�I�V<��8�X2wGDfN�fڤ��z��HD=e�N�/��L8���AS����r�rȰ؛��3�W����	M�b+��5���ºQ��O)��{�?\R}!�I��I��0�r�
�Z}�[>�{2D��-D�.�&)�s����H�I+U��K�~���'�U��?��j�I�l���%X�
�1���e��d_����r��z~Ռ�VZR��לUp���_oӺ��({�]֭��{��2��e,1Ex�_�t�v��!Y��(����K��9���>j�Y�7|��L��_�dAB���ϭg�-	��˂G���*��֚�M�������_n�=�P���LK	R�{;x��V	�ān�f��1�B�u�qK>�S���Ywm�L�<��,����Ǩ�dK}Q�)-�r4�P��dc]�	�{��߳�ZY|(���$��c��~�q)bi�$݋Cp�^��>E�I���1�����A�KYʓ��8qTp�:�U;���_B`JF�=�,��5��S��l���D��!^ �j��`��kG�=I��~A<#�c~6q62m�!4��c�w�Y>�"��Ph+�ZW_����q-�3�Ϟ_/"`\�^��t�9+���c�������M��`�C��U!{K���;�P��q���Δ����O���1C-dĐ޾@�ӑ/UU����e�wU��~���6�5��k����Z;g����\���3��/�Ӑ+W�uAעO���
no�r�'q,	Pf��89�i��S��eM��ݞ4�ҫa�C�i�k��|$��0uq��/��=f��6��츻�+0m�^ጾ#�z�������G���JԻ�d	�t�>��?E�X*�=!��z��W��l�����0n�sO����s�M2��`c�\� C�>G���ڞ����ù���ه�R)�-�t��?�,]n����L����ƞƷf��8��^�Z/�*��?�$1,m�^����À��%S�8�4��ף�H��~	y�7e��n�.*�$�Y��]����_Α��$`�f��:3�|���eJݫQ2�ZY����S$E�Гc��������{&����b�	{j�.YS�Qc�*s���F]��#01J>�)���r�i�^��'B�xD��g���ŀ�=>��߿��2��n&0�=�;���sdjլ�%�.(��(Q�S#10)���K��+{gګN	��Hk�_.�A�����\P��?�P�a::���6�
���F�^-��=�ۥK�>����(]��[�+��		�["#u�� Q�<��$:oc7+OE7���(J(�e��*8uJ4��=菵�d�N
�Hw��i{�7r#hq�&Jۘޗ�ζCh���r�����3 �޻ۊ�ZJ�M�zW�3\��6���� ���#"�M;��I��g<�-��ػ��.�JW��8�	��́]o5pB�l��E�!8��纱r@Rӂ���Shbv�i�	�/�s��H\���^\��؟�i�a΀%4F$�]f�?��M���ΉƩ}��Ǜs]EӋe+5��H�#D�����W7�����
Xf��~���:��i�6�� �9�r�+K?4����������4h�uy��b��j����6-KU�ܕs�"۫)�y�- "p�������i�Q8a��|���V�j���A�E��Z���[�y�`8z�}�?w��"�=M�q]� Q�Bz~�݊-"��K�Ƀϭ>�y����%�y"�czwAv�9R�9[SF�.�c�q�m�P����o��"Q����~�!`x�SOK��N�{%��0ǧ�����V�p)z�<#T	X[}�����~�!1�x�I;Y�m��3����U��I.��H �� ��G���)Z1_��e8{9^'�q
�gR����f�VĿ�X�.m}/��3��Z33
ڕS�����	��2;�l�6���t����޹�Ϛ���,�Xg_��������N�����]���8Ww��ʣ�:��A,��`��m�嬀A�|����$N*�[���y���k�e����r�L���?�e��2x�K*xl�|R�5��|�5��̭|��O��1�=�E�e���n�|���:*EM=�X��'T��죡���A�H�.ێ�GJ�hsy��5V �|vE���mD�4�����0�����Ȱ+'�uz�0_��o<e)v����'��_֚�0��$,��3y�@�q�����af�j"�ͶQ�u�v��Υ��]��~�֡E�p���?E]|'�a��R� {��T�=���[j�ΓZ���f��-l]�s�)Q���I�A~k�*�>A����X�)r3�*_+(��a��%�5p��_��L�[1k5x��81�*;aWf��:1,u3�]�k8uj���2���`�rK�)?KF!�JC�Qw���v�٦���W���9����]/�H4>87�%��iP��������>�"���Hx��C�������P{�#.��_r��������FR�o@��+W�w@�3/�I�44Τ��i oZ���m�i�G�Ӈ���ڶ5����X�
��J}I-�`�n���A�G�d����Ѡ���t����Ju�p��G��O׸�f-����_|�J%�����)dENs���_�f����Lĝ��2���E�U���h,� d��iEԱ=�橘���g^�H4�Zy���k�'v�N��9_��!�T5]���&��]&��q�7��7�Hu�Rn���[Xu��H�H�����-���@ �k<%M૓�Ή��7��fq�b�v���2�a�K{�jn�av�R��,����O×���m�#)�F�b,,����!MPxAk�-��Fzt�<�	�|h��ŀ�aElY�@/{e �N��
��?9�$��z0��-zq�9�A��io��n͈e�EGp��$w:�0v�OA%WPC���{���<�������[�o�9��1��ySpG0&b>��-��W��{�g}E	I䠫�T��X��G> ����S��z���Ne���a՜S)�q��&ȫv��Ao�3A`��	���+�R��ϫ[��H��Jo��A?�!�T����^0x�4Eȯ}�|2�vf�������&D�lՏ=��#�X+GY���-렟�%������1������K��C�E������.'_�������J��<�s�����UE�@:o.�����N�x�!�_u>��̖mĪe��|x���t'� �ܣ �˾�������õjV������7���b"X�z�d�rn�e�3�袖-�����x�GU=͚��Iֵ0�7PJ��ۚ�=��P�r�L��!�6'D���R�?H����I��B��qF�E�����کg\�<D�Ҹ�](��#5H�}z���c�r�ܺ���]f�{����������(���$-]y���qD*Uiw�4�H^�����I��*�W�΢4�\�BԼl�sz���O�ղ�U6g�����J:��G��5�N6Sډ���홱i ��t���	k�'I鴮A���cY�.6m���0�!���sp*w�زYY���kjOh�3W�D��~��-�L����T"��^��G�%+j�ccT�Ś�������R��CtW�!���}�;��Q&dʉ
���dƗb�OZ'�1^�����@��/���/R��ا@�p�<�`6��l����]�p;��ǝ�'2��$L�������Jxq�N����������doY�p','�	k����ΥD�V��e�9ݙ��L��f�^�����8�W���u��5�*CÄ��"�oGa��ɦ[��9|��^TzS�̩�.IGX���pH��tc���ߓ+l=�I{�u�W�s������.���Z�'�U]M��`^�>\G���������Ô#��8RĤC�F�_���� ����L�ȡ�e���r���YJt/EAw��r4�?�m� ݋e�û�%��8�|4�2ݣ��h���yn%���~Un�f�*=dY����m5X��<����:$��_�\�S��֨�BYMeE�2��Z�ږ��/ETcx���)+.�<m�����{%�;YnW>QޞCsb&1F��*���1EҘτ�<���i��[Sx�g�_Y�=9#*�6�2^�nAq;6��;���s����G@c�)R�䃺�S��1K8
)V��Kձxf�c�F��	�v����o_�M�A#�m�r��P��?��j��@O5�q���"
�GMF�`��]�~���KK&��Zi�}�i�RF�+qe	0�ֲ
#P���;��ז��z3�x,7���`-�J�(��)�vu���88i��	�	Vc:�͍�J��,&#�"&��"d�ك��)"e#p�� F�]}D���M�x݊p���Hu�W����b��gN�*e� �-��^�^M����D5�g��8�k������^�����0��]
1�p=[[l��ܯ_�W߱��]���0�bt���/0����J?��Q�\���z��ǜ�L%�5m�XIN?& ���-�Τ�}���NU���X5[2H��JD�)���p�0^���^��~�:�� iȯoT��;��FfA48C�e[���б�Ϙuutc�F>jG'ܦQ3XUM�Cs�B�d��6 �ޅB�hJxiCa%������V㉮k�vA�9ߵ����y�<����X<�w0�G�؁�M�v�[��B�I�~�-�NTK��g�
��������ԑ;c:ՒA (w9ͅ�[.��.�Y��#�5h�ѷ_�o@��Qm+��n`S(O�L�鈣%��N���C-�V�����#/�[�㺽}��߆���Y;�{5wz}�3�R��S����C�ݏ[�Gr5�)u����8V��'��T�Fz��_���
#��iY.��}�T���V3n�~��ZȨ�������]��Q�5�4,)�^���8���z��'ٛg����:��;q��ma'�I�]#Q�3��whal�^��U�w��yQ��\
,T�mg��<;z|�Ÿ�ߋ��v���{��F�K�
x�r~�;�5�?!����@o�f
�l)`��s��׷��5LB~�w�O'@��M��)0U�,>�W�q����E��X��T ���ʻ��о��>ӻ	´�("JW�ZyH�����7�A���DI����E��- #}���:�'�>�z�%����e�����嵻���q��0|SR,擛˲�yط5q�'��I�fN��"8Z�Q����x���ŉxm�q%x���s�����6\]g���CRD���롅=$�[E�����r��K("�F��s���Q�Id}�k��z>|��� &�)�]ǅ���I�a2#��|^p�3%_1����iQ5s�ד�R*���fعq���3�^�ks��͚k)���+�t�K�݅)ZD�!D)nC�����!��O�*��WED�9�x!�ؖ%H��7�?��?�פo�r���bp>��s�;^�S��CYU^�;����<ʹ��k#�P��C�+��eYo��/�
��&�w���/�7XO�ؤ� J��U�m�:'�B�H�YZ��q��ʟ��ӡ��CG��}�RD�[�������3��7��T�O�`�5�E�^�B(DO2�R!�����y|`t���#��;E�9��^�_Hᙲ;��Ν�s`}����<�PU���h'�d1{��$�`�X��=�Bg���Z�̉f�G'�U�ߚi6��H}T�g��׀_���4J�R�2��7?��)p��mlu2ߓ#!O�:�m-N2�@���<�G��N@L���]�W�=��v�E�2%$�a����w�·�N�m��,~�*b�F���d�m�T(>��b���Mˮk�3v�@w��������g3a**Y¤{@��N7�a
>L�9��#�&!)����q2@�hOr��_�o�X�#$EBx�D��:��v�%�nWC���{N�����2�a�5�y[���9���1+HrSK�4&�+��^��c�ݢOg8X~I�
���s�X�G�6楜�6�FH�S�����N2� �B	<�GSd�}��V�Ȧ4�Ĝ�P3��STN	C1S+^3�
�h��w�E�?����?ҙ!���?�*0Sr��}�>�q�P�j���J�&_�
+���+�}F��ُ��`��YF�o����b#ym�ր%������_c�nt����6}������M�UU�Ɲ���o�C)�&������/���ּ�	�eb�Lx�?�t�U��N�-�����ۛ�0��j������72�d�6ѕ�rd7à�@M��#��-7n���PG�ܚ�q3��Ș��떣�����=K!�P�SpL�q��2���<���.f�Ʊ����0B2�FqAv�	��τ쩂��<�#��þ@��=�K{}u߹|r�����]���{w��I`<�(��$��n�S�/q_n�i������^��{kI��+��2��ڬ�w��O�ѐN��nC�p�:U1?����J��d�b��5z�WSZ�֋I,��4a- �����wk�6VI��A2T�c4�<6�U���-�!�N�Ν�wK��Yt����]:h�=}W�
�	�-����T��"�^���j�+E�cc�\�5�:���bԭG�C/F�!���z�;w��F���$fc��3���O�O��1yowĆg:@|{~/��2��������C����6N[�a�8�v;�q��>Y������L��~��e�[��EªX��C����� F�o��H'�A�	�*;�.�u-�٧e��,ݔ���U�!��yTȽa��2$?3^uO6��%	t��P��*x[�")T�!��7��"z�٩���G�[���+Y�O�t�K������L�=D�m�p4ZWAn�S?=��Lܕi�J�5�2됫�Mhə`Y��\��˴�e��̨�����o��OֿR_ñ�8���?ע�v��v�L�V��|L����,��T
/��Ă�Z-�Z��myî�@����f%���8��4Y��F?����y�25��;Un��*�� Y�G����P��:���7)$V<%�7�Ï�9&��#we@����Z�v}��s#E��vcS�ߛd���qٰ�{���Y���QY�hs=��F�tEY2�1@�6�����~��i	+���Px�[Zg�Ŷq=4���u��2,Cn\ҟ�&;n��s������$����CoS��<1f�_)�j�K�pQ��T���	�w����_x��A>�n��� P�97?6{����0�ȷ�U
k�F�U�������KX�A���x^2��Pu+,o	K Qc�#+y�v���r����%��7z� {�����(�!d�)u�/��3y�kK/����~���%�Bj30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��*I�HO�@kQ����^|�e\J4��\2A���;٤����U��'qH��N�,}�(0��qp�2aΖ���I��6 �*�J��#�_���q�W��83CS{`�!��K�$sL!��c��X���/g�BX��w�u�tKN?����K=\J�\%�	�fؠ�X�2�}���I�ɲ�dۓ�YP%���K�_�$)!�)"���������/�1'�g��c���-r,���1���Q�ϐ@�&ٍJК+����L���מ��}��if35zǂ8�������R��*����Yvf�	mKǡx���6�o��aJt��� 8��),�/�Q����x�Z+���E�$�R܉��0;iw�H�l��&5R�S�_���^��g� i�d��t���,�����tm2���ܣg��Jl:Ρ�㻡��OA�f��t?o%1���`�K��.ԩ/��Aj���Ո²i�j���ޮ�κ�����i��A'(ǈ�Ɏ���G�����m�O$,K#$��~6Mm](�6M�� ��i�xu߂�J�ci�5��B!���A��F��b��v�8P3�]���G��1�":03�R��|�-�����sW4��!g'r`��,�%�j%��6>}�bn!ˏM��6�����r�O���G�{��6��Q�9�d�{6����H7��g�rV����1Cx`����M��2��]��枯ΐ�S��Q(�"�Xh��I��٩���A]L��"�^1/�`#.gH7�{��qI����O$���ʑ��@D��5egx�7m�K<�ÉZ���Z����*f�D��j�iS���g�Ûڞu:���<VJP����bsR�Ǯ�Z���i��B�tHH�p+��ſ��g��s9qp�Đ=މo�������������^7��}IL�MKRm&�3�P��Y�-��/㗢H�[1n�	�
  AcR=������d���l��(C�C���ւ�:���0�b3yc�u:��:�u<�Q.(D>TT�B���A�g��Lyj&��PpK��@�9�ST��T�J^S먷�"�K7�<`m���uS��kL������ه���G6b��]_6ʈv�?H�g��<�JY�1߁�~F�Rs
���/Vu]]B����Ɛx�ϵ��"����
��ꕓ�5c�]A�"��/W��.��%7D°��g��}�)O>�\�c��IВD���e�S+7)?�<S�����M�GB9�f��DZ饪�־%b����1��G{�a[oV�$S��}b�%���j얙���C1�DR�0�ZϬ{ ����d��/p)p0�O=�_�G'�ł6��c\��R���9|=���bR)��36Z����w�^�b��x+�űp \G�R����&FdY1 � �j�"�9d��AҮ���4�9w���2��
��HF��z(R��:����z+��D�*p��g�����{øQY�X�W��`y�bW�\�\y���f�riE��.�8��d���و�X�s?��;{M�P|ߺs.���@o̻_�.���,�)�{6X� 	�'̈́c匄�UQ�Җ^&7�JiG���,�	�y9(�E�W2Ut��ڶ'�@X&,)�/�tq�To����G�N�GEd���b<z>�]�j�/I64r\Y�K�
#	�/Z�A��<����O\�VY���X����.�|#		5
YN٭r�^��Z�O���iv�L�{��{�;�|�{�w�m�y����Ah��Y5 6_�lʻ�F>� d{�9[{w�95!�ϰ�J�I+�n��Q�ɂ�'��x?��#�=�Y�˒JO��;�\r���
�9�1�PVp�������q�G�t(�CqK�=2�%�;PrI���6xq�t���7:_��qʤ���C�$���K��L���~��a;6���/�a�X#���p��K���t%��5�\��V%��f�X��Y}�b���ZI��,��9����%��W�\A��3�$`���M��G�
�d���Bȯc�ik�-m5��+Z��4Q븚���g�h(3�f��SVޱ�}��	[�}���fN�������H�ο����*	��i�����f�)KBFSx�4��<�>�
��aEr$�
2�8dМG�č@��xQΕ��h��Y�R\��L�(��� 1�\��R��_w]8^��g0 ���X6^���,����S�At
O���8gEyl�C�����;��A����f�tڱ�,J�����K	�I�/f�.AE�4��]`}�e@�Ss]�:��ǳ����D�e�F2�(b��ɉ*����b��m>�,����Ɠ<6�i�(��M���@3#��#\c������3����Ǟ�+��$���P����R��
��p3e��.y��M��΃�ԫZE!�ֶ`,{���jKBv��j���n|"�MpF:6�:Y�>*-��/{<F��1�ڃ�N���6)�S�6H��g���)��1>fT��ѥ��M���n$�]|�՞�D��WY�L�"?1s��-O���t t]'�"�/6��.b��7�~#�,����4>O}-���i�HH�D�w�ebǕ7�*z<�෉u!zȌ$4a܎�e�rD9���dm��]@ �~ ���V8���K���V����1Sbn7/�uK��~��pl����O�ϫ�\�`�ƙbŪ���.p�_=�{V��ϛš���q�v��Y����#��Os�R�d3u���4w��к��=;��VwT�d�� ���RX�|�e�	dx?�����U�>��1��hv��i�0]y�y>˜:��>�<Q)�>���y���g?8qyE�þ��2KK�X���S�	�T|�� �A�#dn�7Ø`J���xS�]���x��Zdv(-7^n���`9�ն���Q��ƺ��m��.-�A���{��������V�T��j�CAJ�Ɗ��ĩk�4X��45�����o�nY�O���se��AX�Ϲ]Ǧpq���n�v��g���z�t&ږ
�z�#27|�X)r�R��n�R�S4�5K�Ь'�m�i�mi����@�������;�<߈ֱ#��}���Z[�Ϲ,7"����Uҕ��HZ��Qg��Jf�Wo�o3��é"����|�4�3��~�|�t�Gh�oT�t�OX��r( N��IIu
U{|]	!\-���I+��ºp7 p�I �Ɏ,(�T��ëj#rJ�$��g�����w�觔c�K0���o��#�\��Iu���4p5���	m>Ԝ0u�U���DD!C�#���mkI4��������w����׈�TX���j���M���+&;ra���gtob������N)�s�hn�S�vp�r/���6���]�vC&�U��>^L��5?�5MQ��Ps�)�������O	n>Z�Z#�R�P��xo�V��S�9T$��%��AI��7�H��e�}��f���T�ݽ�8�*�|ى��~�5�1�ևne��j*��7���6�ŧ?ʜv���R�h�Wg���MW��׶L��gmjo?7#�D"焑������[��y�L�
���`�T?�VZ��i�y�����Y^!�����j,E�����u�D�M��9,��y��V Wࡨ���ՠ�x��E�QG�b����ii�� ���%'K��g�*�w�Z��@;�[�j�����.ʞ�ᅧ{=(�I(ZQ�\���l�8S�'0��B��{��r&��)��Y�X8���!ӷB4���Ց8Y�)CFցn%����oi1��������$S�'���[^�6\�w��ʴ �K?Z�hݏ]	m�['m@�oF�-x�lIR�5��_v�T`hcg��Ӱ[���Y&��,ea��g�5�ӎ�^�a��\A�i�x�!`��l��'�-�h��s�0S=���c�<:a]�G�o���z�^+Mj��4������#�v������8�.֗����:U�-�7]��a�v���[�\�=ѷ�T�'�$��q�����*�H�t���q�B���x޽k�ВZ4��	�bJn���*б�Hy����b)�o��hnE�w.����u3*��͏ %{<n�ۛ-لRե�N~wS�s|Ž��М|P�Q���iل4 2)ȃn)#��\�+�?��Q�˖X^4#�O���+��_,��d�Ǻ.��p�������^8�!�E��+z�b�}��<
���Fz823\]|���c��)CMs���s8�`)�c�C�8��ֹJ��/�,`+Β���hߗ���YC�#�����V��<���N1�P}p�;����z�}�gg��L~���]�1SF����©��0Y��q���VI��QQ>-�Z�����F���|�eA�$09��o�j.P�� oaEV�{�zM�7��zTE[�E��uE���ݯC��/Ǯ��Hj��z�<5�^3Ռ��A+�L��������#�E̟����;X�z&��b{~T� �y� fI,�E܉:.��a���������*�s��X�4�{��'|�..��+��@q_�r
�H�.)<�{��  -r�(�h��w�U����N��°zt�y]���G$�&
Uư&��'E��&P��/��D�x����G��h���K�в9<3F]��/���4��������.��	BE�eT�<8X�B����j����ɖK�����O	�MkN�e��L@ZĠ��߉��-Ζ^�{�� ��Ǜ`��O�b�0A��[ޱh��5�m����I��$�����Q�8���r���J�'�+�y��/*���h�(@� ���(���J�W�_��\�E��B������t75�&�������-(�Xq�12�Q\�� I�yJ6�_	��f��_)Dqn@ٶ?��C�9��@@K�n0L �F�"�E������/�U�X�4���*�KM�)���`��`B\�F%PJcf7��X=��}��h�wII�B�~Ȍ�75.%CS �#�cTL�H�L������u򲮩l�<����c%E|�-�nE�Ϸ��Q�v��խ��>���^�ۚ���j}ǆ#f�j�!���s<c�'ë�L�*-�-�?���}
f���Kf93x��`�`����d�aiWQ����8����Oı��%4Oι>�D,�"�R ��p2�¦}���:� ��R-�_�?^퍴g�q�C	�ڨ? !-,�k��w��t�'�9g��Bl������_`�A����Bwt~�P����c���S����/�9EA���|%b�������lL�y{��G���d�j�(��ɭg���)���\m��,���j��6��G(L�qM�ĝ���W#�ub[c��-F���h��B�1�*��u�XP�r�u���(���L3:��ܻ�'�7 �r�R���!&�`PVX��F9jovj�u��4�tn ��M��6Y��b������Gx{�bG�U���P$��C�6��w��H��{g�p��[1b�Ã��n�C��k���X] DD�%Ր�=��pZE"�ζ��ꘛ�˘kH]�U�":l�/��.�)q7��l�P��/�O�|��&7�l�D;$Se��7l��<��v��ȰW"tC҉Q�D��/鈒'�
ൢW�4���<$��V�*i�/�Tb�@_�y�9�Ԟ�����抰������������S�rz�p�%�=����~�E�*�O��ý}�n�|�sR,�3����؞����H���)�z,۟� ��R�����3nd��ʬ*���bM���po���U�| �0�sy⺩:t鬴mCQM��>Sџ!����gc��y�
��K� �>A�SS�fT��@�!��G�c�Ơ7*o/`�z�-kS�G��!�}����d3�@-�y,n#�`��q��ߣ��Q���/��	)-V���I��X����E�TֈQ��������́�3k!��W�5��������,YP^����d�/�ڢ~:������d��Ʌ�pn;�Zϋm����&��$���2[5/���vCung)ISX�f��D��������i��%�@��D*^�+G���R����ȩ�7��0Z�2��Pgt"�w���ΕC]�Z�b7g@��f���o[y��!"C�l����4Woӣ.�|Y)��k�(o�Ujt	r����! r��I�
y�|�u�!&��F���m1��f�(7$�AI�ꞎP�t��Κ�#��$��d�zN,��z��K�C/Z90K�:ѓ�#'�D��u?@%4�C�U�|>��0�FUB���A�!gSX���8k:^��L����ϗbe�����,�NX�15�����ڜ�� ;���䘠5��ױ�_��MK)G2{h�OW�hrS���Iщ:��v�OU<!5>o��,���٨��!T��i��wዟ��sK�>�07#ɭPI��o�
9�B�09xqJ����g?ݪ��l͸e;����%Ř�M��j7*B������������en��*>7_�&6��s?nV���x�I�W��/R9��7�LH]lm4c ?�@8DF�8�j�"�L�T�ڝH�Lr�g�Z���t�z~�F�d�_p�^E���L(gjP������& ��p0�)�6������b� ����9��y�=x���E��,��4͐V���� H��%K�������NZ�< ;+-ͫIA�(�b������N��O�(��=Z���!tlw|����g�U�@I�t��Th���88#P΁�znBX0F�y�7Y�^&Fz[�%)�9��Co�X��T���hS<�_�,�[4\0QU�����l ���?~�h�x1	��h[���9E˭��lmA�5V��v���h�������D��YJ����c3��:�5Y����4>j�e��Ay��E���>�',]��)�s��&�=�b�~1�C��a�ꠓ!��BzP��h���k+_�Gm�vt<���'�鹛�.�oj���~:y�����6��v(��[:҈�٧x����ީq��Ì$�H(Y��AԕD띋�)��r�6���C�b��e� �*t�s��vf2bM�woU0ni!�w�t@�lW*�cp�$4u<��ۿ����sܥ�Osw��|��t��t��Q0�T�����)�hTͬ����ϛL?�r�Q�?"�|�b#k�z�5�@+%�3,����k����+A��,�<8����ige+��=����}�ש<.�Z1/�F4r38�/�]��k���)g�l����s\x��ʇ�m�����ݿ����l`2y��l��F礇>�C����e�&����'!���>1X��pĆ㹍�*z'���/�!�0�K~��]�GF�h����j��l��nd���
b���t���m�F�)+�TX���w��렧�;A~}��_�U���S^��6�:mF�p��o����Ŝ��2�g� ��
J��L��mi�22�?��>�-GE`������;_e4�m�߫t�RTE�}u�#FG:6L��p�؄Z�![�?�YBT���� ���C��B�V��B����!��fёk�Y�r���xp��Շ�B
����g�i�#��?RB����pN_��yAM_�6����n;)��e�-	KB���Q�C�b�&C�c�nP��L�>�;Kܦ�ۯ&�"0��|bޤFǭ�t�yMw�r��{��Kѯ$&�|�oW	@����v�J��:�.�a	2N���-!�&���w�w��lΣ�[y���
�Jc�|wd�mo֚���R�(w��G�/�pFNP�sbc�i��Ab���ht�#�=���~˱spTb��	��l�a��d�a׫}��=LQ���^����tx�]��)��/f"܇�-{�V$T��E���=��؆i�(�Ud��E���/$��=ɝ&��� ?�o�~����/��Dmv6�r<���B��%˪"����Y~��ca����'�웒ؽ?�y[�L��
P`�U����/�&Th��5{سh�1ܲj͈���v�25y ��7��cj�ۼwZ|v�c9�� Lhn2��f��b<D�ڎ��������3��%҄�?�E]�f��YcM��V���1�~%Dy��-v��(beG(YJ ���f>+`Ѫs5s3$
�4����L���ze�������@�Ɯ�/�=3Eu(��z/�!��D�����'N`�*@�t�e�a���i1W]�x.�{nZHW�;g[�u�޳���j�h��ߚ�	�&�9�b�?K��"T�d5���X���n9Y�x�}��������t����EC�e\�oN$�5��S���<��1�w���R>��ޜ���N0=3=@�`?n��
Ѩ���It?��4 ����h���Z�uA߀�R$���%u�;:���=3�,�*�C�u�,:�G9�fFȾ�O��x�z��g/�6xaϳ�d1\2'4}`j�O�-T�;X���%���V)�	ꕤ�\l������_��ɸ��/�i~�)�±nMt��V$�z��QgX*'d�����P����M6�ֱ(
�X��[�U(�B��������r�5�΢�$U��ojO�8KX[�!��`�$��F}�L�����8��j��uϧ�,|��~ı��r��C���>	�R�H7��[άR��N��CYiOzV���5	�nkz#�$���1+�OΉc�����g7k0��l TG.M0J*O��x�M��k	y��9���|�suE���pDx�����g�
��(iZ-����j�8�E/�e
v�_iA/�=G�eN7�2�L7�5�������{,���M���:�$s�Rq3�w����8���:��,���A���=���d��2��i���*e>���e�$J��:�i�dԆ��zh�k������P��8�����*]!X�_E%�v��9)��vw�ɩn� Zo@�Rr��xѐ��:�����ͭ�l�rE_�On�~�%��ǜ�>:^,��~�LX���ǡ̔ 7��}�ų:�y���߀H�a�C;"5���Y9H�&�YKvc,�q��O�cva�Ln��H03������e;E�<]D��G��އ� ���H�
l���;���F��z�2L2z��HV|nH �\m,b����97eӢY2�p���������6��y-���0p�8�y�{�C�-�!SJ����)!��N�NR��l�AJ1��.d�C4�������ݡ춎�ܺ+m��V�k�*<�ɚ8����4�.���,�ʤ��-V1C;_�h����U��A2�QZ�Q��9�(uη�u�w���}, }��b%��-�Ո<�B��ȡMH]
=x����s}��B��pO��ON�1�WÏ����
E�ao�#�sǤ�<��d����VbWȩ�\�?��`t�Uv1q�yId��	G��}Mբ�<�8,�3[1���v���D��*{��Z:M����O�П ����9Om�>�/r=��]��,sn>�c�&1"7o�F=U*�X�F	�ڏr�[aS�*����e�d��U�s�r�\��@+r��ב�_�(�#��N̾��z�d��f,�,��!�P������Z�@��h�^q�:1^��=�j&Dڗ����5�6���k��l�@�s�yt�w&�����8¡W�O��!!��Is\��!;�żŸ��QGMg��3�������"d;qʼ�S|���c#MQ�O�����d�'��]1��+�K?����M�[�q�G4�U�� '�%l,�3�y��ո��_��~�i4p��y1���=5����*+�F���Ӳ�fRsy���[��ݎ(�s�����|������w�ԉWuz�a��`��-B�sP��,�;�����}�p>��z[�E�0�yB�z�#R(����	z�<7�4��+����^
��^BG�\�2��T�����m��N!���v�)�?�`� Lzi���*���1-A���.n����~�W�]i�E?��T ;�ňC�wDt���/��r#8�W'���P����C#��Ȏ�T��}�T�
b��^�m%P���uZ�����A�ժ*�i�b�͛��sr��K��/���hq�xj�s���+7��B [ft�m'C%�q��'���e'I+Fڈ�ߘц��C��򡩲�ؖc�u<��^�տ����e�V#���T�"|ł�;����_�^"��CqJVp���	r�v�WY0e[�T��0�)\��4 �M���J��L���#�J�֩M%>�����%�Z�J�}W�+�V�z _j�������ixw� ~$^9È9lܐ��L	�_��%d�Eӱ)�J�9�.7�Mh%l&���j��4���:�:��Xj'�Ͻ9�D�~7!@Q����S�z/��ՕL�����"����z �!��D� �qb���e��$=1$��.��� \*�E��Y��UZ�z��L[����W�\�X���e����m�ۊH7C\z9!�k��Cyg+v�Ի_1��e�P�G�l�5b��X���bȤ����y���fv�bE�2.
J�����`24�w۲s�p��D_�{n�|Ў.��M"<@��_.���5�)�b{3/ ��͕6����NU�� ��k ��\Y�OU}�%�y*�(ⴙ�3-�U�J�s '25)&ݯ�/��Q�Ef���LG������ؓ�b<4�]U�/�.4c��%g��; A	�M;ʲh�<%����=�'8���㖸h��ܐ	���NJw���BZQ9	㷉����G{"��̀���no�<r3����eh�s5����I���X�q�t��T>,K�
������JK�+����G���<�	:���O��j��(J`�T�l�\^U�����ʭ��ĕ�S�y�ɂ��X�(�!q���2Tɤ�LIdC6I���s`��E_6�q
����C"R��FK�FkL�{���l��[}K��/RCX����!nKz����5*��7\���%��Vf��8X*��}xT���	�I����D4-%�3�����Pf��r����B��ʩ�����ē1�cr8;�lx-i������_Q�"��N�ٹR����Xz�hҽ��E>}��|f_���.׫� 4R?��~�y*�',�:E��sIxf�Ks,Cx8�n��������a��۞�8U�FX��ľ�Z����������4R-^}�=��/&T��H፭�5Rb�_d�^z��g"�LlGE!-KB,9�Q�Ēt�+����gNul�m�Q��lG�AG[�!>tk�-�d��&P�����Z��/��~A���aW?�i�|s$%��&���nֳè��������j(��:�t��0�S�Em#)�,�!���@6��Y(9�Ma!z��s�$ň��wc�q�ڂں<;#�/�PƎ��Ϣ[�P�,���?��5�S�N�3���ܨ;f��6ϟ9#Ԝʂ!�D�`]�`�D=Lj�B��b�����nM�Ma�6�)�o��{$���d{�U���㬃}���6:�Z�p�Hc��g2h�����1����8��^wǔ�7,]�Q��[軐�jd��$�"��z!�w�˥�9]x��"�,/��W.1�7�y����'�O�����ޛ��4D(��eM�7�f/<Ö���mȽ���/��+D������.�x�o7��K����*�V��a�Gdb�b�F	�����?��#5��������������p�8�=
s����g���2.����
�/��c��@�R�{�3�KSŅ7�A���S���ޟ5	� ̌�Ri�/���d��V\�������,�u��Yr����0�5�y�C:a���|Q�p�>���������gp�y���hj[K�ݎ��m�S�M�TmZV1M�Tb�N��7w�`�f$���S�����%�ed@�-���np�P`�V������}LQwR��=i�N�-���k��E�z�k�G'���K��T@'��.��kn&�w�5<�X��`�5Y�ϻ�Λ���;��[��s�QΦA�^�ܕ�n�wpϘɇ��s�&KJ3��b2��/�)���C�n��Se��k[�AAAȰ�?i��9�R��@������8�����"�Ȗ4G�r$&Z,ٰ��A"]R�[���Q�Z�?g-�f@�o����x��"�����#4����_|F�,��?�o%��t��j� �� �I��t
Ɠ|���!�T\s��:����=L-;�_�~��Y}�=7Ykr�����5@&�`e�dnYAa��]'�`>�_gm�q�u���=؅��Un,M�ϜO��O��&Oa<����2�ڻ���G�nX�SiC��	l�Ec�4˜i��>���;@���5Pl�<+l����&8�����v�Z�I�!T�"��`�-��td�Z
Pg�w�fDB4o���|/�"4�B����4�����|ʡ5��7�o��dt�����" �G/I^�
�~�|$�=!���M��0�H=�k���Ûs�
�ْM�"�7T��SO��7�T-�0Ϛi{��_^b� C5����]�Ԧ�çN��t���.�0galbf$�5�tJ�y���ݖ@H���{�y���b@=�0� !J�E��[%a�/�NH�-��
;.w/���7���+��[&1ڒ��c)3d8�G^r�#ܬ(��GJ;Up����4cz(��ɔ�bTft��=IS~S��p��o�me|3�abw+��p�$�=��_�5���c� �x��<�ʱPp/��r�h�{q>4$�2�EC����)k�[i*����>���ղnF�$^�P�%TZ�:�j���@~%@.߷����O�6n��Ð��B���2	��n�\~a�c�D�|���t׵�E�Fy��,�k��P�;N�s�w�_��F4�ey��;���!�jU��h>,2�1�F�إ!jY'�w�8Av�)���y �7�2m�$�4�DEݾ�SZ���_�3n,ЄA���%WY�W�9���up�1*�Y̇[��UB�2cG���Y�:� �t+�4Ԫ���3� �4���l�td��i��@-�O�eL3͓�vj����BD@���N�D�@Y�ev��Ҟ�1�T� T{�S��I����ߙa9�;i���h2���������լ�\K�mU��H��
燏���79��xn%��x�@�s�h������g2�́Ee�kN����e2�G�C����X蹛�͜+�xN�E�3�Y�`Ǹ��ب���I��=���$ uĻ�ty��x|�u�1����3�J:�͢��:X���ZS�ٔ�m8u�q:�ŚG���FPlcO��� �4 g�� ���hf\�K�}��O�@T>sK�d��^�)vt��`#\�ں���>��͂	�`��)-5n�7���XJz$I�J�n���~���NȔ��`LQ9���k�D��=SU� �!�~�R=���`�5?�1���3�j��K��>ݩ]@��oD�X����� ��S8?%Dj?D��/)u|�u���d�9t��TX1�
ڇ�dx{	X��H��;��h�R8��[�Li��V J�5�b?��9�E���#����c.#5�`]Ok�/l��?�o[���0���O~Ox���� k�'K��v��[u}|9��E�¶�t�xm��Km�
=�i�h�jwU���E�m�
���`�l�<~'���ݣҺK7ǥ�z�$�=�4,)b�M1�t�$���q�R��~���v��«,3�0ћ^<�qX��;φ>Ì��-�G�	>JB��HJ��������kV~Θod��3h�*�D�i��Ӳ;X�%wV��ڎ�9Y@�Q�S����0Sr$p�I�:n�"=}�4WPr͚S��~-J���E�:�˟p@%L�t��O�w���J�}é�M��Q�َ���]�a>6"�\�zk�9�7�&3X��2Q���MO5a}Oߦ,��3H��) �;�K�<�F�5�fa� ����.HB���m�;D!Z�Φ���1L�[�?�=V~H���m���ڝ�9�L��
���*"���g[~������y!�p��y���95.���S�-��W�:67�tI�wdpA�C��(��^w�'�k�1�	�t48�d�m\�V%\뷲=_�"kr,�����v���+��V�;�;��h*3���l��.'Q�d�Ex�(�ݔ�����"E}�B��&���2��ҷB�:x��_�
ŀw�H�o}6�Brc�O��NF��WKްؘ�
��oqE����-�d�߅f��WP \^g���y��~D1�x���dYl	�����j�*6��L��A^18�QvAT��Y��0�>m��q!�<%{��)��'���Ċ�{���P���F��T]iL��C�Տ&���=��u���	\"�r��S	tg�Ll���R����W���ȿ���@{�rS����Z/#'���FPw��i�y��Ĵ�A�VGP1 ���,~ZLL���qW^@ =i~&�*�3���~��s�TkKH��&Ps7+tt�&0lo8OU8�\�W���(^�!�Is������<�D&��C�M�QA���s�F�����
qR4�����9��M������+
b�'>�G��IڳD�?28��dY����4fyLU�'܏,{��y<Q��1Ma�a���4��M�?�ƘE��͂�G�������F���:S�R���۠��ܞ�f���bs ��rG��,
z��u��ߒ���e`(��-����񬵴W!�-�T����z��aٸ5B�#�ї�7��z1hf������ ��_=�4F�Bσ���Z�Tk���;�G��'���l>��L�?	T �Ki!��*1AƜo޹Af	�.�\u6�2/EWtr�i8��(�,;�Å�G�Cz�D�F��f���H<��''8�PGcD�)�C��)�uZ�K>oT$���>^�P5Z;u�����DA��V�������U����͜�ӳ��	���x����Z���pUV[�ז��G%x�O��=v�WM6I�ƈ���� ϒ�~�W�V�:)��$uĖ�^��5�<����0�]=�i9�";���i�W�^�� C�C/p}�ݏ�����Y�⥫ܰ�0u)<�v~���!텏g�b�_����n�J��کՆ�Ƈ��jݐ���J6��W[(�V,e_�3�� kVj�w�$�{����ld��Ԟ�_�dn]L��1���8�9ly����l���R��>Y�����Yi�'u��93�)~��T�T��0��}��WB�]�����ت�g�k�� &>���_~�p�C=�e�$�bH��*.%s� �N�Ek�˲/���zI�[[4���6e��o�R�X����c��H��tz�Q0���2���U+�9��C����ya��$���9��"X����9�ibPp��u�<y3}�f�I	E1^�.�J���ۡ贆���UsX����4~{��|X�.�(���'@Hq�_�nd��k�)Q@�{��� �P���=?�U*MזWOɈc���:�)�Zy�(�<� û�'UM�E���'��&e�f/Ep���&�-G<7�� ES���1<��?]�;/�z�4�+����Z�Ù*	w�S�:d�<�bs�W�ί栭�3�@�{�5^�	�N�z��w��Z�>m�?@���[���{�l�U;��pz����8�E$_�$oh0L5����%WZ�b{����R��`����A�H$�J��%+���*�(���6���Ҏ)m���8�L�TJ�(����\�'����RB�ŉ�m�ۑV�Q*!���(d�q$^�2�Y�T�I�pJ6Ѵ^^#��[��_���q��g��]C���U|NKI-�LU3����o��/���X<g�����K���N������\~JF%���f.�X�f�} �|�k �IO��sR^���0%x.|�Z�����]���W�I�:����X�ʲ�4�c����16-����
�(��Q�㾐t(�A]�_b�l%ر�/՞bTA}��f�~�Ƕ��٨F��x���*B�l��[Դ�0hf�ǙK��x���5H��#u�a~v��c�8��I��H�F�׍Z�ΎpN���G弆?R������<���|Bۍ5	oR�H_�P ^7�g�=}�K-�5�LA,�	1�L�t!��2'�g��:lnu���I���P7Aϕ����t�se��de�J�i���|/�AJI���jvn�����k�>@�nws�K���2��?J�({���$�54d���m�9,C	���6�j(�1�M��"�n�A����j��c���b�����Ƿ�&�qy�*�}Pg\=�j`�ʘ��Hx38��0`��.�H�'���$!m�`��b�̧�jD�R��=ށIX�nՇ/M�V�6NZ7�� +����{ԁ{U���j�I��T����6�����H�!�g�3АBѬ1wVO�v�eJ����'��]U��㻿�p�ⵅ�0"�q�yZꍿ�-�] K�"O/O0�.�27<J��l��ux,O6��[���A�>D���e�2�7!�\<K���Z�E�.:3��^��DRZ.��ֶ[����y�)���?�"Y͟V~Ց㤫�b��]�ί��Q��O��<�?�(k�Ϥ���y_�����'��p(�'=����?*��z��������4�1���4lR!��3.�����ɐ̗V�$���4��Ǡ T�R�1�9MdQ�������$o�w\��;
��	J�qlQ0��y�d:�7�)�:Qb��>�`vv�uk�g�6y�S����Kdr5�S�YS$bT�������
֭7�<�`!;0ģSI�G�vG8��\d��h-�Wn��X`������:d�Q��غ$�ƛ��-�rX�� _��e	����� �r����wi�̶��k�i`��C5��d����
YE�)�Ve��d6���_"qә���̦ɗ&�deon082� ���Sv�&ӝ糓~�2p%G����ˌIn\��S�r�󉍟ɜ��8\i4@�ڽe@5�9Ö�����Z֪���	N���Z�ﾹ��"�5@EO�xlcZ�X�g���f�{�o�� ڳ"8�Z�?�4���x)@|�~����o��5t^������ �I"��
N�|(p�!;���?���g�[�7�ZI�(�%��3p͚�J�#���$G�o���m�耟�d�0�
HѨ�Q#�+��cSu4�y4)r&����>��.0��7UW�+\k!��L�{��k�.4���׍����b���X�'\���wܘ�ёz;k�B��l���f1�D�Y)<Yh'��O�r(���O"k�O��v��U�!�>�y����E���C��B�o���TI��о>�`�#^�HP~�*o�2򘷮9���M��rBݟ�V���epv�_R?�mU�# �*�J��B~y��lӏcue�LM*>�7�&�6�շ?#���m���>��W _u�i��nJL�nnmI�D?��D�R��_��з,-���r��L����#ޭ�^��.��/):lW�jp^v����je�e�M���ɾ��~Ë��+���h�Ȩ� 舡�H��.ܢx��E{ǔJ�����b�V �S\%`(ߒ�Z��8�KZ���;�����rɒ�+�һ��竧�
�(L��Z�,�8=�l�
#�4�����U'��)�ͬaw��8�0h��mDB-�ڴ�FWYȁ8F/�%~�`~qRo"����9�Ƽ�sS���Ap�[��	\��EJ�+�@� �xE?Sfjh�V�	��@[�^~���B��#Zlq5��xv��h|7č�C��+zY�5�ř��`/75��H�WAS���z�)��7��N2���'���A�s⑴l�=���30k���a�, (�}�w�   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   ;    މF��<->��S(O5f��p��'l��_��p>�� B8   ��A+,ɘ�I'\	~�`%Ϲ>   �   ލp�F˸���ph�'�1�#l����_�)��ToڬrN�'|V�xc���M��.���	��M;5�&��a �*���'l���t��Ԇm�F �V-i]����e
��#��+$�"<��`{Ӭ ؇N_�x�h@�Q�|��mqQ��j� W#f�4��7 ?��-ܷF3�6_b}"Ņ�R�, �b�Z�B	r�m�}����i�����~���y�~Ul���?��p����/W<PS.q���{)$��
˝l���CU�<��ǉrl�+��R~��ؖ"7�`oz�-!��0E��S$�� pZ�zc�t�<�Ív��3�֝N�'T��jC�	;��[�j��@v�)I��H�vC�I�#c����F�� ��@<C�	�98I1��R�iل� 7�љ0�PB�	3d�H�#�MO�{:v�2�δ*"0B�I(X��$y��ɷd�:(�1�^��.B�0d�&�Q�	�U4@��ߞ�B䉩f��Eƫ?W���3@��C��;Y.�LZ%�Q'%���울9�������6�̈́.��s�1$��q����]_ܼ�dyr2�?�F�lZ$���']�T��MS��O�2�(;�)�#U����Y�U�pO")�wؐ/U��'H���ApHy��SK���J}�K�c�'�|�Gx�C	�P�Ha��JX��٥�y�Gɱ[ d  �럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���O����O~��G��Oq���v�	&���b@�9�(�*oR"T�dYH<y�/��V�,4���L� �H�M��Uv���i�>IR   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ���Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   �  �  �  �  �&   ޕ����9���b��3f}�p��'l���4"S
�����?�)O����O��S�`��c��I�@T��#��n
OB5�D  Id���P�`�<��2�Q:�PxRCмnWL9 ��'t����X�;���+���?9O>1,O1�boa�mI!k��.X�#Ħ�yR�N�A��kr W����������'��7��O��LH�M��ᙦ�L.�~<��`�*J�zX��Ɵ�&�\�)�gybES�
S�l��M�5|� u*���yR��	��%�`_7&m�) D"S��yB�D	#��1�2��$�\��v-�y��b�2|��)ߤ��4&gQ8�Px"1S��hc�)GQ��q�*g�&�D}��3�h�*=���VܤyB���H�.�놠�ӟ��cX����ñ]��IrP�K�io�`�� D�|��j��a�X1a��E~7
2�.?D��#O (��2��z�'Y�F)�B��
	����U�� ~��1ၾ=/0���B�'rNHo�V!6�J�*��iъ Z�'^H��4�4�$�O��Kq�4���K��A� �޳M.�	��H�F}{B��J�������:��L�ȓ��0ѡXL���j�y��=D��)��W!���h�N��W�b���;D��sci��7�
�XU���Vj-I2�>}BE?�S�'\#�\#�@�5�bc!�tZȰ��U1$�6-�O����O���|���?үU�.<݁%a�laJM��F�s���x���c}r̄�I
k,.���+�#Sߌ@���`:�f��l꼅����H��Q��&WC�!D{� �	�R�sʍ�A��|�p�R�YP�0��?�f�iR[���}�Yܔ80 ًpv@L�t���:4Y�ȓ%w`�3�M]�5������� F��YR�|�b�F���<I����?9���e�f���3dl�����Ի��N�?�K>��S21��&�\�O�勢/԰��0�1�� /nx]��'c,8�łA�I/D)ZqK�$��x �ʫU������IO��'��I�g�r� j�P��@�¡	��	Пp��D�S��R�Q�c,�(m
�8뒻W<t��	~(%�,G�<���)TH�)���H��?�)Ot���%�aL]���%?�%-���W�XG���� �4@	�Z�'\rE��5k��T>�p���B'�Ŷ@�|��Dc�6VM
�%��kV.*�S�'Al^)�!�;9��u�A@� $�&�(�$C�O\��,�	 �.Hw�%��	Z�y��ya�� }|Q�<��	4�:�)5埠X'
��G�R"@�"=	�O��Fy���T�j 9�D�<@~���#����EyR�Z����?�����Dت,\VI��B�UP�i��~"q���9}+�26V�b?O���E�^�9��i��! H�"F�$I���'J��QB(�3�$�;k�J�Ql��6	2w�� %�p��П��	�s6x}�)�<�ߴnH����Þ!"̈́���� �>L��OI)�	[�F�̢��A2�^e*�>a��I�?�	f}B�^�\|,��_NL�P�혖d�
w0O����ON��+��~�Jd9�66J��৑���p��"G@<yd��4���c*٣x^��r�޽{�܆�����1ƥ��6���� At�*c�[ߟ`��I7<�r�n�����,�*?�B�	���,�%��X5�|� ��O��➔{�4��AZN$͓��D��D6�E;шާ�Dl(c�WO��x�Ip�	��p��c�`�0D^�I�
���e[�N��h`A*<,O����$B�!�n�r��\�|�HyrB�Q�V�ay�(U��?Q���?��4Cj@ز�ux��#��Ĺ`�VB���'�R��	 �Q�ycc_�t��h@$��wD��䙼(�ޅa���X�͊�C��n�]���O�����f�i�B�'��O�&iە�p���!W-Wr`@sf@؅����OR��ƁH-^!`�X�/4?�O��Ӛ�fD�6��7U�$]�%Y.K�*O���g��.O�
]!���Z�����N@�tUH94
rz$O��rT�'��6m��u�	{�6��ŧ�5z���¢H�c���=����<�G�3�Ը �\a��!7Ka8�0����%<�$�RD%pT��@c��%���3� ҟ����|X��� �M#���?������ h�V4'�`a���0z�HӉ�F�[2�0Ǔt�,`K��>hux��3��_]P$�>y��[��p<i�LF�Xȥ3�-�NL��{���F�f6H��}�	�i��)�<9�4w�Bw�˧h��VHn*�p�O����n ��V�37`ØA��
�>��	>s���>�"	*=;�m:�H��*��S��h�9��Cx����O$�d�<����?��O�Fݩ .�o*�q� E��MW(�)d�<�r=1��'ݨ���̐��s�!X)q���U�] �L�jB�'�Nqu� Y��1
4_�TkD�'�?!���?������Ob�T���K�nlhc/�~M�Pc�I;D����T�\���E��Bq��n5�ɰ�M�����C#4�mڰT|�o�V�1 A��=P��ŷEkx������O�d�OQhJ����;O�7mEҨ�Af����`�j����J�ay���
`I��{&l,?�L͛��T&`L�Y@��UJ$��n�D�#u� \rў�Y�D�O��Q����kh�S���.�b����@Lr1z�V���I`�S�'t��!�K�&M�
R�o�Oh@��}��0�UgڧN��5bDA"4��1��.	#�?�O>Q������'��F8�C#*B,L����5�h����4���+j�dX�
�jưi�E�;(C�	pt�s7�U(J1j�A���
/C�I�P�h�u��BT-SC�̮-�C�	�DLX��oN>DYY��U���'��<�E���r�re�ǁ�>
�2 &�V?c��C�����'^W�L��I���E�׬G�����#D�D��?�R�8�e��)�Y�i#D�#!*W+u����d��r[���&"D��s��-�����=o��}��� D�8�5��=(�ЀWO/lh!�v�*}�A3�S�'F��8Z#��1��dG��Wg�O��"���O��3���ۥ��P%�>=�8"䃚��yBL a���:��JI�FM�#GL��y�P�l)�|y�hC�+5܅I�HѢ�y¤�d`�0% �p��˜�y�^�M�bШW/��o�k≖ɸ'r:"?Y���ߟ�iR�S�a���8T�A�@�̃��E��?�N>��S���\.(�b��	=
$�p�Q�H2!�dȨ,��!b�ꉺh'�n�!��FU����c�_���D,ɉG�!�$M/܆�����e���{�� *yݡ�DH8n�(�	g(��� �2�dE�7�^i��d y�>���F|�i4 4R��I&Θ��?i��ΰ>��@ڈP���P���!]>�����QG�<!䒸Z?D�:��ˢ�n�Z��TZ�<q�"тzJ�z��Z� ������S�<�匋� �>q��A2>�<AJ��S8�0���X!���$�N�=T�ɪ3G�(4�D�����H�	U}��:U��XlL�W�4�Ű�y����u���S�jr}����yR�@�v>�T�v���E4�<Ӆ�� �y���	*�����<a*��%�ybD��y��p����c�5D���	<�HO��]���^	~��� $�$`�<M["�>������?�����S�^���H6�O�ad���&ƞAmC�-F	��(�A�\<�r���C���l�M���j�d�=�F�-D������>D��G*Z�[����J+D�$�F�I�2q�����k^�9�/$�	���O�8�f�'En�QE�������۔W��\�U��O��O���<9pJ�en����0�<���@�h�<W'ìb%���d'U��d�@1)�h�<�Pǜ�fو�PƧI��l(uY0C�I0fU�,���.�a-G,[�B��Unv%(1Ҹ�F= am	$(����=m�ޢ}BcmC�hpL �EG�woR���(�
4��'da}
� ���P+R�1���c#�9�Ĩj"O*�� �-es�ʴ��IM�ɢ�"O|A�EgJ(ix�CphN9K)��"OP���ӳ���+Gh�H+�aCc�'0��<!6`�U�67�>;kf�c�O(�~b���O�)�O��ĭ>9���9m�<p1�V%3d��%lc�<!��[�4�[�I�L�ځq�D�<i��E"<���S&� 3����\�<��蟗J@��1ū�hd�hJ�i�U�<9̟�)�R��w���H(IZq�W��h���O�l�ڴ��V��-	�ʣi�J�̠���՟���I�)�	�lR �Eʑ���1�"�T>!���.}�40Sul q3ЯO�3�!�B����Ju�ԝ~�Z��`�<q!��40h��Fb�0"�M)�/�_!��g0� ��.Ys���0�^?7ZqO��G~" R��?u�Z38�Bh�!e	�&�kE	P��|R����ɡ=c��d��5��Ā�!�!7LB䉚a�.A�c��*d��������r�tC�ɴ2|�irQ�B��ф�R�jB�ɜC|�M@7-���c��
=B�	�A�P��_�`	߄D�ԸV��
�Q�Z`�%ڧS P�Y�gT�.����`�XT;�'��'"f�1d_<A����ז2G�I�'�����K��mR��Z�A�1&wR��':L$������� qto��� �'tH�k7+L�,���#4���	��s�O�Q���w�^������D��ୟhۣ�+��|
���?��O
IA��ŪCłY��儋x�V@�#"O8�R�G���P�FV��f�"O����<̝�����O�P%p�"Or�gO�?Vٚ���oz�"O6�#6N��3�Ū�'-��Ң�>���)�9���y`��3YhI@V��6���'�L-i��'|J~:��^[�����L
4JR�<��L�K @��E
��ې��N�<q񦚶C�I�4��:{��2�h�M�<��-�
FFMZ�IQ�F��9���D�<���*TN���$�D!ݼ����@�!��xC��Ol�sĨġE̰`V�%V��ȋ��F�\&���)�gyr��4�i�Yd$���BȖ�y�I,of�x�E�q7�ߏ�y!����SH� _:՚�胰�yb�S� '���I͠}�Ё��@��Px2Fw��g�>V�ZEs"Q�n�ۥnU�'�����i�6C�bMHa,��,y`��cm�;l��ܟh����2X��LG��P6��2H�B�I)>	&4�#�Y0MW���$o�+5q�B�ɩN�6�!F�;Ll�����B��(n�z��J<WrX�(a�K�LH����T�'z�mZ�E���<( X�=*@P�'ќ請�4����O
�FD>��a�C()f6u�!c�d�ȓc>�p���M����&�T�n��؇����Gd�\�H��ui�
��ȓ���k!�,����C٪-��ȓ0����@7t��L�b�RZ��P�O�xFz��ԬΚʔ���L+-p���I&)��!��㟔%������5�?MQ e���Y}�A"O2�� $T&j�ŐWÅ�rC�=[�"O5� b�z,�@��Y�4:���"O��2)2N��Uڄ'B-Q.>��"Ox�A�⟙!�-�E�J�r��1�d�Z�'V�1��x�����ȡb�XZE^0��9���'�'���Y��p�X�,�٨�bcG�׃V!�� 4|Gi�7k�pmaAÅ7��U˱"O� �'�F�C��E Z:Uv��`$"OhUp�G�n��yį�*SnI��
O�Ep�AH*����a��n�U�T/Ҫ��OzY��퓷|&�	`�I" k�e��
"p�^x����?�
�i�PI��ɟXE������)�ޔ�ȓE_,x�w/��Lghb��`��h*�i�t�dL!E��	%Z�H�a,D�l0�,�G�����*،d�p !�$+O��Ey�,� �H���
�.bj� ��[��~��K �O���O����>��gA�`�����M��5X�*�G�<�ČޮE�HiF�H�x0� IGi�<A�"���������|@DR�&T���Ḳ$,��p�<���c��:D���0�����q�r�_v��}��g<}"
3�S��H�1㧧St�*q�nũ�.O����OD�+���cˠL:�H9� �dP���$�+�yҩXf$�S$�
Z��/ܡ�y�j�  f� ���fÈ)z��"�yRJ')�ޕ1��9s1�X��$�y�iLXa`�/#_��uQ��[����\��
�O&y�e&�&P
�J�
_�QQ�d�ߟ $�T�)�gy�l�b�q�m�:PFR7�R��yW}p�;ǋP=K�8����I'�y�Ն�mH�eәw����·�yB	�R4%�I�v8��A!E�PxrkV�������Z���x��㒰P\p�F}B Ñ�h�r��	�w�D0�UM��u�
�[�,W����	GX��1���[��Z
t8�&	8D�� QMZ���R���8dA6D����J�/e]|����3]��P���/D� B��BI������ЎX	n,O��Fyb�Z���Q�$�ː`b������~�`U��O���O���>�&��3["�:d,[����CMQ�<yƧ�*�	{p
ٝ:�,`c��M�<)�� ��i@��oG��3v�p�<���$�H2Ub��~΂����Ol�<A��'~�J�ZV���l� `.�l�D�X���O�����~4}�n�0YI(��L��%ʃ���	p�)���'�l�c���h���eوQb!�64��q�/ӾL����Ɋ>O!�L�s����B���(�R-:!��	X�\U��.��4 �`-��f*!�ĉ�ntYR@F�w5�H ���zqO�}E~m���?i@o�:IreZ�_�8�(�c�A����|r���ɫk>F��'���2qhv�":�C�I�bT�dJ�b�a�伺�d�K�C�	+Z����0e�/+���B�y1vC��3;ު�u�b쮤�`@GC�I�U�� ԍ֛!���'�O//8`b��I�?"��}2�#�&���+�e�7֮B"D\:��'Ha}�a�6nl�<�OW1`��u�I��yb@O ra���g��1��������y��Oy:H˶͊&�+ $d6���rk�=xt�GXK�h:�A�'���	��(O�$S���rP������b�!
��O�ix��i>����`�')0���Ș'��\R'� *M��3�'�,)��'?9�UH���#0̒�'[��q�:@�,i1o��,��A��'Gb��	�&�j͛'
p	BY#�'��5kҬ��ؘ%N�m$�]�O��K���	��\�x������%�8�إO=��^�����?QO>%?�K���0|(�d�
%s��Y0�;D�����OK/L��M�!<a�U�&D�� P�f�ܝ/�dx%%ٟ`�H�yU"O�8A#U
7���C$C�� 0j�"O��F�[����ȡd��-����M�'�����E��������P*�����'��'+��Y�<���������!@�T�:]YD&D��Pc%-+窠j�%�q�
��%D�x3T���98&���hܛcʬ�9�//D���H�����aF%	�ؤyS/�x�#M��B�$@z@jS�`�)�ǉ
_iQ��S�=ڧDh�B�34/�(2��RVT�z��'��'<�:� ԕrh,�@��ㅢ�y��T�RԨ��R;zP�����)�yB�g8�0;��O�}Ӭ�PZ�y/ߧH=���&lفz�4�K��א�p<	P��-X�b�
�%����3�H��UNhx���i~@�
t�'r!�^b�'�?1�����L�'�J4��d��h����4� �3��H�.�*#~�����e��Y@�T�g��<Gg(��	�(}k^�C��V+PAzM�ƻK�Y�$ $D��}{�":�3�D].x��uOz	q�(D�18ri���O&�U`p��i>M��l�R��4%�)R����D
}-X%��mUrH!�M�	/�tu������O�Fz�O�R[����.L�W���x IY��(�S��[W��xmj�����?9M>��8z`��PP�<�&��/�H��G��miؐ	���N7,���o(<Ox,�`jP?L-��N��$L���+��6��]�BتN���!�<<O�Q8���>�~�QTF��T��y�W��cO��'Tў\�>���M898QA��F!<�\�����k�<I"[�p� ��%c�nP��n�iܓ<ț��'z�I�&���I޴D����4fL���UK�&M#��Q�H�45��c��'��I���I�|ʇ�TQ#D�J́��Ƚ��=8�J��_.0A��8>ayB��Cf�G�;/�'�`�zݪDG�1*~
��b#H�M��{˓`W���ܟ��'�`��cφ@FْUO�G�d�ʌ{r�'�ay҈Ռ�4T t��QFJ�Cʛ�Px2��4�J�K��z1��JelQ�s\5B�'��	-np�y1�4Z�r���'�u'OߟD*h�Y�M=E�x���F�����O4�J7(�K�j�k��s^zq��t��S?�P�%�������$8'�h���;�d�p�(�!'�?2�J� ��ZI�Ot�@�oN~aƥ+��Ք&o�uBN<qg ��h��M�OF����Ё���wMʙY�C�l�zB�I�8�Ps�:H��cb�e��-��I%�(O�}K@m�6o(	� �8^"d@ᒉ���h�	��/.��I�O�D�O\�G�EK�+��v�!���۴y���xU�U<rٞ��'�x�w��#���ēN�(#�a���\+��d�t�5ǀ�}��' @���~&�8��/yh���Z�ZnE9����?��O�0�����ɓ9{�x�A��o�@��!�l0C��%�I�R�`1��F�hRp����>��i>Y�II}�@sd|��L�H`k�&���Tg&l���@$���`tY�ꈳB�t�@�
	�a�L�"O$}��lA2>��Ґ,�*�E�q"O�J�B_4G���&^����9�"O@��E@_�F�j%�F�>��[�"O�Pr�+��p��s���*p��x�$�j�'�`�s�:��c�P�*�J��L V�ҙ���'&�'���Y��h��ƕB@�<PF��6
�)���*D�@���N���"���uP��W�,D�,C�V/�D���~ODe�d(D�<��f��D#�t�r�Q��v�Pa�)�<����2c�&��a�3y�,�&�Κj/Q����-�'�� ��#P<P�����D��Xn��Q��'X�'�ֽp$��c��9����#�'��٣F��������U�p��'e�\豁���y�j]�NOȄ��'������V�*l1`�H�V�i�]�Q���S'��5;'�Zy��� �%D��Ą�  ����ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  1  �  G  >)  B4  3?   J  GU  �`  _k  6t  �z  -�  5�  }�  Ҙ  .�  p�  ��  '�  ��  �  ��  ��  J�  ��  ��  '�  j�  ��  ��  !�  v Z �  �# a+ �2  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!�O\e�'C~�kc �<��Q�̥,���'��Ap�՞IpLa��وA��tj�'����T� �Є�Ь�#����'(�� F�M!6�"<r j�"q�lPR�'���EWtl� �g�ʟb>ұi�'�AGF
6�%�V��T����'C�X�%PT�Q��܉��'��xV�U�X����vm
�'oЊ2FE:d@I{���)��)Z	�'8jMQ6��2X�n�"�&V��	�'�h!g���&&��`���c���	�'�L�cp (TP|H����b	x�'Ҩ��W�6�9x ,�Z�DJ��y�Yi�F,�0C�����F,�yB�H�>�����\�8w�ct�O��ybD�/֥Y�`��3F���V��y�BZ0b�$])�' .��p�è̢�yr�\�n^� 2�]<,U�A�w��0�y�O�!Xi㇄��#�ʌ*��@�y�W�3U�!hunP�h��i��I�yҬL	��\�P36B@� A�'���eW�e� ir�c�2T>جC�'����D�gF`ag�}�����'���%%�us�Q��L��a$����'�bX��и8�N��bA�#n&E��'�z5{�?��8GGD�f�B�A
�'��Qr��־5.�A��ȓi�V�	�'{0E�C�Wvj�@s��4=�]��'kp�r]�^����؟�,���'�" J�f�{l.h�k[�7�pЋy��)������)W�]�p{��þ4�"C�I�~X�H�S�^�:%2mP�ca}�C䉅&�`�P�>^K�	�Ek�M��C�� X�,����krZ8�RA=G�PC�ɓ
�*@2���2�-�#K�0a�B�	�o,(�Z�'�7t*�33e\�Z�C��"o��	����r�"��V�O-��C��4t|� i��Й��!P��m��C�	�qib��k�!��1腍*7��C�1�R-r�b��a(VH�	 �C䉭z���Z�'�4"����J��b�C�	�k��R O�?l���X5i\�n�C�ɼPQ�����_�0e�)r���fC�)� 4�2�GLjz Rf�
� 2��@�"Od!1��J�AW��i�6"O�LѢ� P,r�cg-E3v�6��'�ў"~R%f��:qn@�d�H�5�@��y�C 3i ���%Y�E�eE��d0�S�O��ً �\*�QZHQ*F�Ju��'F��ZB�,.n�u�4:�%��y"�'�Ҁ��E�E�H����3"zi��'��>�*O1�剞]&�T��g �Jц%�vc�{F�t��Ft��E���$,���%Ɏ1_���lv}��'U��N�'J��U/�4j�N�"W`�1����
�'�dxR
�i�(1�k�}�L��'�*6�$�O���s�--0� �ޞa�h<Q��'5�	I���,C6��W����:�k"�1Ox��$Ag&l�c�T,�v�§��Z�!�$ČA�
HP��Đ(,�U7韵<�!��2>��!����#Ti��'�1�!�$6=�ڵX$V���{�aY77�!�dǻ;I��YQY�b�<mZ+�-ٱOP6-:,Oޖ�!�����ލ%c|�A����y�	�����C�
%��eZ�$���y�+4n/���C L��P0a�'�y	���j3�ش?]P�bW���y�g�tN
� �iM=g�сǹa�!�DJ�;�� E�*�ʔc��Y�'<!�$ʤ!,� ��Ʊ6��0�.M0$-!�D�x�j�q��Dɘ�	��#|!�E";.�*�lڭ-�|y��FS� !�d� X"x�"��A���,�ve*R
!�$o�ai�����կ��BJB�j1"O]QV���y'J݀d���<��"O�{�c�3B���,�8Ϡ�`"O����(ŵ5T�0r���$�����"O���	��jnX�wI�z�|�bb"O2��B'�"B[l(�c	
��\�"O��I����L�REPeq#�"O"5����=:��9sr۱O��5J�"O�}	������F�9I��t"O��'�Xm�9�@H`�p��"O0�ѕ_�,R��6n���s"O� #vE��4�Z�$����c"O^� �	�"88eQCA?׈��'"O��ز�'D�Q�YYW�:F"O���E��5$
�H��WG2���"O<��hu����EˬNP����y�.�}���;�+�1+@&L��� ��y�B�	w��ʦG��}�]�%���y��C�n�6���(��(�bА�y�,�&�P�����SS���y¨�!O �L��O��J4%(�J�y��R1zO(9��v�l(Rh�0�ybbB=6X��0C��j��T

�y��0���*@o�Yr�	��+Q��y�`]��ʢ��L�T��G��
�y"���(SmQ�A*q��2�y�m-|�m���H�x� [7�y2�O2[�p�����J�����y2��>@��T�Ѡ����K����y$	�v">��1���D$��&��y��J�(y�@
�qib-Y�ۨ�y��i`�i�A��N�9�D���y �����o�5�M)���y�( I��x���P��w� �y�.H�,��83�@y%J��$ �y
� \1p�Ӳ���1xz*���"O��;HS�H��<��%yH @��"O�@x��U^h��F�F�U��c�"O��rV)F�!B��#���[f�q�R"O��$[�pY~e�p`.?�l����'���'"b�'B�'+��'�b�'����f$��'U`�4m|z|�e�I(�?��?	���?Y���?���?A��?a�/����a�Ϗ^6��.Y�?��?9��?y���?Y��?I��?q0����0�.ʳZ�Z<��Z��?���?q��?a���?���?����?�qc[`�R���L�[f�����?���?a���?I��?����?���?��[>
5�����pQW�@�?a��?!���?����?���?��?ae�x[.�pA��`���*�?!��?����?���?����?����?���G�{n�J�CE�@N�T�C��?����?��?����?����?A��?	�AsEsp攞:��H�P
7�F�$�O����O���O��$�O ���OR��Z&~ZHJ��C�/8�ӦJ��f���d�O �d�O��O<�d�O���O����`)�0	�B����1DBA���OP�d�O.�$�O��d�O���O���EW\���"ߕ,��p3�%B;t�@�$�O����O(���Oh���O��d�OT���w���8�HQ0]E4�!iƚ%���O��$�Ol�D�O
��l7�Ӧ��	ßC��+X6v�D%�al5L��'��P�b>�)��f$	�o@��[� .C�@=��G�:�yT�b�4��'�@��?q�D*n�𤨶 �4q��5S�.��?I�3�bs�4���x>!H�����C�pr�5�l��vLV�. b���	Xy�퓃|P<�Api�4<RaPR�;2���H�O��?1���m����$��!Sw��5��b#%�t'����O:��h}��$�<<4�6O��[t� ��a[��VxJLA�1Op�I6�?��D ��|��P��Q\�~U:� HJt�HF�b�,�'<�'��b?����,1Z����kX���G��2���?ѤR���	������� #<�l�	p��"B�2%b� ���ҟ�ە�C�A�c>�Ӆ�'��I�S$�f��[Q��yƎV�O]���'w�	џ"~Γ/N��5e^9L�кB�'!��y�Ac��my�@h���y��\P@��x.��d-Q�U���՟p��͟,xq)J˦�';�	��?�2gQp~I���^.P�����E�r�'��i>e��۟$����h�	.�:(�w��:S�6q)t�L�`i�y�'�,��?����?iO~��A0�ׅH{�h"EN�M�6���P�@�	ɟd&�b>Ux�-_�J�H@�#D�L�(�#kI� �lx�T@�Vy�#�%�����'��	�p���C!,��0CȈ�P6|��$�U}R�'��9c� $���Ba����nB��'+�63�������O��$�O60���^)\��(�v"Z 1�R���(�b#�7�;?A��ޢ�l�SJ���=��\�y]�&��ǊH���{����	O��d:�(��Bhz4n�>>?V��	柜������?�Jܴ��	�5;D/�����D	���H>���?ͧj>ɡ�4����5�C��?��r�'�6��po��6�$���䓴��<�	�K�����
jUV�D�n$z#<!�^���Iȟd��L�Ԫ�='B�"��-��M�3�H���$E}2�'�R�|ʟ�q���<ĖYCg��g_\��	{��@����c�y?�H>1F��90 d�V���El��r���6�?	���?����?�|�.O�m& zȚ�a�)3�J�"*��Dg��ퟜ�	&�M����>��L���S��
 �JG��m�����?y0Ȏ��M��O��	
*}��	����$��C��P�A#Ќd�Iq2	]+F��<q�2����`#
�>��}s �P���RY���I؟���X�'=\��w�2Pj�BЙ$������F>	��'�r�|��4��>x�f8O�����,~Q�i��ý:��0R9O����6�~��|R]�l��ş��@� A�mA�G�dTƚҟt��ߟ���Oy�B�>!���?1��z�bdFǈ!zܹ0bU^����>a���?�H>��� �~��zƈق@����k�C~Ҍ�W4m�W�W���O@6y�ɨ$>RM�R] Q��	؇ls~-r�P���'�R�'�2����l;�EW���=i���-]'�Tp�B�����Oh�EK��4�.j2��S������iZ�|R�3O����On��Z�0 7�&?�����=���S4=Ti���Bb$��� �:ml$A'�������'3�'�R�'�p�����Q`��')T;Ph���[�D9�O��d�O���,�9Ox��\R��ץ�;kz�b���hm���?�����S�'͖h���E�`��3dʰr'X���2�M��Oȝ a��~��|�W�X�@
̼	�Z���'׭c�ڐ�U�U����	韀�	Ο�hy�>��25����*H��RԀ�W#H�8�P囦�$^z}��'oR�'j�x��Q�\���3꙯sy� �7O [�柟�"��y.�4&�u���� �a�A�K@/XZ�?��Q�;O����O���O����O�?Y{PM�m-�����^��d!���`��͟P��O�i�O�4lZg�	�1Z�$	r�H�x���؈A\&c����xybe�!��f���Æˈ�M� H�z{PL�"mW�)xԬ( �'��%���'q��'"�'�	['nʴ|߸�a0�Y�XP��8C�'��\����O���O��D�|�R+H*L������<p�����K~�>�������|z M��J�#k�pT15�Y�x�q��$�"=���<�'?�*�����HV��AtHϱC�B����d����?����?��S�'��$�٦e���E2B�|�6-����t* l�0���l��4��'J�듬?It���*��d'

j�@���T��?���(�J(A޴����� ݩ�O��I#9�rъJ��6Dj��<`����my�'��'�R�'��\>9�c����ha�B:!)��į��D�O��$�O���d[��%FlD1`��
, �{�D�DP�Iğ�$�b>1Y�KLĦ��bۢĠ
�4�Z��q��"\l�Γj��@͵��&�����4�'�z��MM[(�mhf!ԲDzhYq$�'��'"U��ӪO�d�O|�$\�i�=Y�EĳˀP�'.�K*�㟀��O��D�O��OZ��C��9M���S+�iy!Ӏ���ѣ<YG|pnڇ��'p���	˟��G!�������;t����j�ş�	�����PD���'�@��0i�PS�;#�_��̸���'����?��j��&�4說ƘN�`*3kAgV�t��?O���O��V'u�H7�7?APƑ ���d�	�v�G�J�Y�&��^}	$���'2�'��'/"�'OH����ûG���1��&T�l�¢U�`ӪO�$�O�<�ӈ�0jQ��r߄�2���6�ș�O���-�)��q3�<�@�@��0��	ō3*����	��Ԕ'6�p  �Wɟ�|b^����@�:T�,�X��$&��	�L���`�IşX�	͟��jyr��>)�3F6���ձZ�9h��͏kX�ϓ6����D}��'���'�z-�1C	*�-EO�s���K�/>�6���A���/^O�d�����*�b%	)�\���A4]Ғ9O$���ON�D�Or�D�O��?�	����yN=Y@�G�sk���S�Nܟ���П���O�i�O<lI�I��� ��F�+�H�{Ƅ��n��$�������=g�D<m�X~r`��&���iE���?ZPr@Q#�����jߟ��3�|�Z��� �I������� <��˥ �1>W$|�g��ǟ��uy�Ƹ>1��?i���I�f�8�S�Y/��E��I�h��	���D�OT��"��?uq��<F�� ��L D���)������Cܦ]���á�l%�D�0��7�q�
��իƟ(�I���I��b>��'`R6m�<mB~qۥ�P`sh	���� ��D�O�$����?�%X�����ba,M(F����z� �A���HI�Iğ\x�i�Ҧ��'��{��xr*O�AYJ?8���B7�59�@9O�ʓ�?	���?����?�����|W�����5(�.�`�Nų[����';b�'!r��T�'{�7=�IQ0�	;}|H��G2ܬ�Ec�O��b>!����Ҧ�͓/@h]�W뗗r2�i� �IT��~�yi���O���N>y/O���O^PȑcΙ��)�e֞�D����Ox�$�O��$�<ipU���	���ILF.�Q��IK$�K��];{X��?�_�@�	Q�pz��H��|,µ����'8,!XT���XeR-"�����8"��'��)�L	f՚ SD����S4�'���'�R�'��>1�	�-~�X .Y�d��i��("�1�	�����O:�$���y�?�;^�H�d# ��8�V��|�N���?��?�tnȫ�M�O�U����)�rQ�N�`i��Cǘv���`�Ł���O���|���?���?�jU�ТjZ0Zk2�z��^�H�S.O
m�'���'����(��K1�]$��m:@Oًu���'-��'�ɧ�O(��õ��p4 ;�8��� �ȱXӎ�2�Of���T�?�eJ#���<It�Q^���'M�3K���^%�?����?y��?�'����^}��'A�p%Q+����nACy؝[�'�7M$�I:����O��$�O
�2Ϙ�?�r<s��T�pn�=������7�>?i��7Ey��|
�;Y�Pː�ܿ$6�����ɛ_: ��?a���?���?�����O#=s��4r�,���4j��@d�'���'Ԡ��|���~�Ɲ|BKQ�=�D�RA�<{tb�ui�:4��'r���T*�#T;����RgO#;>�i�#�B�FP�� 
>n�ri���O��O2˓�?����?A�� �X�փ���ן=a��(�v
�O����<ɢW������D�I[��	/M��	7�Fj���b�!��D�N}��'�|ʟ6ݒ7邟AА"��<�TY)WK�-n�����eh�~��|Z�Ƿ�%��R���B]$ �e�֛zph�h���Iğ,����b>ٕ'�t7ML~�Z�c&�A�j��asE�}x���O�$����?�]���	�Zn�x�昕@rV9v��}J�������pr)�Ȧ]�'׾Q9���?5���  �D��qƥ
D�n�i�1O�ʓ�?���?1��?����)I�A�~\���Q(l�q`FV��4�'���'�2���'�26=�z)k��#%B}�`�R�W�X���Oz�$5��i��GX�6�y�H����/�290ϟ�e�z�)��t����.�S���\�I@y�O�RGM�PƼ����X�o3
��%��[R�'��'v�	5����O����O��Ҡ�Q]TE[�A�W�P�=�	����OT�D!����mh���U/���XA���2Y��� Ey�W�ݒe��%?-�'�'��5��!��da�T;m��� �\�O�����ݟ��	ៈ�	V�Os"��%h�DTqS�M)<��H&"�Z�H�>���?��i��O�ǎ|����7�(Z���p��>����O����O~�Jh�,�Ӻ{r*D����[F������	g�"�0I�/�*�O.��?���?���?��#D��b3 �|v�@�ڠ���{+O40�'
��'`"���'/����8XY@D�]:����Ǳ>���?9H>�|Z�.޻0uBt�D�CS���I��O�(~�}�Rg�V~�N�*\���I-��'^剡f�08��\	�C�OH4h��ß��I��t�i>}�'����?	����T8`P�B��.Y�ibb�<�?�G�i	�OD��'��Z�t0j�'l���q�Q�!xL,[W��;0�ʼn�O~�l� k���S,<��O�Wʒ�7���3d��P-P�C��ͺ�y"�'��'"�'���Ў�0U�މ�X�x5ɛ7����O����D}rX��Zٴ��jT��c���j�����
i����N>���?ͧ1QDM0�4����P�|���Ɇ+J�cĦM�<�Q��E(�~�|�R���	П������r��,(Jz�4��ސ�t+M�x��EyRm�>����?�����	S�_v�p$V�v�X�t��6�	�����Op�D ��?%K%�v���  �!^H��F�ڲD�A��uc����4��� _�O��Q$�]2"�����?���z���O����O^�D�O1� ʓ7C����RD�`S�{���Q#�yb�'bhӚ��y�O��d���R�1�޻�����(u$vʓv1����4��E�S�����.˓p���2%؎ �,�#���R�̓���Oj���Or���O~��|B��Jb
&�	F�a�v��X�,���Ɵ�I���%?�	"�M�;�RKE�E�d��#��&��8A���?iN>�|2d���MK�'[r=ʰk��-(e�V'�����'�&�� ��ß\2!�|rY��ß�F ���0-6`�h���!x�H@�Iş��IٟЖ'$^ꓳ?���?-u;`��5�<�h�oz�$��?)�_� ��韐$���fꈜ��Y�Ď�Y�8�0(?� ��t�X�A!�A̧u��d��?1t��'Cz�	Q�g2[.�KB%U;�?���?q���?���9���臧�S͐4b�S��6,P��O��'���'�t6�8�i��h��׏���)ը	$����3�y���	}yrgǸk
����DRqjO?��Ģ:Gb��y�Y"(�h|��$��s{Ȅ&�h�'���'��']��'�2�0���|i��à�г	s�J�Z�`�O����O���-���O�|����}Tt��fB�G~%�� �D}��'s��|��$+\@
�Q�N6�&���[2s�^��$�@����շL�
�P��?���O˓)�zp)&��Cp>�%���)����?����?	��|b,O���'Wr/�w���"�)�h0H�������n���,ëO �D+�G�R3U�Z0hT�� ��d�0Ή�0f��o�Z~�EC5'����D�O�g��o	��Cud�7?V�H��ƪ�y��'	�'���'F����u9��c�֑`΀���7c9(�$�Ox��d}�OHniӬ�Ovٳr�W�W9��1h%V�+��7��OV�4�����C{�L�\�܋sD�:�\*���;	�Pxt�
3F��$�%�䓲�4�P���O���ZM&��R-��\��eRI�>xr����O.ʓi����H�I����OS�!qb���>]ʕ"��/H��O��'�2�'�ɧ��Љ��9�p�?C�J�P�J�B ���ʚ�A��6�7?�'l� �	i�I5TGЩ��		Qt��tcиP��7(�I����I��b>�'�07�I�x?��:5$əC�b�)!�>Hh��O����ߦ��?�5W���	�0��[ň� ��p��9u�0���PA�(�Ǧ�ug�����kyriSQQ���A�ռB�m���8�yRU����,�Iş ��џ��O�jM��M�9y8�!� M
G������>����?9���O��7=����n\��a�d�h�b�[/�O&��?���:�6�v�l$ IL�q��G��dÂ�}���\/Ʉ������$�O����9���s���#<4�z��I�����ON���O�ʓ��	hy��'K@��풽_*�*r�D0:�j��DH~}��'�R�|�D� kB����F�~�1Q7A�����S�!-h8x�k�Px��F0@�Ux���bMr�@N�Hƪ��@��=t���O���O��d=�'�?�2�D�pb����f|.�%��?YT�<�'~6M%�i�0$��<�j!
W$��9H�I���m���	��8���V���lr~�`��m](��g�? ���0i] x���	ع>x�x�E(�d�<ͧ�?y���?����?�J�-L�q�&��cƒ�ᅣ<���H}��'��'���y��ѕ;���6��5� x鲣�t,��?�����ŞZ�axWA�5�j�����A��A�q,��M��O2�1�~Ғ|BS�� �GV,���C?)�HP@F�L������Iɟ�@y�I�>1����K�;� )����;R��\�Q�f�dIW}��'$b�'`����,��v��09�+S���} ��	9F������ț'�Q>���!M��xA�]�r���#�TM�,�	˟��IꟄ�Iܟ��	N�������O�R�-��
=������?q�� �i>��	=�MKJ>	�甹I�ёs�ޤ>�8�+F%ژ�䓎?)��|Ru��M��O��IdK�\`e����I���1u��&�����'w�'W�i>��؟�	�Y?�YֆF� �H����,=�n��՟ �'��ꓩ?Q���?�-��Y���	�2np�1D�RM�����p��Of��%�)�HS�"?P�Yp�GZ�iYd��N�X��r���>Gr�/O�iK��?�!�6��P�E�H @�\2-��k �
�{ ���Of���O���<��i���E 5��9q�Ɗ���!�'\B�'Kv6m8�������O.���dԈ��LP�ϵ�e���OB�&t�7�+?��%��Dh���V�V�Q� חgk������9.1�����d�O��$�OR�D�O$�$�|#M�=Rkf�
�×'��"�U)��I�8��럘%?1�I=�Mϻl�F�3r��R�zl�W����H������O!�Z!�iU�dZ!�Yv��/kM B���)��zp���"���O|˓�?y��<TQ�C	K�_J�}���Y8V�H����?Q��?�,O���'/��':�#�NA��"ʠ!6��ҧ���62�O���'���'>�'HL�t�ʬ �����Q�c�0��O8%��w�lah��_�?9��O�M�cA����� �Q�S�*$+�D�O����Oj�$�OΣ}�;3�B$b§S�c��x�$3H�MS��<L�	㟜�ɍ�M��wf�}z�	4%�\Y�L�*b���'9�'���O�R!���� �
X��T�)5�0�KĠ��d�f�3���S���&�藧�d�'�'s��'�xb$A�'X."P"S�j��:�^��9�OB��O���+����p)�#b�y��	3"�-.��O���O��O1�� ��hK�N�=S��B�
�*d�G��^s&6-AlyB!�>��������D�8P�v J���:p�pC� �~S��$�O`�$�O:�4�����ߟ�qD�T1  ى7���L����؟`��4��'�8��?���?�K �G:��F�>K�6m�3�7O���P�4���ΠB��2�O��O��)���B�ԅ�8m�P�c�aݶ�y��'R�'^��'����K �~i�
.eό��ANL���D�O����g}�U��ݴ��7^D�8�-� BR� �oF�Ct��3K>!���?�'_�N�Pش����M�0 Z'nV��A�5�,�2��,
Bf�x�Ily�OIb�'�2i�pc6��cV+F�n��剐U���'�ɛ���<)����	ϼ4o�����K��1�����ɣ����Op��|�2lx��ݱ3�\BM�
��ņs�b!c��$��4��ɣ�-���OhPz"�T@Z܋K�$�p0���O���OJ�d�O1�ʓ��v�/E�LS�F� �<����y��'bJrӊ���ON���u��j�(@6Jf��v�>BxJ�a��	�4��D�=��I��i��u��� P�Y#ļؔ�5z��Γ��D�O����Ox�D�ON�D�|2㦀�)U2��&Ҟ�\���샞+^�I̟��Iퟜ%?��I��M�;'L���&I���!��K�4.R0r���?�I>�|*Vꂵ�M[�'Y>�)�"ؒ}"��k�,�	j�-��',�E�G#�� �0�|bS����П��&iYgq:w��~S�I!�ܟ|�	�����My�¤>1-O�����?�2��U4J�lӑM�75�B�O2��%��.gV��5��R�l��$�Ԛ)}��3��ْ�i�7S�p�O~����O�p���{LBI:�V,���:�,���\���?���?���h����N�<�AG�W.�~��D�]�x����R}��'�r�g�^��]	���W��Wnu��T8"��	����I��|±g�զ�'ۂ� U���?���_��*��ØR*�M��h�3h��')�i>M��ҟ����<�	=UT��AMG�d����@�D�'|��?���?IJ~Γ2VQ�&�3L�i�E	\�?��P�S�`�����%�b>5i4�V�4��F���RG ��,��}lZW~�K��tU�\���䓨�ʸYC$�A�A�l2룃.ܺ���?a���?���|
,O���'Q��k�N�8%ьg)����"R�ouӪ⟴:�O����O��$ھK���P����&�����.���{�e���7�|!+�o�?�'?M��6t�>t����
x�8$������	ן|����\�I���I~���X�#G�W��Tc!�J�/qz�9���?)��
��)�Ǻi�'�X�g;I��<ʐ"�Չ�y��'h�	�_v�o�W~R]�� ����(�,p��qBԂR'R}�Vj�?)��6�į<����?����?a���^���O;]6����C��?������v}��'/��'>��?�����&��@��8AJ�>6s�����֟<��x�)��# �I�~�4#��]�+ӭ>8�Z'�͏`3F����o^ڟ��Q�|�N���� '�i��
+"�2�'���'���T_�x�4�e@�rڲ��'ɃMҹ̓���ݦE�?��W��ɹ[pv:� �����>� �2sg�ٟ���52lR9m�Q~�?�b$�}°�P-<�&D�r��+S�n�#"��<�+ON���O ���O����O��'3������L���h�����<�r^�h�I꟔��Y�s������K���NA���,�:A��P\��?�����ŞL!ʈ��4�ybj�t��)���ܑ������yl��{���ɒ��'��i>��	���Q(d���܉�e��I?V��՟��I�̖'fj��?���?QR�LQNZ��4��8�A����'�"��?����Z�$-y#��;�Դye�'�9�'0�h��ۈ�	J���˛ɟ JT�'�|3$G�w�r�D�A4.��$�'Y��'/b�'��>��I��0��e�*4a�𲶦�3dv4�ɇ����O��RǦM�?�;�R쨡��3L�HR/��UΓ�?����?�F`���M��O�!�DI���㑨m%���eN�o�^U�v�#Q��OX��|*���?����?���K�\4�q�4��E�@��!�~�.O���'Ar�'>"�i�&ZF�<���3̒�Q��9,�d]�'���'�ɧ�O���3��&k��z���G@P0+���4ZE���A!�܄s���<��<A5Ő�}^�8"�!]V���?���?I��?�'���Y}��'NB<�⮌�
� H�G��k7x�`�'��6-!�I�����O����O�4p�`@I�̉U�,�"ؓ��&A�64?��J
<��|����Ђ� �2� )q�0`��0̓�?i���?A���?�(O1��x#$/�G�X�����JN��Hc��OX���O�A�'g�I?�M�O>����;G�&�f�ɮ1[f��f	���䓑?���|
+��M��O�l[�N� -������JZ֚�	dORE���'W�'E�i>M�I�l��44��d �5:T؃eO^)w}��������'����?���?-���mO�B.��p�3I�,�ӝ��Ol��O��O��,y�2�jkE'1��5q�,�Œ�.�8w����3?ͧy�8���'��.�Hk��B�4T��y�����(��?����?��S�'�����o�	Ǌ8���Y��	A�D����ҟd�ݴ��'�f��?��@C)J��$`4��:�ҍ�wE[4�?���d���H�4���ҷ	0	��O��ɅO�f����Ót���yQm��R�~�	hy��'��'��'Q�S>�sJ�	O���2S���R��]�ENV�����O��d�O������X���R�aI�|n2`��@ i�x$Ç��O�d#���F��6�w�h�t��+����H�R-nuq�@~�d���\���"�D�<����?a�`D�+~����� �졖�:�?����?)���d�S}R����*`��;�( �0�[5�W�Cm���b-�>i���' �s%яX^4�uO��1�p}r�O ��ǋؼey��Ҕ-��Y<�?��.�O���g��*w?�˂��'���x��O����O�D�O��}��B���
� 	H�,�EF5����9���_yR�i�����@�
d�%�}���q�X$A>�Iޟx�	蟨����	�'�j�;&$�P���%=C�c�L��k/�q�&������4�D��O���O���3DV�!��#���hs��&'�˓t��I��l��ɟD��A��6�Ԍ��-T��L����5����� �	O�)�&m$H�2�O�	�T�A�<B
P��,_�(�v�'4�`( ���L���|P����B	�a=*���6X���cRi�ڟ$�I֟ �I����{y��>���nu�d���B�Bm�`P�G<P_�d���v��f���f}��' �	��tÕ�P4`^�)��~��щ�"��'��yJ&���?� �����wS�ű�o����$�%Ȁ �'���'x�'k��'��hU�����iQ���kP��f�R�'�R
�>�-O��n�k�	fȢ�zEB�Px&�H7�R29aH�$���I��ӟV��Qmu~���h�dd��A=犱��	�;�$�S m�V?1O>�.O���O����Ot�d��j��QCgG2@Ԙ���O����<�PP�ܗ'7�R>�:2雨_^|�вg��J�D�<?1cU����˟�&��'6���ء I��b�	&�ƦF��Dsso�Pw���kL~�O���I,��'�X��E�^5p �`�YcL	���'}��'B���O$�	�McU�ӕ~���#�m����JVm��<����?��i��O��'LB-��V�A�E�i�� ��FŽz4�ɓ|�X�n�t~� �)Xz��S!J%��58�(J&�^�1�1{d���	cy��'r��'�b�'��Q>�e#��	N�!У ��{��,;<�X�,�	���	n�s�hZ������\�	u�4+Z1��4���Y��d�O��O1� �j�.j�<�)� ���!�
�k�*�?&�"��4O�`�����?122�D�<ͧ�?��(�
*��}�C�W�E���+���?���?����ąd}B�'I"�'M<��wn�1"1$�ٲAۉt:�kp�dMA}r�'��O���1J5�@A���W�c�@ue�������B���d*�e��C�2*���<xEM[F�N�Pr�ˌ̸e�e�]џp��۟���ğXD���'�R9�ؖh��E����d�h��&�'����?���g%���4� ��5��D������:#�ĉ[�=O����O��J���7�0?1�N��v�^��ְZ�t�c'�5d���f��(9��x�M>�.O�I�O��D�O����O|��S�^�(^�h) �k�� В��<�0P� ������K�s�H���L�p���W��e� ��0��d�Oh�)����I0�f~�u�f���3����x����8I'G��w?b-@|��ly"m�D}8��R��%g�x�r�L�]��'��'��Ok�I ���OTث����"v��"�!e�R�)�l�OPIl]��|�I��˟�"�Z�A���8u�����$zP״[�rqm�k~��A	\ը\��pܧΰS�Z2�<���AبN8<�)��<���?���?����?���t��
�����N�"����9j�B�'#�(�>ͧ�?ɣ�i��'Z���R5J�<qt�7�^� �yr�'G�P[ơmZr~�eN�i����ɉ2�2�zB��5���E�����(��|bY�l�Iğ���쟴b�o�#T�9A&�2d��Z�������Ay�h�>���?	����Ζ"|�er��2i�0BB�Ψ=���ON$�'�R�4���I�8	���Չ�]� 囀k�rf�8�@ʎPŮ����<9�'-9H�Dף��k)r��'��9��k�J��/$6����?����?a�Ş���\Ʀ����C?M�X��"�WD(�cCm���	ş`ݴ��'I\��?�
�
[h\���5=�� ��%���dO��6�9?���=P������I��a`#���F�bt�E�{"B��B�<�(���K����3� � ����R�����B�g��L��-GIC3*�ϒ�K
��/����p��*����	-dN*A	��[֙�W���^�ؔ������Yq�s�R��tK$wi�H���s�yQ֬��B��4�W��H�%+٘�B��c�²F8�Џئn1l,���32�;����
װ��p���-�͠����j�f�i!�BB$LŁB&�:9���s��)���tӊ��O��D�O���'���,
�m	GID�:�d�iCCN�4���Qش6�h�1�����Oބ��@�{n$�aR�a�ƭ#������埈��؟��'�b�'���O.��еi�䩳�څIP�7�#�dRk.��'>�����X�I�.ϐ%��P�U����q�Æ
@���4�?�������O���O�Okl�!k$p����6!�}�v���|���2HH�%���������u�)�#DXz}�v��+��u�hy�d�>�*O��d,�d�O��d�1a�4m�rjN'0J]PC�9:�X&k3��O���O䒟<��@ht�����h8iԅ6i�^6��O4��O��O6�$�OP�i�j�� �׋R!��9����,&"�=���>���?��$�OGL�'�?�E�'mѦ��%����6�[-���'�'[��'h�@g�'��� �w���Р�'�hJ�Hm�ӟ��IZy"�'�맶?��?Q,�!x&89P�C�3s���@�̏|4�'f��'!�YF�D�?��j�?�<��= t*���Ad�^˓�?	ey:�'�b�'����>�1�U ��?�0��e&�k���@�i>��'�Hm15�d6�0*11"�d&�qQ��M45�7-�O�l���|�����	1��D�<� �h�F�-Sf	li�fEؾ*�����O���|"���O�m�S�ó%��U�bn ה}3ՠ���%�	���ҟT��O�˓�?��'VFU���o��"2%�����}�͝���'���'�B冓�(�@�o�|� g�z#�7�O�$�W}bR� ��|�i�-���D_��!y�� .���>��9�䓥?���?yI?�rw�Q�Xp	�e�6��s�c{��p�'^��p%� ���`qBF�5���R��Z�'E�@�B,7�b�%�������	m�����ᖏ��WnI�3�N�y�CN#�M�)O���+�d�O���C8T�Iv��i�ό�u���4cԦZF���?���?92���))�S 6����*m���G�_���l�T$������'U�3l*P
 �1�4�x�e��b��<l�ɟ���Fy��'�.�����Ok�17��u�DGĄ`3(]��f^�C��'��	���n�s�֝�A1�E �'F����t �LyF7�<	��eZ�e�~����?���p��Kݬ��eӳ���\�ȩB�d�x��?���w'�Oh��M��iT�A=vx������E�@}��'YB�'�2�'m�)e����%�o���13H�N��	Wf@#<E��X"Q��4FSf�e�O ^��7��O����OL�ĵ<�O��a��QFj�#@V����U6a�&��1�	���O���Or�ِ[�Ȣ�A��/o�@2��i2�'"�	��I ��������F2)"�Uj��,ꔤO<��EU̓�?Y/O��)� ��4�H�8~��d�E�d9�uP��i����D��r��?Q�'�TU�3nՃO��۰�����i�4u�8P�<!���<��OyP�C�%����	J��셹ݴ�?����'R\�xBb��Op�:e^��> �d��1����J<����$�<I.�J�$�1T�謓�m�(מ�3bHR=,�lZM���?�)O`ȕ�x��� V�T�qt�Kp�g�ŷ�M���?I-O��d�k����t�i�)S�)���a	��_;��8k�2˓�?���?�����<��Q�9�p90���ޒ{���'��|�����	֟<��u�L25\�<A�`�:��2ʎ,�MC����/.���Na�s/��0�ޠ� f�\#&�#P�iub�vӰ�$�O ���O\�&���{ͬ����!,��k�� ����ٴ�?A��?	����İ|�']�͉4	e���:�f��i�#dӸ��O���O��$��'�~R�. ��`Wl�b����Q�M���� �s�$�	���I.v`4�p��= ��\��]�¹	�4�?���w0��Yyb�'���ٟ�ثɦ=��)p|�ҥ���7��O|=�1O���?Y���?�*OkL��;�̽��.��d� �:a�̱k)���>	.Ol���<��?���dÒ�3��1�H(g	��z�X��Q�<��?a��?�����q��vV�~�"��SD�K��2�[� �6-�O��D�O����O,˓�?�4�Z�|�i�“����.�R��E1�	П��	ៈ�'yR�~R�� �J�͏,$e۷�31�V�0P�i��T������$�	�����Y���0E]�q�`-0���J�����'j�U�4����i�Ox���O4u���4Zr^,b���"H�b��E}��'	R�'��1�'+�s����?}+��޸<�]C'�D�%?B(lZayR�'�$7��O���OJ��Od}Zw0B�0��	����1�ᅾ>J��0ߴ�?��XA�͓��s���}� ɕ�t�u0d���͉����Q���Mk���?	��?�Q�h�'���0�E�����5|�j���|�ĥSS���'Z������$��,�#�0xv��O�}�Xo�ӟ�������	���$�<����~r�.<*��z䧉#}��Y��
�M�M>�g��<�O��'7��,g+&�����1�ĭ���V5d�7M�O~�dHx}�V�x�	Ty���5 ŷZl�9��P"k���DN����՝$��<)��?���tɝ�
٪!Z��<M��k]���m�7��d�<�����D�O��$�O��pFӅ!~f����Ze�Df_;i1O(���O�D&�i��|���0f>șHq&���5*�K��A�'��_�D�I��d��-g��i��ɗ��F��� �&��*��RnkӰ��O��d�O�m�O�H`Ӥ���O��eB��t7���^X-��ٟP�6�'}��'���$�cg>���Ο ��7z���a��,%��Pyí���M[��?����?�3���'���'���5O�RЊ&*��:`đ�iN2>6��O���?�4eE�|����4���
��.X���P���~�"����M���?��iX�f�'�b�'{��Og��_*|��H�78�ڦ�	�~�P��?!��Y��?�����4�V�OԎar�E1 q�А0�ѭF����4�?�0�i��'���'��d�'I2�'�(1P�R�fm�T�� "d`P�1��d<Xq��<	+O��Ο��jJ8W�&��&�S%w�"���m��Mc��?���?Q�^���'?��O��)�@�w.��K���+���S^���'}��b~�O��'_BD�
x��y�S否w�<(�l���7��Oj��JG}rW�P�IQyb��5�.�
FM�-A0/E�7 |�d�Z����1i�D�O��$�O����O6�Ӻ�'M��2��+7�V�@� <�����ˮO~˓�?I/O|�$�O@���w�1��0zm��;�%���yF���Iҟ0�	�t����m>�1���HI�N��8��<�w�<�X-O�D�<Q��?Q��I��QΓV�d�(D�҉+�f����̶yid�`�[�����t�I��ħ,�S�"�@i���%�H[¼���M�������Oj���O��)��������"�\wu`�jQ��7,WvDmZԟ(�I���I���ٴ�?���?	��<;�%
���h%���*ϵ#�ܠ��i �R��	+.��'��i>7��^��� �DC��
��wM��6ś�[�`�I
�M��?	��?�v]���$]n�&ʕ�PSz9bL��=�6��OF�$ʣ'�D�O����O� r��c�� Bq��*l�,5iڴ�?YA�i��'F��'��t�'T��'�Ș�I�! �b��eFC|m����e�F�au&6�i>c��	)e6�����0&�����.e
�@��4�?!���?��T�	{y��'���[�.��%�Ksֽ���є�Inyb����4�����OT��_��e;ЧՎQn�y�6N�l-�4nZ��4�ɂ�M����?���?��U?���p����'ήXR����ǭt�H�'&Y�O���OL��O|�Ӻ����p`<#lF9V�H$9cK��=خOvʓ�?�(Ot���O����0{�~���cU�NF��#�DŃ-� p"�>OR˓�?9��?AM~B�9�h(�����p�6P���%ߜtHs�i�����|�'��'���ƒ�y��&&��TI�:3\EX#��D�7��OX���O��d�<ͧu�������
� ��#Q��?Du��6JF"'Ƽ�J��iE�Y�<�	ڟ��<���'�~�HX à����эP:��uT��M#��?���?���t#�F�'>��'��5`(5�+�
V��d�Q��8H:6m�O���?�I��|Z���4��6�[# \�0@N��a�n��JP��M�+O���I���	ݟ������O�.��(R~�c��o�l��SkL5O��'mb����y�)�~��O�%[�B��K@q�)�M7�ɲ�4�?iA�iz"�'���'�.Of��ٺa�p��9b>-9Pc�()x��l�)K���	g�`���?�"R#��\"�͊Q
�00�V�'b��'Q��#�	̟$��:J���2R2`񰳥���@��>Y��q̓�?I��?!�k��$t E��KZ;ε�p�>j#���'��'�	��t%��X�R"X ��3o�:���36�u�'}@5C�'��Iß<��������1 �[.��Hg��)k��SW�ixvO��d�OҒO��D�O �A���|� �IG@��̀�@���Dy�'�r�'�OU��9X5�5�[N/��2&A�3����?q����On���Oҝ����O~�ڳ�\�1.q�)��v	��3�L�y}"�'�B�'�����$>��&�"oJ-"	 ��X�Θ��M���䓝?���=h45����ɐp��) �l��8�V��"�KmV6��O���<A�-ډOv��'�����Licv�Q%�-k�m*��>�d�O��ַH��,��?�ȧ���V�ȰQ�%�><	�d|Ӗ˓�?q±i��'�?9�[�I� �>%1D�I� ]�҄(H��7-�O����G��$7��	ф�b\��4K�<mk`/� L1�v�'v7m�O���O��$n�I�X��R�j��e�U�԰v�h1؅��;�M����<	N>�����'Z�9#��ԀV��]Ђn�
a�`�9U�y�����O����O:<�>q��~�R�.UH1�Uf-��ݣfF���M3J>AP	V��O�2�'�ˏ5�rd(7�Up�ҩ��+L�xI27��O&�d�z��?�K>��=q�ҏQ�v�&ŲuLؾ4��q�'	DQI'�'��I�������������ZCLz#�^�+�EJѳi��O���Ob�O��$�O��C�J,\0�����1���ɖG�4�D�<Q��?y����'SX�32�z8/�BaZd�cR���S�p����\'�t���� c�i�G?1-	&FT|W�	=F��t�O}��'X��'|�L�'>!�t�Y|i$8	@�s`�UzV���M���$�<����I=C詺Ү��RӪ��rg���+4!+(�ؑq�*g��9��۸H��b]��q�3�N�	��}k�#[-u-�r6L�2V���vI��e3���6]8�� ��!V�x���^3IE�3�A�p��놚eÒ�s��#0gp8#'N��lo�pz��K2M3X�� �˪G��,���D>
� Pru ��>�\ڵ+�?O&T`� Yi���7=�\��OW9t���P!�9ѓ�̰�L���/-�� �Ta�#���MR3L�@r���D	����	#2��@�fqd��w���hhl5"ɧ?� � �'��~)F�*1���M���?!���O>Lx� �ņ:;2� K�-�g^�b�<2`�%<O���;�6|��瑇x��I&�$�
;�y2n�9�2m�cۓ<��KfD$�1O�	KP�����MBXɉ�d�?�f��'$�e�X,�ȓ(Y(Q�DL69��HGN��D�'�"=E�4�J�f�xU
g��rRxIqU�x�|�Su�g����O`��<���?��Ony;_*D���j`P%˖�[$x9"UM��2`�� �)��<��ˎ30�T@�'ʸ��Uf��nTD�z�(�WX2b3��.��<A�(ϛ *@��,S~9bD)T�[��<��؟F{"��OCP<е.6|�l�J���:!�N�\��5�F
7:� | �R�]~1O���'h�b�@��OB���'A8DI �r��m�э�31N���<���?9�O���iѪ\�8@jj��\#B���v�!���.p���c�-O�d�.��+��x!��E?��CH6bH�8��?a�\��dB
B8��9q�O��d�<1�ˇ�BJ��
��l��;�T̓��=y�ύ�p�h�Cn�$2̐��O<�C�i�ґ"�(Q�[�����NAN�,:�'���8|�=!�On��0���O�eÔ��\��csȅ�����B*�O:�D�����R�W�<�`�ʯO�St�虏J+��+Ĕ@TI��Hٰ��I���I�q������)>G���4�ϒAk��:3���qn�&��T��ş�F�t�'~ڈ�p��&�L�{�gG:��9
�'4���ǹ1�������4��:Ój����A��<~��'C�42���@��C����O��DR1w�i�OF�D�O�[����WAB"���)��[+	*U���>M{��O���1���m�g�	�G���T)ޓh�z�;�a��,��J�b�{��Ʌ8�n82��|rV$(�{6ַ ��UFU�~%b��4*�K�O�I$�c+R�Q�OC�䨢)ɒږ���7D�%S4�U��p�Z/�A�'�"=�O��)� �Ɇ��5���1��G�,v�9��C:�oڟ���񟠔'dR�'��cG*���L�I�R��$ �y�"_�J����d�}l�"@+�r�R�,�6����& �4�Xd�#+�;)�az�o	a�@pr׀�>���ۑp5xɑ��?���i<�^�|�Iay�^��ñjӕc[�P����Y��u���)D���X.���@�ֻ1�!pA
_��M���i�I�Fu���ܴ�?y��X5Z�C�)G%��J�Ǩ)�6�'����I�|�f%�˟'������N�"��UI<j�`�&3O�����E���� @�%'�@�)ܲv��x�G� �?�O>���pJ��!^����AUAD_�<�gJ�r�� ��%�6s�D�G�(�|شH��ܑф%ʮ��0��>����<yKԊ>����'x����'��a�@�s��["iN+�� �'���Ǣ�B�T>�Z�ԁ"V� �VF�d*��(B1� �O��)��Vv�LH�JًxlJ���N��CS��Otb��?�*Tn��-��i&���mR��y D��q3D�}�}㣀6c���Q"+?O�!Gz���>lܨ����B�i�4�AU�AA��6��On�D�OxaX�=����O����<�%V2܈K�gI���m��Lз��'�pݸ�
E�Q;��W:A�V��;2a�=&d�^x�0���ѡh�	�p�ŦWD�k5�Na�|SD��)�3��FC@��)Ї	�v�p8���%�!�$��e��aJF��l�@d蒞��	��HO>a�#���q[��p��5��0�"���.PPߴ�?A��?y)Oh�D�O8擆�I�7�ū �P�3FY`�3�a<�T���̶.�\�E�OVH���ҥ�f	B�	�,���O�@NpM��	Ӓj�����O����T�4�"tjPj	:0�Vb�痀$�!�c��ᲄ��y��SB��1O(�>d�v�'����s2��� �&s�\��4��S�"R���I꟠�'���l�I�x���c��z�k1,�d�����W�Sh�O8�C��	R�,��a�>(J�(��'�.H�����v��1P�G�F�x�e�	&Fl1�ȓy mX2ᑨg9R�����}�輅�`���Nɠa�����RŮ���c�;��'LX)*�C�>�����?��_M�>8@3$|�d�;�`C�?��<�����˰mv�(]���
�^�dT>�	-�?Kά�j˸VJ�Cs�*}��E�������ze�զ�A�O�r�� !n|x1��βGE�H0J��z�'���S��D��ևN�:�aq 	+ ����0D�\�+��P�j��Wh��P��� +OyEzR��0,��
�N�7:�s'?w�6��O ���O���4�L�D�O��Ĳ<9e��/�:	���E:�
,1��Ә'�ԜϓP�v�ǀM.i	�����O;~0�=y �~x�b��T9�A�	RH�V�sBc̓K�V��)�3�ė,bl�0	�b"Q�]��o��U!�,��()�(�dh�ԁ��ɯ�HO>�pdm�BE�8A6"��<}�"�)78])ܴ�?a���?�-O����O���,�d��o29����A�Z�&����:����IA�[�<2tL	�" �ȑ�3��B���Yݚ����PPB Љ�%�.��+f.�O��D�jG�X�F�ǥEL|t����1�!�$ʠШa�C98hP�z�ǅ	1O�0�>Q���+M���'{b�3qzI���E -��HiS+�"Y�P���	���'w:���*A� �_=���1c*aV��` ��>	'l���	�!�`��gO�+��ɣF���Z�iڀl�Bb^4L����ha2�'���'�ֽ�"@���ڑ䍔Zs��2�Z��IT�S�Or��[�m��eV�$ڀ�%~5���	�'�^6MΰC��4h��x,���]:�����<������'A�Y>��ޟ0ˆ`J��Zh�bM-�	H��$����`��@�S��O.�0�	Q�2�I��E�l�<-��>��m�I���Ol:D�.^�M��Y�E�HY>>�L��$�Olb��?!"�V3r�(t�#�8>[0)Se)2D�Ȣd�;YZ�Q�
N(	>0X��/O 4Ez��Ңzc�A�ŀN�-KPP!�
X��y
� T�k f����u� wv��0"O�)x�g�	�\��&1�-��"Of���D�f-бeoC�h��BF"O�Ȫ�O?�ȵ��@E
�JL�`"O��:=��l�FY
w8�-0'"Ofͺ�#��#�l\�f�Ĩ��"ON�BS��p;��I�E�8Mct�0""O*�#���`�r� J���j�"O�3
T��U'aL�\62�va]p�<)��@�a���Q��_�n#:43��F�<1��ƞ*���p� vf���VGF�<��*�	)v"��׃B?J)<xZ@�^E�<U���=� |`b�2��l�b�OE�<�q�Ĭq��1
��ߓ=P� ��A�<YwÁ�e2:��#&�Z�@!��C�<q`�B*F-��1��>���OB�<�����))�����(
)����d�<��jʈP��CmZ~ኰA'�]Z�<I"�H�`�,�)�dT�	�h�hd-@[�<�CwpB1E�6
���8@*�`�<a�c�i.�$�wM]�l*�Õ� [�<!7�N+�YkfMYQ	�T;V��X�<�E�_Du�YS@�;	��6�Y�ȓ^  ����U����#��U�Te��ȓjdY���C3���舤N�D��A�A�vE�F2rI�f��,R���X��@��һ,��!Щ6'�����
��a���+̌�!�-4�l4��s�~)�QE��!��� �tv�$��]�\��V�7����7���Ub�E�ȓY~8l!����]�%��)��W�<H�ȓ1V��Ya�x�`�:2D�4H�y�ȓ0trI����D�:�a��G�]�ȓGZ��3$1=V�S�E�:ƚ���R�>#�(�gW���� H����T�b���E�-�"ɒAEO�g�ل�s	��[��A� Cʍ�M�P3&���p��49��2��X���1\4\�ȓ/3z�0�FV�]4����H�� |��BR��k�%Q	��<��	�.�4�ȓY�4�R��+oN^��",ڶO����ȓ9b�:2敢`�m���Ũ�:��ȓ���V3\ �P���,�6���J��=��O��6���Y�<5�ȓU�}�Q���X��u�Ζ���ȓN^��"4FI+OB��+��3W����5�X�ȑ*�!*` ��%�~�H���I�"M�Oz�lx�&ĝ=t^��s�\�9a�Ot �&S�p����e ���12"OH�p�#`]�Ȓa
�F��T���I�l�X�0���+/
�c���\6��2���L��B䉰j!����G2�B��M�I�z�#K�n�"~�I�n����W�Ƕ��A4�8�XB�}��DA@���2]�a���Q0&l�	 ������'Z���dU�Z,�A(�@,^D��$�H�Ȣ;On)§Pr��c���-��2�"O�c ˌ>LTr�9%��
"�q�r"O�8�k��r4T})ЧW��h�"Om{�#G�=�-!���A(~1a�"O&��!O)�V�# i�*+�0S�"O2���$ � ��1��V,[-�&"OVu�F�
?��i7g�Z�	%D�dAP$[KzT�c��F�M�&�	��.D�`��λo�>��+��i,{��>D�� ��kG�}��qaW�d�0�'I8b�ON�裇VC��D�eNЕiB���"O@9��L�O��܈ n��/O@U��	�JqB�p��I���l#��BՖp��˽Jg!��L�@�@u0�Ǒ�Aʀ��B��eΕPD'Ӹ����DN��Uc@K�H��QP���>?d!�䆎S�<U��HC�s�:����|I��C�z4�p>��
Eb�!�*B�� x��
	E��ӄ����3���P��b���O��r!��ҳx�4jŏ||��j�Z�7��@i�'�Q?�3���4�R�;f��0|�Pix�F#D�|��Ӥ+$ɈaI&e�mGܧp<L�F��s��"�%�1��Z�d�Sl� �8���E��a�����%V42D:|
�	�F�tI�F�)�bD!G�Ӈ@��х��
��	�Xz,��eޗ_X��� ����h4ls����b�(���c_�"ń7`ӝw�@E9$K��Px�%�w�|�!��F�'<�Ki�"������Y(&�eZ�Ǝ�w���4�?iN������:��X��y���I�m1�!��� ����q�Q��h�6C���r�f�h�[��䄀o�$W�p" �i��Y$[ڱ�5-�c�~��ָ�¨$L��u�^�a0�������ß�J$�XS�U8F�Zy)$�گ_������v+��y��Y�4S�L�U�[ўT¤�ͪn�:�,ܶj�|�,|l�	g�z@ڐH�k�t�U+p&��sB
OX�GT$,��˧���_Ă����'�DD�����<����$جIX�O1���%� ���EcT�z&�1D�(b����c>��tI��V�X���e�&��h�4���~��%l���(Hkї>��%0�`�!6��d~�] T��~��T��Gӷp��p�`�Uj��@��;uT�q��H���S����AT��aTOExX��{�+X�h~:���=�ĵ��j%�� %���$.�t<�ӊF�Uv^���)`�xF�N�Nچ	�7�G'��C�	/f�`�V,�'UW�m�E�
j��"�>��fg�RgTQ�č!sװt�)�S��Y�˟G�!!���IޘB䉥��t���i!��0�/�iMtYx��Z�@?|�c~⬓�L'�$%���$�����(���ł�kP�`~������d>��aT`	<z���mT���`b��	����'��^F��eC��<�dE2w��i���(|�z�0�Z�'I��Xd�	##�����0��9[�F�XqVx�Y�j����u�0q�`C�I ��IBh��r9�p�����Eer%0�"<A�fP	�	�	��l:��snY�@ԯf�Y��i�
׺C��!T!B�zP��!���L��F�@*ԌG%�x�H|ӔȐ���q�'<B�'��x �E.SF޽ bB����Ĥ:�O�0`�	=a�i��O�T(+��D�d�1��v
�UI��B�2YJ���n�D�r �,��sr�?�D���!H8�}����9 $�e�W�
{��X6�њN����k��Pj
LUHC�I�<�.���g�>��W��.<�2�kN�|姐���d��̅`�Yl:�����"s�'n�@��U) C䉤r0hQr�4,�������T��I(�W@�A�֧q��S��CX̧q��'r��H 'Z;�����j��p�V=2
�'��Jt�0XϞ�ƌ�2~���-���� ���	 L`(��>mP����i���嬊�{("h��KU">�ax�OT'���AI�*��S��C�]�䆰^���p�#Y�N5Z}� �����D��\Ia{rтrj��fjZf`!q�(���
l4��@��-� XtI^�q_�3}F�j�(���"��s"	��9s"Od�b�J�0��2��=:�R��qOVF.��O>�uW�8L~�;%�t԰�nϚz,0l�$���!A� ��_���9��\i0�ʕ�U�Cz��oZ=��$E�%r<�Ӻ;��L>S�0���4}����� ����Jx8m���^�0>��aӅduj���ݡ+�؜�v���^�^L�hD���Q��'���x�jR� �j$ڳ�2O6P�!JM53i.p����i>����ɧ6��l��K��.��}���S�S�`�Kb�E\�����4�0�F���?1֫ڒI����s�� ����s�K
#=�,��C�{�K$@ڞ~'���'�.�aX>�ݓ?�Xi�GEE�+�JT�I��FB�ɕs�\�c(�Q�`�F	̧�\;��%?Ʌ��K��	ϧC�D�7��H8��(O�4R /"-��dߡ���'{��# ؝�(�� �Е�@�$� ちU9cP��(�"Y!95ID*^�Z�1�����?�F���%��%yv��v�#�E۟�Z��J�'wahS�Pp�\��B�0�7���1P&�~ޱЁB�=~Mq��I=��?a`N֝b�c��E��Z)Ffd��$�'��� Jɼ�R��*9��������:�2�jDL�'�V����'д%���!�bE+�4@+�}��Uh"�T�1m�!���Gy"� ��|��E4(��U�5e��򄏓v�P�$'ۋ3K-���[%+����:�,��)l�T�v���68�4�gԸ-�0����"v�p���J��F��C�
n(�e/'X��5G �T�j陶�T6^)�㭐.�r�C�����0?�/�(U�-����.�[dŁ8>z����k���9�Ɂa�� �kse+�`�>��!��,�Ui_�v�V��v�>y���33 %�mk�/����;�J%�s��R6���vx���e�N�S,T��ə^ٴy��~E�K���q��o[��kFY�D����`ǹY�x�^)|���&0��_&^��umZ��D �#.K/�$D�+K�ј�.^apXxՍ�S/ў8S!�O�JIbh� �t�˅H�UB�ū�,��!ƠJEƞذ<� �S�(�X���T5Q�p"$+B0Mp<��ք��ayB@F�d��X�k�<+�̰(uǒK����ڐn�VC�ɥ3y��`D�ї
|���nDz\�����4���r	*�AV�&Ӹ�'_�aKR�ND�P��vA����6�����	(���э�
l��JE�
�(���']��E
j�`D;TMU0T�\���䅾.纙�r�ʬ0!���f��}�a���+=���˵��R�nI*�g��d���Fcٟ���"��Dx�,��l��æ��,YB`ty_�"?��.
�`�Un�a��˧�X�3k_�����n�+��̆�*���*��B
y�����M��ʭO*��cឰ
~�E��D���Z0�&fP���Qm�9Q��ڳ"O.}�bҏ|�|���].0��kt��^�剳69�QA��u�3��=9�H]RTAD(jFl	fӓ�rC�	#fш�H�	�x�e��>1\ZC�	�}�8� �(Qg��d/j%m�	�')JM��1��M���a(	�'�$H�`�"k�싇���*����'Ѱ����"X���'�8e�'��v\ƌȥ�'Kդ��'�8��ևZ(�Dq��$>�P��'�
���l�=h�&y��8�@
�'>�t�BèP�RCU]�h���'� ��! $e
��CB��U��@j�'H��%gM:{UB�/�H�<i��'���ѧN�/	%A�/8/���'WLт��Ɂ&�$x��(1��IC�'M��K��9w�&��A���\;	�'or��c��j�t-Y���K���a�'�ұr�fO�iiL �Cl���L�2�'��f��duh�1���x���
�'&̐b�Ά�z��m��I ���	�'E'%����AU�Gv�0	�dU��yrT��	Y� K.h��H�-�5�y����:d�)��/�-�Y[Q�yB'�g$h'bQQg�� ��H��y�f� �F���5O��Pd��,�y2 L�&<Bx8���$B}$��C!Ø�y2M�l��`�2��3z�M(�`_��y��P�{b@¡�6Xy����y��J��!:�DC��\���>�y� B����#����p��H;OQ��y��s�ЍpB���k̝sP�M��y�BʔMj$8ufu��Ђ�C;�y� �YN������>��a(w�B��y�NH�4k�Q�`;>	h �F((�yrk��^�x�񮒚<8Xt�E/�+�y2��4\����L�`��N�y��0I���җ$�g�!+��(�yK,~�V��)Z/���y
� d�k �Y��%�K33Z�hc"Ob�y���nm�)g�̉
�(�C�"O0�����x���s��F�8���"OH�c1�5`XH�wG�U�Nu�F"O�DZs���|����	�F���-D���`�X�p���c� �~�X��'-D�`�� ݥ�\�ߦ_�� (��7D�p:D�<#�BPc�ɵ)��,�5!5D��Ɗ,I�`�� ����Y�1D�h���Z�K��ə���Y�� �! <D�� ����0̻���[������/D��Z��A3x��)�ڐ!�.��Sr�<	w�� z`� �ejӨcF pxshq�<A$G؎(p8["
��t
�hh���n�<��e�7�"���M.*0e��b�<9A ��,���NC�P�α�DQf�<�Х�2Y�ܔ�c�M�R�|5�7+�e�<��(�&����d�ٛ:e^Ct'd�<ᄠ�R`���؏U��]c���]�<���1ag���ǁ�GFD`Cs�V�<i� J�&Lfk��z��	��ǈ\�<� �X.D��]�S�_4c�h����O�<���E�y�r<�1͜%M�����t�<I��A*k°-H�mK1I��}�Mp�<�V ����.0Ip�;$c@Q�<A�N
ɡ�-_�V�N�{��L�<� �S�WG�5�Ձ^%,����w�EL�<���8@c�dzs,�#e1z$o�K�<qvl��_BV�{�H�_Y�H���C�<y5��G�(����6�T�����v�<)�MҌiKd��f/F�\��d���Ds�<�u�S�)ٰ�
�E�,!^�ure�F�<���^w�(x��΂%I������L�<��j̗
J��u	�M�xD�oK]�<4\#y΢�Ƀ���L�d5��&�Y�<a�۵uHB1��בo��!
���J�<y���H�t�+sD�K�҉xP'�G�<9� �
�@䡅톊/{Ti�ƄD�<i �ķ9tNP�G�X�JSZ�6�F~�<���T�V�>\�hO��|Y�h	{�<�e�ˡJC6��a�݋ �n@���v�<�MWL����ɇ2��H�CPN�<�-Ո�-k��C�5�.�&�Y^�<A�ѣH���tM-����#�^�<�5�W=Z��;q+Q,!}ȩ@#l@�<I�#�&Og�q�5��jlzm@�d g�<��T�8:�m�A�ƽ)���c��G�<9��R�{�@ �$�X����f(V}�<IrÔw	z�R����E䈵,�z�<iEhц�&���ީ5�Jz�<��C��1��<�̙�X�pH*���~�<1#O��U� QR���c�|@���b��p�>�k�>h�gF�$ 榙��]�<�G�\�T��]B��	bj(���V�'r�?�����/u �E�{
b���)D�0���Q>4�����L��O(D���� �\��7!��p�E	(D����A�hdhx⧆>I"$2�a8D�X!�� Y���P'�ٞ8	,�*�:D������(��e ��'R��e�U�8D�D��H��N��T*S�̋p�p���/8D��c �:�t@�i̓Q���)%6D�0ke�@�h�"`�Ȃ��,	@!�$�-6Զ1�"��#���s4��d!�� ��w��O��l�W�
=^��q"O��"�T�)�E�"�V=Y6���"O4DI"ʌ�Ax�fM\6Lز"O�X��X ��51 ,t,%�7"O�U��%!5���3���j�Q� E{���_?�@!��$I�t��O��)!�D��ۨ�2֥f�dف�N%!�̉(ێ��!�_�4T���-S�p'!���Qe�&��_>2M����K'!�D�d?��Zt�I��m��*N	j!�W���K��1�((�ǍN�dm��'�n�3�:o�v,S�e��Iu�<��'���tc2v�`N�FӚ�9P�(�S��?��K�*��eC��R�10A�z�<!��]�,e��Vd5m�5zwl�t�<���
�:[�8��,�(!�	��jPo�<��d��Gm���iD{1ƠY��S�<���
����" :�\h9��U�<�G�?A��8��
77V��3iCR�<���(<�T�IE����x+��9D����A�0��To�.|L9�DE4D��Q���Z(BS�G?&�X �/D�P(��	��|̱E(9  �H�O��=E��M �t��G�&��b�χ OV!�d�:vJԚD�E]�V��g@G30?!��K����/��B�� i	�};!��ֈeC5��&3�D����U9!�dQ)5"@J�'N�N�buX�346!�ٖ#�h����M�T�H3�Ңp|!�D�7sF�J�&6�`��h���!����E2� �����r�I+h�!�dH�t����m8M�<<G�C�]o!��,C�&�)D��Xkt� �b�-uX!�A[ � $2���CǾsB!�Dɡ�D�	�̐�e$���a��>!�dO8'�T�Bʐ �aSu�J�9!���nFh���ׂ')���W����|��H��&�@ 6.���*I�cM@p��"OJh��B�eW��9�	�<f砍�t"OH�@�l���(�����V,੉G"O�x�� Cu�|�WA�' �AB"Op�C�jZ#��Ȣ2�(~��)��"OY���ܛ[rD"�ˢZ�l�p&"O�@c���c��T�W	�SwƠ��"O,9ˇ��;I�.���)�_lp(�"O�8���@1:���6|W�a�"O��Q@g�]���;��K)39�
�"O�0�eS�E��4p�FJ1�b�"O�E�D��eXt���Ɲ9o�F� w"OV���Z�VF�:�č�3��L"�"OX�Q%+C���͹��Y��� ��'��ي��֙v�D���!f��IS�'�����Dv��	�b���'N�8��#  �j�k5�r����'~&,��Ʉ�{$��Թj�����'϶���%T E��j�hN��a�'BZā0&�}|Q��n�1m�}9�'(*�0 �	��ȃ�k?n���'�F� Ÿ(e��2`(��@
�'��U�,*�j��2�VW�B�(
�'��D��:G6H!b�)z���	�'�8�Zĭ��j����2r�Q��'�4< �
l�6x��=G�>i0�'���q�DA�e��P��M�%7�:]���� �4c�㚕	��0���׃B.Q2"Oڸ�c��m�$P���+���"O$IQ�ѰKi�0����:nm��"OB���	���ڤ'9`U�$�T"O��@p�Y���`��Ѱ/�d�"O�e�`k�+��azFl�#��EA7�Iz�'���܆f=������U���Č^�kW!��G�&��p�f�!L�Vqb$F�<d!�$�d5����;�
��U�>Ea~bZ��VB6GK ��U��az�,(�)�	q���'8�����O"F8��ɑL�t<G|��'2�>�{�ԡS`���c�R�\���*D���ˏ*w��𻓡+jl0 � -D�h�(�a�.iq�m�]�4܁fA0D�${���B� qj��ZN� ��K<�	����^�K~��"� �O��ͅ�^�*6ە��]���@�6���l��~Ҋ�+&�%0���P%��Î*�y��b���p� �dsk���yr��&��3*�NNx�`�`���y��=�ƈR�_J����@��yb,��p�~�"Q�(;��!��g���K���OgZr�B#J�Z����5����'�N`�v�#v�D1;҃	5��p2�'����w/��s��A�~z��A�'1A��X�A���%�V	|���'ޒ��vG�~��� ��r���
�'~��Jw �,~l+��ǃ;�b��	����/Qd������Q�iز�y2��7�z8��F>J�.ݳkբ�y�>P��AW�ӮB�hR�K#�yrϙ�t!�䣖`،
���[�쒡�y���g
l�)W(%�L�	E�+�yb�Y+��	Bƈ�~�,\īK�y	\�sQf��2U�@���# $�y�@�!rl��hF/���Sm���y�֐6v�E����]�ՙA�:�y_�B:�{��
P(�( Q� ��y�ӠI5T���"�EN��⃋�yGB�V`�x��SDj���X�y ��hv��Q"ġ�m�#�y����>k����v�,���W2�y2�_*%y���
.�b��Ĭ�yB�	%R��T�G-����D��=�yR&��E���86NK3K����pO�u�<y����;���x�%)�`�^�<��)F�|%T���\�;�(<(toHo�<!RL�tDZ<)Q�۸$s��RC��<ɲV(��9��O�Lma��f�<1�D� ®q�7���\>Y��0D�t�bэE�֠�m�]��E+�L;D�l�2�ޒ0|P�{ M)�kP�$D�`�qڃ'��@@e���|�hA`��!D��ɳ�u؜��'�B2c:�zՄ*D����AT�}z�Bu�������+D�+��C�b�4*�ҥ!լ��Df=D��93OT�!�p��LS�@`��<D�R��+j�(+��+?x���9D��i�͋;�8���T.��-�s�7D�����M�n}i���x�ط,4D� ��0�ŀ�(�*}�6��"#�C䉜�6�\Y�ޕ�4/ ������'��9ᐮ�AW��1 X���'w"�b#�Q�{@�Sv�� N�&]�	��� 8���	��6|t��8$���;�*O�C�a�  /jp��NG.L=��'�<�1dH'�u�m�8*�:�'/൙so!��1b�	J�4��
�'�
�z�D�B�ƅڢ��+se�'��Y�`�pW@�K���
/��H�	�'��HjD�зR�^4�%
^6!~dl8�'9t�҄b\#���
@# � >���'y$�����]4�Q��\�:��i�'QvY�&��{����7{�v y�'V:� ��YW@bDMBuOxt0
�'��;A�]�O��8j�og����	�'Y��c��@�(	�C�S�UcB])	�'wb��JJA�f��1�ڿO!$�H�'/f����,]�F�2"���NhxE �'�z�`�ݶy�Π�d��\�@A�'���h �K�P�<�S��'k�1!
�'i���5�[�:�3C�	$n��'eް2�kE�?�BL���LB�!`�'�R,�F޾a%N@ۡ��E��݋�'�	{E�*u� ��ɲ-�����'�}���ϲ>�捠 -K)G40��'=���r$��<�]��䊫'�\)�'�B�:�^"6R��7j֜%l����'閔��M��l)�&�y�и	�'lP�D�H�|�Y��Jة�\@j�'G�d��������5�։~t��ʓ9�Z�)ak�)8�aZ�;p�.��4��t��Ҩ<�t5��Q$���F�v%"�/�vf�$�P�گ-�hU��V��|��ǔ�&�h=J�!��6���������Y�N# ���H0BI^��V<�j�F�/1Ŏ$x�%��U�r���d\훲�
h���Aʖ&u|L��Sۖ��,�=4�|2q�] 6�꽅�3V�K3o�$3�rH�׏V�����ȓ#lB�	� !tYvH�O �ȓ_ڑ9rh�cm>aH��DP
0�ȓzb�آ���,D��9xg杀W�`|�ȓx�A	��Y+x����ᒷ&搅ȓW箴[ �ӥ(��T��D�Z`�8�ȓz>���-0>�̠�"CSWF��SK��үҌA� � o]�t�^̈́ȓ@iz�jE�_�8�L,h�
.�j��0 �O�Ij`�;�X�HU�4�ȓM�P�:4/��-�͙��ޟ#���}xfl�W�=TS����h?��ȓ]�l��EԔ3qn��㛁~��D�ȓ&���&$VV�p�<Ypчȓ��pr��U(E���h�f ч�5���j��fn�p:b!A�#�����W��q��B�{�6]"�V�2��ȓ �K"�S/(7<aJ�@C=Q���ȓe���$���N����W;Rfj���c�$ �K�/Q���S��?K��1�ȓ�@�vJ�8M����='"��ȓ'�rM�kJ 0>8֍��kh��ȓ4���aX�;���b��O2)��cbA��I.�j��ՄQ�R)��ȓq�0ٸDo�Iz�HT��-Dw���U6�iի	8��֨vd����W���Rg�D�����r�����E���5�2)�cL�!�R���}���f�& ����G�4=��S�? �0B�Rj8QIˮq7�a2G"O
=S���8�G��z����u"OE�ŧյe�\I�GgB�YA���"O��@�m[+f�����5lβ	�`"O�t٠���L����n�-g�ʑ��"O��� 홈^�r�CGC�R�֗�<i�^<@(��gSIa�y���}�<�k�� �:�\�]I������w�<� �V4T|C�H��d�eMt�< �S.G��هD/&���s�<YըY��hx����v}�ųtJ�c�<9#hմ!d@��/�7��e��c�<��`��v4�Zc��7ِt*�Qb�<�w�)|�`c/�:{O~�9a�]�<a��;y �LH��5g�8�`�Z�<	1�_�|a�F�48�~�{P��~�<aqd�,sl��(�&�NH.��3��w�<ѡ%  J|`Q+�`z�� ׂN�<q�E(��|8lQ�/ F<���
G�<Q�w���1�� aT}5��E�<��+��}��ӆ!Hl�G�}�<�2a�@|�<��%(N�l)U��c�<��%�:�<(���	Y�ąJ�CV�<!UJ�L}��dF=�x�D�h�<3����2qqa�>,�d0r��^e�<�F�#j�0�
:%˲�ɦ�`�<q�&Z�i:�`�ιH�%AH�U�<����o���T"�7vRٰ��U�<�t��$GnB�K��q�*�(���g�<a�d�x�fyxP$&���Q��k�<�Ԭ����qx�e�8cxl����o�<!��F�M����j�>���b�Bm�<�r�Y|!���6b�e�Q*ǀ�d�<Ѥ#��TJ��r�̚(�\�@�MX�<�P)�
E|*�L]k�䙢E
|�<��BX��8��:nZR�ר�z�<� MV	E#���OƵDю��3 �]�<�g"	!&�~%4.0O��r���t�<aAL�
��Y�kM�y�z��t�<�Vb��<�j��	)[��ʑ�Y�<����L>^�@�OG�D��0��.�n�<��J��m�.Q�/��� �<�wmB�"�TM�@�,��X��B�<�1-I:lձ���o�z[5D{�<1UQ�7\�]�%�H�
$����x�<	�-תr`(k#��.'*�D�B��z�<��+�?��ѻ�LJ[����w�<)dC��:]���- ����_�<	�c ^������
Q�Hp'c�Y�<y���>�x���@\D�S��}�<aV��4�ЄXEK#���a�x�<��Mǟ8H�J�	��|���(A(�L�<ـGT�pWT"sc�c 6��	UB�<�H�q!"(cr�E�Þ����d�<��*��[�ƨ {����M�a�<A���^�p`0�Bۗ|T,�S��C�<���Z� ��ٕB�6sA�\}�<�b��k�Ҩ[
����%L�u�<�pkΐ(�h�����;�ⰸwH�s�<�E�M��}(�I�
t�$,Y��N{�<a3@N�S�`Z�­��M���u�<�a,��Y����.:#*�*�F�[�<A%�)xȔc7&@.U�%
K�V�<Y��:1t��yR�51�*uHV��T�<� �	�ӫ[Y ʝ���H�M���4"O�q���'\J�(�HV���xc"O��&䀌bG��M�l�t�؁"O�;�T''il�IӬ�{�ܕYG"O
��J�U�+ʫKWFyBB��M�<��F@)t+�mr�&�&�H�U�<iN\�w�}���� `�̤" �I�<!��:�ͩE�L�XR�B�B�<1ClšI^b�����I�"#l�|��hO�o&��4	Yi�@*K�R��������f��9�=@6ᛃ!k نȓ5���#��/q�x`��n�vцȓ{xzd�&�7k1R��ʚ=����&��s��ܼq.�;�Z�Vu�]��.���!��ςN�.g���)��x�ȓu�Q�ҍT<�(Z�H��)�μ���XȨt�{�`M�qI�D�*<����M�'e�"��*c!ܲ&T��?��/����0��������"P
��ȓa��"����R��i{G�B�
���ȓB��q����+S��J$,�!�^5�ȓu�-z� ��pe�q��S>
9�]�Ik<!C��>��5	�ėw�ұ���c�<���"�2�;dNN$ d���Ri�<�AA�q'�i+T㘃	���YKUc�<���T��y�A�D�Κ<����V�<��J�-;�,����]2��RC�G�<)�IX$�3�bFK$�ɀ"��D�<�,�*�����iљY�R}��F�<9�[�l�v �Q�Mz�`h��Ɵ�D{��)�>�-��) =?zd���o�.��)?��E�U���A� ��44���Y�<�&�*Ssh����G�\��v�}�<����
����M�MsR$Z%EUy�<���#ئien�Y���t�<ɳ�ۍ5�r��PT��{è�sh<9��żVҤ�kӑ*Xh�Q����y��VU�ج)P�C  �u;���)�y"
@�K��LRH#KP� �-ђ�y"��]e@�I��L=B��Z�E��yr��@�2D�1�<Z�`v�ȗ�y�G�^~�s		�E�@�x4HG4�yR+�$KT	��,8���^6��xR��*X~e`��E�%����PFݨD���e�'��ؓe���ĳ�Oԥ��bn4D��86)��4سoD���yS��O�=E��E˹<�<q��N�0(L`��" �Q�!��L;MY�	�v4j�l��硘�M!��'�J0j�EP;���u��b�!�$�yb�I�&����q)��/ў��?�˟\�j A!(lp��Ba��X����"O��I4
ܖ�ƏJ�k�q�r"O�A����4�p��2e[�{٠�Q�6LO��+ec��qx8h+ ����,�S"On�+d+��	o��xd*$�x�"O�p@BʬrJ���b	�<�$�{a"OXs�̔�Q��(dhG�aۘd"O��K�W���c��c�B���"O�%��/�8���VFӭ6���g�'*�䆉1Ӹ�4��cbxX���7SX�'ў�>�rDP���pE�I�u��q۶f3D�h��I/������f����$D����T�9��2wB'g����6D��-W$s����$)DD��gL&D�� i;q ^�rJ�!���x�I�F�|��'wR�B��ؒ9������Bm^h{�'���!+�3e:=*3��8�=�
�'&
D{ ƀs���s���/��Dc�'_�����R8Ɯ�j�/���'U��P.L���$���;{�D��'������� l�$8ʁń_�^�a�'�h�q!)p]nē1�����1�'fx�15'߉~��]ja$�.��)�'��x��Q�i�:�s`ũpX8D��$-� I*��7A�ֵ�SO�'[�8M�"OZ9PQnֈN7�$!tn��2W\TZ�"O,�֡��T#谧*ƕ�z�""OB�[�X���:ӆܑBK����I~>�[�hZ9���N_�L%|p{b�1D� �M�8�D��6^;z���[��)ړ�0<����&j̉�i�rcj�8�nPq�'-B�'�1��I����#Kc���aON���䘃"O�Dj�J�?�T�H���;�a�"O$��O�(B�v�2�9Jń��"OD�[`��$z_J$���:I���"O�m	f�KH��e�g�X�1K���1�'���U~B�)%�<Y+��ǂL1��P�l��y͖�="L��-E�>�hP7�W�y�FP'T`�ISeH�/3��!�� d�B�I+zl0`A`�Zr��h���DB�Ii�h !3gI$b�(��/�y�FB�ɹ������B7>N���t�;Z��D*��D�����)��*�an�
V�>B�ɉ2�bbw F�ivX�+s��*fA�ʓ��O b����	$
�d��}�j�-D�d9��4,��l���'x��+c�,D����o���i¤��}��L+B /D��z�J��6��p@Y*bPzp"wh7D��  By"�	�m�|_�Q��� |O2c��Ga�D���ǁ%k%�)k��>D���"(N3rtV A4G^����@�)D���U.��) ��Gn M�MS��5D��sa�^-�� �2�V����@�l2D�l@s@��5A@(Rf�7:���d+D��s%B�of���Δ�u>��%>D�42�A(�<��!��R�0��h9D�,A�V#h��Q�����}b!�:D�8B
�����3K�le1$�-���'1�)G�7����!E�]AD���G�
_�!�Ć-�L��V�]�\�б�Gf�;I�!��$���C�f�:�� ��8'�!���30}#2��7t<�� �
,�!�Ϟd�(S����Tq<�XѠ��u�!�d�	}yp��J31A��*�@�(jy��)�<�yS��5Q��QoB�u����!�'q����9|��ҋ� �.��?����h��� �")�Y����/�<�)v��d�!�$љ!�d8*`�1�h]�b�q�B��5S$=��
r��С�E��B�I8^Ej��>W���-B�B�I�s��k�T�P�5�J	JtB䉢ABԭ9���&�� ��
ǹPJ�C�ɡD�d�Ą�E���1Gc��a��C�I-�a�g�(SxlH`%��#B�	3\xE���L-nl*�RdX�C��(1M��a�!W_ �IP�m?�C䉈	���� �=4$�Ȁ�M� k�����O�1 P�T(�3wI�ı$��SW���S�? lE��4Pc�I���Z�3�(�S""O���C7KA\�%e�GVN�R�"O����ָ*o�ș�f��@��r�"O:y��KZ�Jx���)M,0QR"Od9��Z|�|ȁkŇ�*�ʂ"O��B'�ΙME�X���!.��2�'�!�$F)ǘH�b�W?5�M����%r�!�Qn�xPNL|D
e������'X�$���#;�@�C�\��C��-hSD#�B��~z�kFk�4��C�Ɍ���Ҡb�n)3 �6?/~B�Ɂ=��!�O�zVT�+A@߉2�C��_n�-C�SĀ鱃�ɏih��OD��$�s��æ����)�JK�Z!��$�&�P�`E+��Y�P$�
~��	O��(��	ц %�&���K�L9@�Q�d$LOj��֮�!!8`��*��^	ܘ�"O���d*FDBxJ"`J9�dj�"ON<:��/YN�{�l\'��d��"O��[�F���#�ӻ���9t�|��)�PoؙR�"F�Kf��ԫ�HyXB�I�*AH���XbM� hJB�IF�D̳eE�+鶸��+�
&:�B��o�0��c�30��x��Ѯ.u�B�ɰqj���B��a�
��6T��AR�Q�0�\U�f�B=Xg�	"O�h�5펏C�h�o�-.&p%�s'�O���f���Sh��w̰���☗	[���$D��P�AL��R���e<�N5yS�!4�<��˅�)�`�Q���a�zDR�|�P�'���
�F�§���5��ɖ��C�C�ie�[��Ɖ���̏)M<S�'k═�,P� ����!HL�Jr��*	��O��B����^��3��;4�n����'�R��((�Q�J�:�k�
�6(�(�N+D���3lʿ3�
e�&�'$/p(`fI)D�0��gۮ
q*��K9VFlI2e'�D.�O(,3�ț�?����� ��X��y�"O`@�q�O�-�pT�
�-1H�5�Q"O��bC�y.!�&"ĚsE�4��"O*q
��îCG� ��.��_M�!�e"On�r� L"@�0v��<elXs�"O�1�r ?_u"�3V■RMnA�"Oh�q`�γ$�}Bw �,X��x�"O�qakM1>T"�V��:e�5"O�т�Tp7`�'�ͪd{2 ��"OFq'%�~�R�S�B��ak�M��"O��(��[�@ z���#I �S��'i�	�J��@�A3)F��tL�t�NC�I�b��mS�at
d'H-��B�	� �Z sSBìC�i���4��B�I�+�n�K��Ն@E�)��g�6t��C�I�V���Q��oŌ��5�j�C�I����0Ī�4��8��+ �zC�ɤq�p*��-$Z1��A��j/R��$�O�J�*�����4�¥J�%$���rW�m*g��N7Q���Y�\�ȓZJ�c�R�
t�Yq��u�F��ȓ#�����ǣ@13�� ����;2PrIW�[0�ڇ�ǍX��ԇȓ׺�0n��u�h �r��	k����ȓx��1�ʄg1.��6GֱM�����`���.Dp�aQ�_̘|�ȓ#3P�q�5�����O��Ʉ�S�? 0I���z>ٚ�٤Y����"Oޤ����Y��ՂgbW9Z4�!"OH��amŅ"����#�"m�~��E"O�S�-�;�`��GZ"#<l{W"O��#�O /+��xP@�"9�)���'�ў"~ʇܘ1V�1[p��m�lJ�e^��yr��c�R����^�v)��J&�yR�2X}&��$�9 �bL�#i��y��ޜS#p�s`����̚we�%�yr���*f��t�M�
�n� G'<�yB��(x���ۆn{����AX���hOq�Nu�!c֥$Gh���l�'�mҒ�|��)��S%�d��>D��Y���n *B�4PsRqa2%Њ+t����˔�V{�C㉼�tq�`�E5	�"�R�D���l$�xG{��- Sz@ ��&!?J��eș�yB��J7��*Ц�c:�)Y eǾ�y�m�{p��'F�_m�I�g�V�y�@]�	��i���jEh�kgiF(���0>��@�+<Xne��Ɉ�s!�$�BȄj�<�BB�*QV9@�,��EQ�G{�<I`#�j�@��!ݾ���H�'	q�<��+��DH4Q�!�Z:�٨Q�j�<����"ƌ�$�4ryf<�v�j�<�E�	� �Q�-f��Z6i�z�<Yd��.XjtjX�{i����z�<�өZ>����$z�t�@x�<i�o�9Y�^�"C&n��Sri�M��@���O&��AVfj����'�����':��yoL�@j�,
�$r%��'�(|;�hޙ]��yA�0md(*�'�i:B(��jT�P���%ː}	�'�f)҅T�(M,1+�NV=φ�S�'�.�9be��O)���4� ���9�
�'���f�ÀC�v8��H":���ϓ�Oxe����0\�r��A�|5 PH��d �S��R�_�:�I��3�6���޿�!��<w�5m��2n:�����!|!�J�򍩳�
/q5�aKfC�o!�kih�0�꓏2&�2�'�oT!�D X�*�r���$&����f�P!�$N�^T���	pؒ��P�C���Dm���w�O[{H�*G22T)�%D��iR΅�B%�2(�V���8a�'D��ks�c4 ]#E"N$\@�¥2D��Zeh�#"S�豠$L&b5ݪ�H2�ON��tv������|S�M�TK�B�8O��tQ9P�~����"&�B䉥v�4<�EZH\"�3O�
G%�B�I<�v��V� ��;5ė�v��B��<�Tb1I�.��7B�$��B�	�
h��	�)zF i5Ɲ��B��/?���)5��R��ȸT��B�I$8���pnށ֌�X5%�B��1q�������I�l�I�h��ۂB�	�HZTͱQHFs�����6	BFB�I� t�x��o��礝�e`��Y���l��'-�.��ҠT%%px5Q`��C�I�E~
�����8�B���\��C�	q���k�EQ�dnh違 ��ZC�y� �X��J�q2x\��պ2O�d5�h�ϙ�Z��؀�#�=N�HY�f�$D��I%਽��   �i��!�D'�S�'p�}iOM�0M��ե
!+�i��S�? �4��JM-]H�A��A����A"O�}�q% >K]aP�e�Š$�"O(X�Q �@����=U�5h"OB	��D� 0]!`�8�.L p"O�m3���S��x�nܦg$��k�"O��C�����P�D���4��=�S�	�Cm40㧯�"-(�����º)ў��i���;s��t|�'��& *B�	
E��aȣl�Z�|	���X&�B�	*x��0�ԁ{t��Z�hW�F�����~��"�a3+!Nt �@ƄVZHF:D���j�?�
��gP �P����6D����4"��I9c��|��D3D���@�/|ܩ��뙪q0�(��/D��b�$2H9K�1"JP�H��'D�ՉB��p��)$p�|)c�'D��W�U�r'~	 ��}�b!I�,�<q����\ Rxˆi��}�۵���N��0?yf� 	󼱂���1/��XS�G�<!��J?��5;A*�,LEh�0z����<Q$@�%5���Pi��0�U8�.�w�<��G9�49s���$(8���EFv�<���FR��<�s��2�;ӎ[n�<�1(�>�HQ�dCQ}�SP�@A�<�iI>�0-ѓ�I�g�p��������`���A!=�\A�m[ ��]�ȓ2��!I�*H��$�K�BA�o;��1R�(pTQ�5���`E�.0=�'�ў�|B�F�(��*B���''^C�<�ӏ�T
�AED��q���YS��f�<�%]�ʜ��Ϟ����	A�\d�<!��ͱ>"	S��1.���ei�Y�<y���^�5*E>�r$nZq�<�B�ʃ��Bc�ZB� -T���ȓ2馉RG+&2\%Pg���u|(��ȓG����E@�7�2p�g�/�|��ȓ
w�|�QD�S�R���h��g���ȓ.b��IsB-r�X�tǃ�z^z4�ȓ1����OQ*,4�eC�O�?1�%�'�a~�À�(Wp���3~,5Q�ꂍ�y2@zAmz�=,��94č0�y"(��XV��`@"\���3��0�yR�U`y�d��H��%� ���C��y�"K�<�ܘ��I�|��"�
�y�I�fF��#����@I��Ϡ�y�N]4G�f���JϦF�f�ʵf��y2	ҙW�pD��
�=?�9�E�y��m~t@�@ݜ�%,���y���F��B4:�	���L�y"lF=Q�$�㐢�"6H��!�`�%�y�C�3���B�� �)�f�s*�,�y���5o"��@�)ũ8���� ��>�,O.��7tήa����L�IW@'D��� ��hLt��J�Z���)D��*�BA.�i`��1	t�8WL&�OP�:�Ă"��fȝxU���}�J��ȓ!���CJ)7�1�3/ċ7V��ȓ�+�cY�nE�e�A�S>�ȓ`mJ��#��ke����f��Ąȓ7��anXF��IsT  �D{B�Ofjl9�KB�d����\��	�'�8LqÄ��
���Ɵ.�9�'j���m d��R���� b��3�'��\���pn����f��E8	��� v�8 �W)��#�$I�d�l�S"O���\	B�ze13��y���B�"OVX[�%��Nt��e�%�ވ*�"O��RG�K),��ڳ�	���ۅ"Otq��L�"N����#	����V"O�q��QT)h��W
0^|�QV"O�A`�Ȏk���c*\�7�x9��"OFq�D�R�5�����'�$�RC7"O��3��,G�����fğZ�¼�0�'���Q2
~�� ���yKx�飤�!򄏨+��!2c@�^8���'U!�ܚ&O���f���_2DL��#�6F!�$�.YgZ@+ژ_R�I�E7N0!�����4"UNϔR�X��Ӷ�!�D����g�8�(���!�DK� �=iBL��S�G�;i���i>�Gx��8K�4�!��[��`
�"�$�hOT���ۃv�(�s��I�~���Ce653!�D�
^�c�FR�n=4��f�ő2!�U��1��,N�=,�F��0!���*EV�w�^A<��ZCD�!�I)8��}J�ƍN(�� Ñ�S!�Dݦ%5��C��	���h! �:!�ț�
�e�;KB���  +�!�I�,X c#j��Cf�hb���&�!���,I0���A�(3`dIDK�a�!�D�5k�&�s`M�z�i��ʔ�^�<���B3�N�H�A��b�F@J��o�<��[�p@t���S�3��y��^k�<�b����5*��K�r)
�ADe�<єC��K���(a���Qh����j�<a�B`h��$�!p;���&Co�<��� ?P��gԔk��Ћ2LZm�<��D�89�H9�4,��f7L�&nh�<!D�U�t��a�u��k��\ѡ�Nf�<���4fZ����ɵC�TX����x�<�V���SL�*Џ�<t�\YU�Pr�<��)'�Y���Z:4L Y��F�<)�-�,f���R1,G;[\P���[�<�'/ť׈ @� _9N>P�A�[�<1�ϭ8�AS�,1��	 ��DW�<نU��>p��b�$C�Yh��VV�<����6J��[��"J`y�k^R�<9Q���FB��C��|�f��fDH�<� K0;����mK�����qFi�<ٷL��h7B�y���
�. �b�z�<a O�r��9J��@�a�����}�<a'������db�Pb��t�<��%�z���f�a��8A)IJ�<�p-�g+�p+f&��m����.�I�<!OĪd��+�i<a6��q1%C�<�H۽p���3�Y;q܀	5�A�<	�iN�p�!/U��yA�@V@�<	��# 8D9aJ��0SNL���E�<�K��r#Le�6���g����U�<��厯�8*�(�{&�qFcP�< �؝YNxi毜,���rd�E�<��ˌ#=�1��g[�r�`5��I�w�<�E��X�YF�?1mru���q�<��醝n���'��K�*<�,��ȓ
��yu�U�fxpG�'�f���BJ��$���1c-ޫ@0م��h ���@�U����o&iwP5��]0r9Ѕ��H��Y�iVD���S�? FA�D��!�d��Dǎ$v��@w"O\*�2�BI�Ff�Lt &"O��r���<���]�T	ʰ�7"Op](��S�zZ\8��L�y�$`��"O�pQ3#�'F���x�F�|1&"O|q׊��2a�g��X�T��"O0YeL�yFzYa�Hv�Y�R"O��04,�5XMD��7N� q�"O�]�t�̉Z����1��j=`t"O� �#
��P��8BF>0���T"Oh蒳/I�U�������Z��"O
�˕aڅv�|��b(��y���"O|L����(	r1y��7m��v"O�8(�҆C���@��J3��H�s"OVM���	W2(2@��3bB�jb"O&�4�!WIF���Q�s�iR"O����L_�Q�s��8kT>�yU"On|{ �]�,k6U+�� &��"O��a�˞ o`��&łb�����"O*<S���b�2�[ NY�2 .�Z�"O�P���V'7V�H�GL�1>d�5"O��s��ѕh�~���\Q�ܹ�"O���4�v�d5�
U�$y��"O�<�������H��Ɇ�$���#"OP��`!If�(�0�X�-Һ)�C"O��P��=��<��Ą&�3�"O4�Se�ۊ5>��3lR��j"O��i�N߳]d�!�i�f��i�"O �i��]��S#��0�"O$��F��a�a3!��0�����"O�# ^�(��W��h�1�"OHh��Վ`\�݁�-B�^*l�'"ONd�""�r0
<�4�8&��U"O0m�3��y�D�`��\
 T��"OVE���+�*�����g���ړ"OF�s򥂄P�0f'�(t2M�"O�8���^�8 D`��f�)�vABu��Q>�K���n"���A��??^Qck(D���r&��8�	����#\�=��<D�x@Pc�	C��0Q�@�"D���9D�L`j.]dl�
��:��Ic�H+D�ԃD�J�X������p���X��)D���6o^�4#c"V=��uR1�&D���"�O0d�� f���E9�*&D���Q!�yV�FF�jpb	�)9D���ǥ>�h9&撛c�by"�*D����@��t���d\��P┯-D�(�VjG�rE �Z�L�|��QN6D�@��E\=������"$:�>D��:�n�'����$(\�7C�q9��=D�x£
9m�5��9 n�)�.)D�Ԛ�N�w������;5I���pL(D��R"kڝv��8����ki^�ے�$D�<� ޤof�{����<�W�"D�h��0M�ʸ���.04�����;D�jg��"X�$$�۴9cj��@j9D��P7�S�FO��F"U2:��}�Ԍ"D�t�@�H�jF�|�)�}�n�ؑ'+D���e�f;��i1 F�Ap����)'D��P�,�;_����F�5`PLydl0D�D8!D�]�,�BS"@ �0"*D�(
� ݘ~�J�ɳM۪pL�H�K$D��җ	D�TL35��4d,�]�g@$D����!O�xD a�?_E<-+��6�Ij���3� 2���-#TC4; �@�0aZ�3'"Ox}�ҡD���*�Jn�J��"OF�V�R"7���� tx�;$"OL1��U1T��4YSK��kʙ�v"O���e`I1,�1����N\�l�"OJvM|4Ψ�3�Ѹky¥�"O�E��f�#X�
�Ǥݯ!c��"O�HP�G9yx��)T���g"O���gH�%b'pK��$mY\@�"O���/�3mz�x[���UG��"O��@�(�sD)a�$EJ���"O^%{%@��-����Ɋ�x�0��"OFd�.ȦL�U�ӮD�	&Tt;s"Od��@>-�.�)KW�=�R�;�"O�r�8,��4��$�Z(@�"O��A�k}����ǅ�x ��y�"O��CU�IL@mJC�Y06بx&"O8c� �W��:Q��iϠ�a"O
�!��"�����X�P���cd"O3�a�y�����K
\�(��0"O��h��X��-ˣ�Ӫ9`�Q��|�)�S�E�e�Ό!=�Z�p&�	\C�I����q/ݭ�J�b�)dHB�	Ld.�4�®e�V$1��|HB�I=k��I["�B�,�J$�U��>�B�I�$D�PQ�
M `ɅH�>/�
B�	*��PQ���
"J�d��S��B�	 �V��p'	(� 1h"c*Q	tC��l��#u��8'���[�k�qVB�	�-��<keB��|��MQ�'ŧ8B�I�]�p�����j��ՠC䉅1�`�sܳs���
WF"<�|C�8��"��|충�A@66s C�ɤh�䭠`�٧y)D���W?J_�C�	�R/��ؤ`~������NW
C�	�Ss22 ��E_j��!�Ц��B䉳ih9�����{�6�d��M�ZC�	!�x�)��V��R������B�	4k�}����"�H��*��~. B�S�>ii# �y��yr&DqK�C�	�)�8��f���ٰ��a�C�I=A$d!I�#4����O�"�C�I�M�� �7]�{$@>C�	�m@��B�����HuܯL��B��tƘ�B��t*��uJZ�g�B��$�x�@�/l���
3x�B�Ʌ-���c%��}2�@f�(�C�	 7�H�҂��Co��b�f<9�B�	�y)�i���[�̣�d�_��㟴G{J?���I%J�d(
��ϡ:�3W�1D�d#��,�E	Ã�)0�Ҙ�`�0D���d�6%�biꔋ�V��sB+D���R�@�,�Z��ת"|�}R�*D���soB�}�&� [2ȝa��:D�����<s��X�
�,rN�-���4D�� B�&�����'G�2����b3D�4@� S���1� ;Hk �#�#3D��P�eM�n��(t�u��G'/D�H��T	1��J�lJ�U,����)D��c��91.0��A-�d̼�8��&D������0m�FY3oǨ1��7�#D� BQ72ɈT��XEwa��"D��!�I�&,y>=��m�$*^��!?D��@�/^5w�4�eꕈ>e{�:D�� �%����IAh��f*�*inXP�"O��8vE_�$(�1�BGu�	B"O"(��X�,(�XS)��h&"O��cH��&-�< hņ%OD���"O�貓*�U���$mH}?�<C�"O̔Sf�6�36Fۋp�����"O0L�%ҭc��Q�w$�?�X!"O�rC�K�B#ҀY悛�'�P��3"Od��Po�")+
� ǁ�YcV�s"O|Y��*�|]�$B ��$8t��R"O�4�tG t�8\��eρf�Lzq"O�0¨f>�C�%�)T��0"O�P�e`OiЊ��
R1��Ň�7u����!�nP��e\JŲЄ�Y8�������Iڰz��y%}��Bؚ�i�!�B��ۓ rp��>m�����	)x�1�Ď&��5�ȓ�B���fT�^IP9au	L4
 �}�ȓ>B� �N�U���ڮ+�d���80T�ve	^fX	�1�H=�H���$�h��&�>%\  E�V�c�:��ȓ}^LX�#��Z}��j�W��a�ȓ<��)�@��4�d���y��>&����)f�@c�-��=�ȓ5�" sj\�M�*t��dH+��T��7���[�jߤ�تa�@�j��Y�ȓd����C��.(�܈���#�Ҩ��yz�����hJ�-j�C֠7blԆ�Q���Jtk�)&	je9e�VX$��ȓ��=�����Y�>�1�a	�o ����ؔ�n������@��i~�l��4����s	 <�Aǆ�����a�N͈Ө�;��ui�P�3r(,��X�|P��L4.[���5�L�h~0��
#��D,�"F��xqS+,S��)�ȓ?X��cC�:m��49��,-4.��ȓy0�԰'@АB�"Qa�K�P��U�ȓ>	`�j��2`Tب�� o�%��l� -�6 �9���1���=tn��ȓq7j��U��#N�D�cK��c|t�ȓ{�4;T�Z�ȃ�ȑ�9
��ȓT��qH�G�u�tL�r�%l ||��r��YsG�Z/[I ��wA�$PfR`��"* ��V�G&�-%w�t�u.+D�p��E´���ɤ"�u_pq�P %D��+w��9\�0�k�B��o(D�h�R�
(H1�&o
U�|���%D�ܨ�"�)RS�yڗe�?r	��$D��cЎ��9
�@b��f�<��q�#D����LD�<Nh�A#)���R?D��֩�e=Xy3�b�z����A!D�DR'&�a�`@�FƶaC�� �� D�|(Ѭē*�LA9�Gà�0E<D��Z�ƍŎ&��YYv�R�;D�D�B�K�AVƋԺOL�$l-D��1n��|�><����`���a�I8D��:�ā1�Pr�,ƮM����*D��:u�C�y�9� �;q=���b/;D�hZ������"�^���:&�.D����Z���jƢ9U,p=Q N"D���$�D�����/�!�����?D��i���T���J��/Ը�@�0D���	K{ lpc�$cz���0D� �Ek��V��B`Nٽ,V �F0D�� Lt�1A�Q�����DY(
**u��"O���T��E�90�$M	�x�q�"O p�uA��@�؉BV�)t�$f"OL��c(2�8����7 ظ�"O��Z���T7�x5��;�4M"O���դW:w1�|��.N)>܆,+Q"O|̛3��.H7��R�P�,C�"O2��A�x�ꉑm��3�)�3"O�Ƀq냅I�@�lڹ${L3�"ONQa��+J9�0b�@R�#:A��"O�=8��G�TEH`��q�|��"O�(�)C�Z� IF!�r㪥�"Ot��Y#s�l�Y2V�,��6"O�������_f|(��@-dH��"O��ۄo����m���ɍ�6�8D��B�؆ Uĝ�qkݹe<��+:D�����M�~�В3��Ks�<D�,�0�͉ir�}��j�~���D5D���6��.6:�鑤���Q�ƪ6D� ��:��IF�B�^�q��5D�x O�4fw����"J�E>0ѡk3D�4pQ ԣ1,0i��[�����`$D���qf��PQ�ĤI>$���,D�PX�L�h��
	"px��M�rO!�d,A��;%#[9�,��7��Z�!�d�.��Y@n�X�p���F�{�!��09:6eB�L#��-a�i��?�!�D�/0L��)&�[ J|ʡ�S"�!��~r�%�)��H�P�;>�!�D,F�V�y�G��Z%�a�R�0!���+_~<�kbd��1��d pb�u!�D�Pcr��ak�&+���� >!�ƦdH�#��NI��ĩ��	�4
!�T>B��}I�R�%C(t�d�܆�!�$K)Zzq�1��&�x3�<:O!�$�i�p���1��@n"!��=�`�EGԧ6�>�aՏ.�!�d�bTL)�E+Z���2=A!�D��@���,�$	o�ԉCc�&"W!�$�5eG,���
Хo�Pq@�Q8DB!�ĬE�Fu�A̴h6h�`T4~�!�׃ ؎h����4��@��cq!�dS -nБ�@["�t`��G�I!�� o�R��-P�e�F�D$Ƭ6�!�D?EU�	�֏&-������P!�[�aZ��Hbo�jD`�YBȖ$j9!�1>*A�B:�ق�݊$!��<Yz�`3���B��BA���!�$��Z���v��{L�b��b<!�>@I���N��.<�T�">�!�D@' �U��H<	9���Nʁc�!�$�=.y:��,��p�:3��$1�!�$��)̥;g�Ӝ?�X �'e��'0!�<K�$Ƞ�D˾)�H�A$O1!��*18���Ɂ$�رa(J��!�䏄�0��v��a�0�y
��!�ĝ)I�(��Y� �W�Y�!��[*����T�D�J�f=�Az�!��M7qD���F��=+������L~!�dαlE(��hz��P�E��!�D��Ne�&@\�@��@ �+q~!�}^�0���%*j*Кaϐ	t!�<i��-:�B83=�-���-lA!���C�.�����Oj����v#!�� 0d��ڱxt�QpÖ�	 1@�"O���$ e#l\i��,��[�"Oz@�����+���;�!��/�8��"O�p@�Dѭq�X��eR:���"O�I;�"��Y{D�	�8�h��c"Ov�����5���͊� 8��"O��
!�0�>xS�̝
p�BP"O���u�� B���%�����g"O� �f&�f!:-��ɘ>`���"O A���_(y��'Y�1V�XV"O���S�#6�&�N� #b�P�'eHѕD�@�SEG	�@�)�'�|} ��,4�0`:�!��s�'� ��B�2�Y���"u�A��'���4�S]9�(2��m6,���'��l���4j�8���ʹ��e;�'�D�xs�5v��਱���

�'�t�z���+3ٞ�hb\�U�"�i	�'"���i�D�!�G��I8	������2�.�єcU.!�P
�"O��i�B�"���#�{��h`5"OR���1E�������|H���2"Ob��d��`�����I�4D��	*O.�(W˄�'$�9s�BW@���'��<���-6��X[� ���a��'�� D��(�"�[r�DpAi�m�<q�e؁��tB�`FWV�ҷ�Cm�<7*B�v`] �� 6`^j�<�㎟4g�`����J��L�<Y�+P:K��a�Íh����A�L�<Y&��	?�tm�p�jo���b��\�<Q�e:	��	[�R�a�n�Y�<Q 䓛ɂP�P�T�R� �a�F�l�<y�J{6��(��=#��w.�@�<Q��T�Sl(����	!��q�%�e�<���NL8{.��M� %3Fh�E�<�R̞�9'�9���-�B�<��e�c4��"E�nƀ��ŔF�<�c�ƋB8NQQ�	T�_l�t:�h�E�<q�K�7Y*�5��Q�J�����[�<i2G�r�V5c��Rl9�9�R��Z�<�I[�G��p���;��5�Ed�W�<�� %���e��z��\H��S�<AD��S=> ؃�Һi��H�ƍF�<i�È��6x�u��3"_H����~�<yP��3|��т&		"^��6O@�<!�mӔI�%iЂD=T*TȓB�<1�^�b���QR��1�$����_�<�TkR.ReҼ;p�C�Q��k�a�<�WC�$jfi��˸{�y�A+�`�<iD@-8�����ͱX0P�S4��Z�<A��Rȝ�����&��T�`��O�<S�q*}X���2v��Ņ�H�<1D��'��K���"�������E�<�r��!�&m+�Q�0~��F.�|�<�22� Lrc*W�9|��$��<a��^��pa�$ڿ1bpL�pb�r�<��
�w�Y��@��@K�I
���r�'��xRǑ�v�4�b�e�6bf�Д�â�0=���B�<81*X�^���+���y�+�e�|�C�*ӫWȎyHu��'�ўb>EIb��4Ȩp��C9�J]8ł8D��u�M�<'�q v�~��8ғ�p<Q�'hGp�&��B�\鱗�Ca�<� L١��]d(���ĳ,�j��!�'E�'��Y��)��=y"U�����'�|�@�(������J�(+&�c��<�S�T��h����r��	�퍂�y�-�*Ĉ"]"{w�9�Q��/�y���\�[��ͬ?h�
��5�yr(.���b#�K�6�Zx���I����#�O$�[C��#9�*I �J�g谲�x�T�(&�1�S��ޕ�i�V�#���@�d�;ΰ?��'.��!&
�7WH͸ �H2�,��MÑ�"~"�K�,Hp���`��a������y"�Y�$�ISd�Uf���%��Ħ<��o�2e�	v��d�>��ȓ0�fJ�+ԡ,�@ZG�b�9�ȓR=�U#o�J���_�(�*�Dzr�'�z��%��K�e�DɏZ,h�	����0�(a�>�f#���(��,�S�O��j�!|��8Y�#i���a��	]����=�Y�Q��U��&������0?!��]B�����6���tl�R�<�ŅՈV�2%���~8l�`pkZX�4��4O06MI�4Q���P�j0LH�G_!򤉺sy�U Y����z�ɑ�J�!�Ē��9�NW4��Y��� �!�DN[Т�0�Ɩ�	�P�B(��9�!�$�?�t[�L&�Lx(TƄ#�!��ηD7�Ԫ��<�.Q1���!���2d�l����daYk�!��<���B���p����]���{��<34dA3l����.Y�r�t(�H;�O��HL�ء�;��M4iW@@�B"O�0w��8��{C�R�AJtLa���R����ЧL���rp͚2#D,ѧ��!�d�� \�q
Q,�L�H�ï�H	�Ic��(���Z2B�
?��1�B�	�y��"OF|�ЫG�K�r ����1ؐ�	B"O&��f�
7�F�r�� ���#"O��2�%%M $�m[�5g"D@C�>!
�老�����gM����`��a���)�S�`����n�(%0�c[�SL"p �n�Yf�B�	�BbV@y��J��+E=$U�xϓ�'1�)Gy"6����`
�>'�m B�ʜaV�4��ɐ��_�*%P�@�4Y�FͺE�*0���8�S�O����c�R�6�ށJ�؞�F���"O0<
���%7f���J>i�~(�U��ٴ�~"�)�#�\5@0��#)+�������Nx��R.OR8k�f ��qgɛ��[R�|"�'6:8P-̩^���VL\�@մᨍ��-������Ģ����x��t���Q��y�^1"�x��&N�+a�Ԝ!�	N%fN"�<y���O���GdP+ � zJ�>
m�(�"Op�Afjڨ��d	ňp����q�'����	�E��}���N�L�
1ؠ�Ԫ!Wx���<扔_<�yr�H޳���`��2G"bB�I�
�m�� Z�a�ޜ��σ�&���,ʓ����ժM�>�fT&�E=<�,݇�Ip�	3,�$�r"�s�`�W,�	(�C�ɦY�Ae�	j��Q�`�e�FC��3y���,�R��)3��%v
�O���$<&�9����Юrm�}�측G�RH�1Q ]��v�q�',D���!�P���p��[�X����?��0|��B?Z������/��:S	f�<a�E�l� rͅ
;"蒠Na�<� ��l�"M���Ag�L����OZ��!&'T�LQ�c���p�'K	\�<Ia@�nm\Ų�e\^�p����W�<�E�I�#$rt���H^xbS�<�A�|�"͸âȒB��U
N��hO1��X"r�F��A+���/�a�3"O(��q�l��d�r���
�¡K�"OH0��̵KU}Y� #��0� "OCq@�%_R��������g"O����]�^�&5B1�A�s���b�"O\Q�W��	TxF�r3d�����!"O�yR�	ִO^P"Q�ǎ_�z)Ɇ�l>��Ԭ�*J2܀T#>D��AbqO%D��k``\%0�Bl�CC��2�|9�f%D�@���iK^�bq���~�2��!D��&�ܬ7��3m�jBB�*D���$q�Ty�֥�3��Ѷ�(D�p�ce�$mE:]s#�?���Ç�!��A��h���R[Xm��MаG�� �?�������GY�V���ژp�Z��t��{�<)w��"�.�0�O)�~[%�[{�<����Z���,� 4���6�B�<��CB�K?ę
P
P?*=�惇{�<�!U�v��H�0�B�<���"s'Ez�<񁍁�j%�Pˇg"Ú��! �z�<���O�����.}��"WMK[<9��eza�?d�$�c�դ0F҉�ȓ�bL�� 6;����p/֜8Ǵȅ�IR�'L��P �i�~pY�EX�e�����'��my���C~��q1'��)G��1�' $yR�H">I]��f�6nL;�'���RI��b`���bЪ�b�'^.I��k�u�.(+#fH%+�ұ����<�Dǘ��S��B3bҚP��[��>����O��Ć�6�|��]e��U;%j��9��4G{ʟ��قL0.x���U敔s�����'�ў(*�m�~��K!dޕ<,��U&�pyR�|ʟ��(A���C6�5*>�4r��*D��0��Ku Z�C�apL��,��p���';�\���_�(��8�`
C}�=Y�'zvY�C�	\��؉��I�=�~t��'(�8B �5s�V�+iT�.X�X�'w�y9dƆ� 7@p@���s��M��'����t��2\X�Hx�������D-lOF�h�i��i����Ο/Y��)q�i�ў�}�ڴ1?\Y��˟."H�ڶ�	+�dl��O���Reb�F�DX�P	��ȓD��3,6b�H�f(��3Z���22h���3}�P`�sj���L���
>x�1AAg�����ϮuUHl��Cb��s
��ux
 &�h�~t�ȓU>�$�$�T6%[ �s���]�@L�ȓ�^5�p*�!(��rGJ�1p.i��m��%�V��t�H�Z0)Ҡx���Q0���H��j�aaәq�\U�ȓR�*3h��1��T�.\��܄�k����),X%rI���ǌ�挄ȓ3̝��oCp �5�^	E�=�����+Q+ʞ	P*@8��F����tL(+�((�P�)��_�%�ȓ��IS�)E)��ȸ�M�Q��ȓ>z:=i��ޔ#> '�ð�����Q�)���$RD�sө��r̄ȓ*B`���	�t���X"��y��S�? Ni@���)�҅С���kt��3"O��G��%{d�jrJPt���"O�t3Di�"���e���A��i3"O�b�dY*a}��X&�'/�b�"O��9!hZ��4딡Qd��"OT��%ۛ��A�ނr	���6"O@���x�m��F�$��4��"O��zrj�L����d�N�BV"O�u��ܵ=;0��R�N���Q��"O p�'a�f~fTAt	��FL����"O9YqEY)O��a��O,����e"O�mP�)en� �A�-g�J�kw"Od�ae�$ڼ��D N,N���"O�;�.�&%�T̑D��� ��YYS"O�̂@	�<e|v%j�ɍ'����1"O P��MG�<�=H����m��e��"Oh�i`��y�5
��O�����"O.t)rI�i���z��|�h��"O���L��.�Cq��z@@�"O�u�'IS�"�zQ6���*k�t(6"O��q"**,�
4�e`�5EcN�R�"O�ʛ*,J��A��A7��"O`�6J��%8V.�����4"ObQ�U�ZJh���+9���1"O�y��n�)f7J�`!��#>��x"OL��Q�]�7���#wlǄJy�Y�U"O8 cg��`�'KE�FtD�(�"O���X�Z�	
7kQ�p��É�ޞ���Q#w�����'�h�*��G�{
�,z��M(2�0�	�'@����I�h�tH�t"
5Y-��j�'ۆ�r�G�X0P=1�ČY�d�'��(s�G��qCGM[ۮ���'
��s��kU�5��(]5HTtA�	�'[��z�BJ8�i�t�N.G��H
�'��	s#��(	�ĭJ�� fN<(	�'��F� V���� ��&�*�''h��v�]�<(�LCC�گ��T��'}�q�o{�&�[�kǽ��<��'���&�)d�i��FL'
�H�'h��b ��;�8h��H(�؈�'�&��FI�6p��I�c�
��d1�'>��k!�:��ͫcNF� պ��	�'�Mk�g��8��kc/�V� 	�'
ȸeYsp9���Y�{��r�'�d�E5�FdY�e�,iu��'A�+��4drq��ΚjΞdH�'�ꐰ2�W�#5u0��K�nr��'h�DCHC�D�$@ c��J�'_d)�/
�XK��U�g�D��'���S�Wa�x���� 5\D��'�H�Kɐoy$�C�Y"h�,�*�'P}q���\�@��jU
���'�b�&�ãSD�)��[/s��\��'W�I�É�[*���C�B�З�y2��g}ַp�B�)y,-��¯�yҤ�(A��)f�X�!o�<��+���y2K�0�h����P
S�"<"V픣�y�Y�!F�T��Cp��B�B�=�yۖ)�B|
�C_ X۔�(�y�lӃ�dp���/i�vz����y�d?`T���3��7�D��f���y�E�#~,��"N+{�efB��y�#\�=c���d��phʖ-��yb'�#��[�O��	H��*�E��y
� �pCRϚ=M�]�' R&l���I"O5�D!]�}1��83�
� q҅b"OfdPB�/�0ጘ�ei��X�"Of0˂���B%��RvM�BF5�"Ob�kr͆+R�6fl�	����"Ot��B.ݝsx��$j��dx��"O��;@
T�6P!bJIm�*���"O4�9��=gV	����g�N��"O�	��@_�E�<P�s&�5�̍!%"O.Qh�C,βqj���]��� �"O�Hj��EQ��H�R�b����"O�r���]�R<�"���1�dA�Q"O����7(5Rr���T����"Od0㒠V�V"9�eMT7(��%�"O>�"�Ԏ��W+�z�(�#�"O�3��9i��	�)�"��q"O�E�����B"����V<�D�A"O��`ƫ�fK�)���B�p��P�s"O$��'��=@�^�P��%"�h��"O��jQ� 4��C��C�_�u�g"Oti�G��<s��5 �b� e�R9�E"O����@�)O�����>l����"O�P
���8�]qS���M��44"O��R�?#��k�H�(w�=K�"O�Pҷ"��M�q	�=2kB�q"O"q�uN�6t~8�bS�aFBxs�"Oj1�r���(D�X�D�G�AM��"O� ��̍�1&x��U�՛
+:�d"OR$s�`3,	3s@�m/H�*�"O����� ��g��"a�%Y�"Oaȧ�ιr���VB_�k�2m�V�xr��>��a�=�~zAF �W�ȼ"U ��~��K4K�W�<�*&p��##�����l��&�(/���'DM�&c��ИϘ'i>�ò@���Պ��Y�7V��3
��rG�p�ǥU�$<��)cD�>6�`���D�&�R�h�c��3GV����v���bf�L��yt��5�Q��{W�N�+c�1��LF��Oɘ��HM;zm�6��'s]���ٟ\��➈E��'��9W����TP�6����[�'=�(�BB6B�����jq�?��NQ&G�p9�]%>)(�Gx��!�B,e������_�t�� �ʇl�p����H��U,�b�pж�G	W���?Q���;��s�	t� F��x��Y#��,�n�:e,<�OR�F��1V'���7i�8j��E D�v���Iq�y�F�����@��PI��}�ɹ�����Ҟ~*�eF�J��8@랗� �ڐ�G�'�l�qH07���GE@�C�:8�aL��%�#b �rmpE���b7�����Q�=.RM)p[���Bf�F�g�$L�i�HT!�7"������}"�D�d.]sB�؛4��G!͆l�XL#�)جE����E�2xH�)CJN0Z�j�ȑ�VL ��4�O@��? ܐPc7	�0|�z���i��g��c-�5v�� ���l���7'��abC�!]4�EΓ���7�]g��d���X��P���Y��L�0� �@,H�@O S �{�{#��{4B���Z0`5�: ����⋸C%\��'�`�#�?q�EG�S%&2'D��Fk60
�D>ړy~��D���O��=1,Й���g�WL�.y�$\�iT��Y7�'6�y�dI�HD�M�.O�rD�I�q��^+�9�#m�7�(�c��R�����#8��e��ʃ9 !(�q���Z!��C͟6
�*b>1�d �#v���ISV:�Y���J �	k�'Yc���� zY~|j��� r�Pk6D�7��!��%&>�Q2gI6cH�)�~�&d��m��O�D(�	W 2y;�l�)Kk	Iz��XM(qS��ޠT�Z�xD*��@$����ϝ5��-rEE���H��ɜ�M�N>1�ȅ;X��ϧ*$���ҩ'�`�j�14��F|B Eu��]zuD�hR���_Lx'c����Pk��Kw8� o�P:,��{���(���D|rE�*I���sdF]&G,4�ڕID��~"�"1�>!Z�aU�O'����U�Z_�	bӎç6���c�ʃ�y瀹� e*vT�-�ȓJ�J���A@�)�X�r扂kF��ɔ(��bI�b�4�6�Q^�I�Z�(y�O@�b�͓-��[��0:�m���a����iZ��Y�L\M0ON4K��"ԇ�����䕴��td�-AyL���	�\ה�k��u���f�"Mf�աÓe�}k��Z6�7�ݝHIf���  Q�u�ٱ8���c��&�b�S�RZ�!���.g��u:�l��#��p�.^�P���,NC@)��|?yFJ&A�nq2���^ext�Q��]ڜ��٦�y���?{��K����|�u��;X�	�-�h�˴h[����%?�ۤ�x��Q��V�{�b�*�X��v����?y�Q� ������(th�F�*6�~��������!G ��rǑ-R@tX�$�W�џ�d��A�\�A��d!9V�J!K� �i�,��f���y"�P8'���{���yd���~�)O�I�2gP�%�D��M��|�q%����s�ҝ&�@��V�O�<���o��d�$�6@����ϗ�
�l3�p�C����g�E�d1��"}c<���^�����	(G�L�`��A^"Œ��*'��|�s*L�	�C\a�azwp�p�e�8��e	�\���O����#�:y�肷eؘs�\�%1\䬔�1ݶ ��H+z��C�	��:daW�Y"|��d�7*�2k���ӂ��N�N�RF�R��}���	�>����P�x�j5#��Y�!�Dɒ\�"h�Fػ�@1*)�3-��8��B7Oe���I�c��1����|���0Kz8���;T'OH<�y�C���2�a�8q1�O].�?Q���(f��SG1lO�)"2f�6sA�ر�f
/�lh�4�'m�l��L��O�!n�?%�z�[2��9EG�-h�� v�,B䉄U�j��kB0a�t5:� :	Wx⟈iW���&��'�ӑ1���3%+�"z0�x� ��I�0B�	���@#��?��<�bG�n��pi7D$���K��G��'|��� K�}��9bCG�T�!@
�'�&D8���
K�hq &B�1{��Ī�����d�a&����R�n�8#E�K�� $�{2!���B���b"�ΠM8�-s��D5�x:��$D�( f@�T�e#
k���҄.1Y��1zL ��h�����/&��y$E\�hZ�	u"O
����:�x� �2�b��a��k[h��C���O��  O�?-��T�ٹJ>y��"OlP�aU�Q�`D�㒻2A�=(�"O�q)���V�DAXGW�}"@"O���'�R�>�� �lE8���"O
 �A%���/�.e!:|K�"O\�Bf
�YF��2��A�6"O�ؒ����l��)��Ѱ"O��ӦC��S��P3흧#�p3v"OZ��L�J��4ٓl�}�P}h�"O����'���:A��1i��{B"O@�y�`D�e�Ā�+ql�@p�"O����aϊbR��r)�U��:"OрԠC1{��聎�
^���"OV@��w>\�� �.(#�"O�MY�%�V�hz���A�bEaF"O~��b?QF���MT�z&�S"O����oC.AK�;��̲6h ;&"O�S��E6x�Pl3�]7'c�h۵"O�p��EN�n�`T�`��%XxY�B"O�cR��d���a6�.A��M�r"O��H���Fʍr�bÔk�-pF"O�&��`��|�p�B�rU�c"O2A2g�R�adByY�	�rՂ�"O�];�ڿG*��$�g�.}�"O�e�C�J;| ��c�9�lE)D"OV���;�BX��bSs�(�0�"O樨!Jڣ�&|�6t�K�"O.A�5$�P����F5}�y��"O�͡%c\�/�R�q����})�k�"O����(�0cٌ$�`C���X�"O���S�]=�~ٱF���]��"O��h�a��f���� -�.5	�i3"O� �]�n��<8�9��ܳx�)Y�"O���kL/�4���9f��u�u"O���E�G{(`#W��; �te��"O�ePӃ�&PF��Pp�_�h��=�Q"On��Wf�+3��җ�G�Fiz|�'"O��f!�c\�����E<8��"Ox]!�f-�T9{4%�� j��@"O��Q�$��!H���B�H(1o�q"O��sd��:O���Q`I�HF�J�"O(���N�s�*b�c�D7����"Of]���z��+�a��%HL"O�AȲ.��:���Ô��%l@�)r�"OH)�U���c�����%4f}�Q"O�!I4�>L����PA�6#X)��"Od�@��:E{�Q��ڟ��41W"OՑ��@�~��̈$aA+e蠬�#"O�Q���$fx�HT�I?H���"O\�:���;7b�Ԛ�Ҷk74Mk�']R�0#C�7�^(�� �L��3	�'}����>m4�H8�U�	r�-#�'E<襇P,Nl\�э�S�)C�'�8�	�6���/O�2x��'nNd��N�,���9�ƶP��(��'h�2��e&�g�?#�i�
�'���@���Ƹ��o�&C2�`	�'�Pa�A�7i-���U��o����'� 1�j�MO�*�/Xe�R��'j��W���(4��#��]�Be��'�� A�;S��Q��*PX�	�'+��ҬH!f�����O��t��'*�%���P�"j���$	�:���'�Ę"efJ1��@�ï�,FT����'o���$�Sy��I�q�:�ʡ8�'V�]�q�Ɗ#�E@�"�,jdu��'�`5r��9M�<P�)��~{�'��ѣ@��r������'�h9�4.�lP~�z�K,e�z�R�'�D�Q�ϥ;k�Y�V)��[Rd�'��J׆Q=H�|4�'+ľ[���@�'B�I2�H[�?�"�R�O�Rx@$A�'K�|(#��\<����JǠ?���P�'�0U�!��	����
N�6��� 	�'�|%�E撣ϖ�(3B�*"�����'<���ɏ<,����sK�tS�'I�p�BΙ�]1�d��m�`j�'脑��C�8�I�$�-[!�u��'3j��ҪK���P��K+B�b-[�'�xš�kX� ���՗1����'��X�p �!\�%��f@L�!�'��g�m�@���C� i�����'(^!�2$\�
���pgh���'Ӻ�k�b�W��Z@��m�YR�'�|�`%���.�0��W��u�l:�'�*�"$��Ze��Lal6��'��u���69�V�I����Pd���'��y���Y�"��H�G	L��u�	�'�<Xs�#I'?�1s��Ԇ1�4���'"�m��#�)�%N69��'�(���۔d؁���(���#�'e�@��	D+/,r1���1�]s�'����E��yH��	�DLB�'3�h����&Zsr	�D��1��'��E�#�(7,D!Bf��+U����'��@�E;�|�4�W�r̠��� ��h6�S�7j���Ȋ29�u{�"O`a�O�1��S!���&����"Oh�Z0�7r�Ny�7��!N�	�A"O8��T��	"����R+��V:V5��"O��dD	A�6<�ë�;*>h �"Or<�%ʤX��I�����"Od͙�l�QA��BF�I?O<	��"O����<?��M;�I�6o*�hb"O@X	��[�-�yRDg�^�� "O~yv!"���+��B=k0 ��y��˸th�[r�^'|���7�(�yb�,(���Ir�x�{ L��yRÖ1pئ(Da��0��[��y�)���DA�N�n��X�V�.�y"@�
'*e�a�FphQ�����y�*�:=.)S�)W�q��jGW��yB.�tt|�5ؖ~���2��6�y�o� �@P���Ѥxb,lJ����y��V�.�H��S�t(�1��yR�K$b�>drVoتp1��*ӁҞ�y��{v:�Zj�B�@S�yB�P�-�Nab����i��xԉQ�y���7
6%A�Z�a�`#�!˺�y��DS��4��?�l���Aڲ�y�E00uj-�	��e���y�͇�l��yg
A*��Y�Bʎ��y�&�K��Z�h�9y�>Ik�#��yr�؟ ˾XŋO;
Q�Idlű�y� A�y�4�x&�!aZ�@��yR�
F�$h�3�������!�y��H;�}�V�
�(�7FQ�y�/ϮSED@��	�6T���
�y�� )ᄽ�w�tA���_��y�L��ZWK
 �m�����J���� �@���c �͂wM�����ȓd���`�C�>iR�
��c; ��ȓ>`��u'2I�>@�@�
$M 0 ��H�n!��X�u�8�[�ü����^:j`@⩄�0ݔ�#�ǹ""�1��@4���L*Sj���C�2ytp�ȓ3b`m @
�RU>5� "R���(FV�qOl�}��<�����cR�4+��
;`:�(�ȓ@���7 ["[��l)�ӯd��$mڼ�pc$KX8��3�R�[�l����݄�F��c �8"m,ݩՉF;��IR�	�tD�"���y����d�a��l�P-2%�3�y�FD�V�:X��-�'��-�><m�R���1g�����@P�"`H���O�A!K?��	�$������ �1���Y2�%\O�i��(.~�X�ʌ�\q�l�)F*�"�wKG�ֆ���G�lб*O4P3`7�3}�oU,�lB�n�m�#�G���'܉��T{IL�"A�b�'T��0Ä�_|�����ԚB���AJ1I2�i�aGڛ�0>9 (�)�����e�:a�L����ڄ�J���KK�_|��}�(ʧ:��2�L�*9�U��'�@�!A˞_NJ�xG(��Y��'��\X"tY"�K6���4H)j�&�&(7���c\�՘���'��Xp*O�e���'*�M� ��3��܇>ᰘH��M��$��N;**Ӈ��' b����-a&*�Kv�Ub�d���G�5k��vR�h�a_��q��X-
���m]���k�߹+���=a�/�Y�D�:���oΚ�*E��O�78�mh���r�}��X�KOZDI�\�3�`�`1�'��$ѓʃM,��C�.*A��i��
��>�2餢X�'�x�l���i��c螴����0���@NZ���`�Y&'z��R��g�!򄜦|���C��ũ��� -����7CP
i
2���<��� ش��g{>UsQ���|*��Mm�����N�/H�r�jB�^����djר'��yC,L�"�I�0���� T&:p`��M�"����	�g��t���߾P�ܵ��T�o �U�/�*M��k�M܉]tNc>��2��#@��2IDE���/'D�� "m�E�b��y�"������'�O�(�E�0���M��}�S��a�P4�ʼF��]�G�O[�<�֌:{7�d Áz��i��Q_�D� �уbA��0<�#gL�m��h���������L8�K`�݂#��d�v�1���~{�I"��I�����B�&���'H"�F�
�2�1�)�ΠA�O�mh3B����O�#�)�r��>���'�
2�Ւ����T�)b�<D���w�Oi3�A4��'��$�.�~���x�<��H�%j��O�8$�̐�(+�HQ��l�����ҁ�-�O�ܠdhGx��\�MY���)�A�!���2�&�O��R��p;���%|:z��W���&X��(�J�5]��Olf�T/$]�9{c���r
�'�ԐA��@z�0r�Գ_���)O�aC	�U�Xh�K��|bh�>�����X���rsOLJ�<�h	\Tx���υ�X]�t��B��
�n��Di���gܓKo^<��LD-5����]�,��	�IiN�C�لX��Qt����ڧē9��U�%�'�,�R�Q+i4N5�GcѺP������)E��� ���E�F]S,f>���&PV�PA���%�\�!G�#D��U��0uU��x�����,5���#?�ъ�<�Qb ���B�����PR@�3_��H�h�m !�D@�~`S$&N59��Y�c�[� �;q�7Fg�P�ɕ;T�M ���|Rd4iO�u�`��G�aa�@Q+�y�I�p���G88���R��?�$ɗ�l�l��30lOF����k�f�`P(��MĬ��'��U�t��I�L�l�5��H�G'�5e(����d�^C��7�RX¶j��4P�S,go�t���L!h.ڹ���=��İ�4N;��㚠m�C�<FL���q��M�@%M����[d�?�u�L��E��'�e���O����'��֝�
�'�μ�d�����A"t�@�t�����Ib�	�k&AS���*M|�y��E7L됐��O�A�{�NI,�� ��Sꦉb��ӉM�0ܛ�h�24�S�f0D���S���#^*0�A��^�f*�A�DTq'���h�Lpx���?n[\B*�-,|��"OFm��
�2�(a�I�&f�A�Bc�69�d!3����O�h��I�c�H�Ҋˀz���Y""O`��&���x�*&�T�Vx�"O���0GEK�p�R�M�Nנ-��"O�����ʴ*�qaJW%L���"O\��d�׼D�ܠ+�Ύ�]x����"O�ѰV�N����z�LàGl�4c"OX\�a�K ��A�P G�c\J���"Ov����\(O��u�SnB�Ŋ�"O���f �	0Ȑ7�;PB�t��"ODx� ��G� 9B��(3�@q�d"OHi(��T��H8X��J$h�L('"O�ձ�����@��X��PE�"O�4�� ,�����(����&"O&�J%�@ E@IY��$��"O��#	�w����Dq�n#�"O����ߡ|u�`�t�G<`��y�"O�DH��##q�V�8a*�{p"O�h�ԋ��(�,��Di�wEh Z�"O2�Auā�AC @Z��B�Q0(�T"O�ř�ߙ.��K�� �:JT"O�\`b�rE<!A*̞Q�t iQ"O�@ȵ^�.5z��&&k�>tkC"O(2��X�tq�H�jx���"O��6^*��d/ڵV����@M��y�K��KN����.K����6lW�y2Ø�s�f���'8s�ʹ�pfH�y��K�E�nH;�ɚ�Z�Ys�J8�yҍ�17�x�C��[(�1�b��;�y
� ��{�a�=%H�hI̠Y+�i�"OZl �Z�!-:P�h�=/$���"O2�(j�+W͌�*&E ?�ҭ"O4\;a�ڑP�ApP�J$]��D�0"O4�q��=�lX3w�_!l�
��G"OL���K4;*Aرh��1֨R@"O�=B7
N�n�₇H�~�$�X�"O*TSV��:��ah�
e�!�"O��Q��Xdj��[�G��C�Ű2"O2Y��C�F�:���eװ}�	K"O�P��EE����gcO!;D��I$"OL�Z/�_�ĥ1wÊGR�w"O �3�搱uϒ���B��vO���"Ovh�f��'?�U����=0�h�"O��uG�8�X�š��U����b*OP���n� B����V��4!��iy�'�z����[�0Ts�a
��T���'���"0��+}�^�Z��I�Р��'��@{q�ێ"2�,KAŦ��!�'��� !�0I�`���3��h��'�p㖀� [t�z'ǵpy(uz�'4�A��͌�X�&�e�X!b��'?ps$��#i��Z5��体
�'[t�74�f���B&[��Q
�'ŖQ"AB�>k[�J]��*as�'��Xꆙ#?�xP7��(r)��'.0��B&^��m���*�8��'��l���΅
�z��Q���&�

�'o���Q�8�&)a���6�x	�'E� q��?t�0�g�ٙ� � �'��UiuF�_s�	ˇ+V�=Z.س�'9����4pf���'G�>���'*�3���w�P���}+���'n�D����|�ڕAv燷j���
�'t�����@�����WO�<�����N��peB#w��-cq�P�~� ��!�X8
w�q����Ё��X5^Y���$�8�3Wf/D�$pm�*Q,��8DJ@	<2ɨ�e8D���AL	�/gμq�ݓp�(%c� +D��ٳ��B$I�1����D��9�tB�I�0�������@טᰲ��5F�B䉺H"�P�*	� 5)E�˥,���RR�	�Z���{�x��!�
�^4��:"�`h�?E���G�{lZ,��HX	k���AمH	r���&%�ICz4͑q�<؜�i�듦vq�5���}� ��M	���	��b@����:�i?�xy�MV)/Z�y��
B���j�Bi	���"+X ��'3O�e@#,ݙ=Zl�D)��,RBu�I6�ڍ��'ŷK�Y�bU�b>��61�vo�O�꽊aH�)�Mb��i�����-ު���<�8-����9v�Hd��c�����;�`i�O&��Ӫ_Dԕ�F!D�H�V�����}����]x~�����o����`�n_I��`��j�� ��M˶��%	�h�֪l���&ҧt� DJ�F��1�)[�l}�6�J�����h�"2�6u+ڴ;T��ݦ˧ny�>J`�UC��SY�,�qJ�`�����X1��e�3�0(�ji�9�����KׅL�W5�U�f��uڔ�2́�vY�$XM>1
çc*����S$	gЏ
�!6!�^�Ɏ�1��S�+zl�j���v$x����D$@N8�Op���nD%BJ0�'�@�O!b,�� 4�]y`�����12�?�~o�9{�͘�͏�k4��֔~�I?5�Vğ\�<@:�aN.b�(��I�?��ɝ^�0��ER�)§_(}�ƂR��}� (T�>�b!�Ke$X�؆��=	���c��zB(��_ml|0-l�<�!� X�"��=��|˴�i�<�pN3   ��   
  d  o  y   �(  2  �<  �G  	S  )^  (i  �t  ^�  +�  \�  ��  ��  !�  ��  ��  ��  �  _�  ��  ��  6�  ��  ��  !�  ��   u �  b �$ H+ �1 �7 > �D �J GQ  X �^ �d Zm bw �} م ^� -� n� �� � ��  x�y�C˸��%�RhO5d��p��'l"�I�By��@0�'�F��L��|�t���pd��46����e�X8��Gߡr.����F�EΙ:��-Rש�-�u��[�}	��@Izn�$��Q��v�m}����"e
���m�� St����S�A�dCg�K�б[w� ���O��6�J�tRTb	��@1'��|rw��Q�^M��6n����7��6%�47�>�*��?Q��?1�R8n��G��
_�D���Z�oD)���?���?�,O�˓�?����?��#���b꜋C���rt@��?q�o��FX�8��ڟ���!:��'� ��О
�P�B��#DBLZ�'�Nm��O�Y�v��A��3;�`���~TA`ؓ`{��H$�%���,Q1`�io�\���d���b����j5#H�y1�&^៌�I���I՟x�����H�M��$SS�U�v1��f_�O���I��M���i|�7��c}�m�`�n��Mk4Y��%"��y���M�K�l��b�~�'�f�
T���bF�3c��t��U+�.	~x��Gx�::uY��J�~ِ�ӥg��?����3���_�MsB�#�O�T���'a~�aޒ��}3����B��A{e ���O2ʓŘO��)P �1J�9���(S�����hO?E�RC�`flJJ����!)n�'��I�{�j<x�4E�8�&����E^�p�LƑ!�:L����D�O��dg>�c�3Ob�GAz��E�'���W�,pZ�o/O�Tڏ��;
��M�d*�)P�<�M�Pax�-���?�����D� U��9����_]R�-T�6N�X�HE{���dW �����!1o(���P���?AG�'���8��^ԴB�dʎ"��<J����'׶���	��Z���Hi�`�EQ=P�Ha"��O��d3�O�-9A�)�n�I�.޳?3�0"OԱ[Q
XVS�)곧��ax�x�"On}���[NZ�{U��d|2""O>x��\��tJpeɯJ���S�	5�h�� (3�
V\���DٱU���'L�L[��4�����O�T0�a����|��c�Är϶5�ȓ|K�𘰫��3���_����ȓS��E��+];Ҩ�ԦԜP�`0��[�xV�����I$���@��! �yj4��,O��Ռ	f�f)�'L�"=E�$�^H�^%re@�h��-ʣ��*z����O��Oq�Ay`D�:\�����(�X�""OL@i��Ur��0��D4w�h�� "OfuI��ݺ.��YɣP���B"O�sa�QO�������S���)c"O��E��S�$� ��"y����|B�:�ɢ ��ٰ޴�?���}�E%[m7��0��ѥ8�~�����D�O��d�Od�e�$i���7?OD睘\{���kR�$B��#Ec��/�V��䆵j�꤉�J�5({�����hH�!�<�\x+�l�|?����FjD�=q�����M�6[�(���`Fx���b�O�N�,O���2�)�'�2�!�%�R��7	�P������MKV�)�Z����ݗXO��b$�W&�?i+O�q���O���!�9O���"6�E���B�bq��N�Z�D�O\��7��$uqO>!��fS=rw���*�*sE� zBA6?Q7H�,c�n�"|�E�Zm�	 �3�2A��c~���?�����OI&]R���"�J$C槀wDO>��0=9c�ɶ#%l��.%���떎�_�'$p�}�Q�N�v+�]"Ca*-��,���1�M#���?)��v�h(������?I(O:1��
�6��
�0Q`��	T�m̓pJ�鉩2�Mb�捧h�,�QBdS��\c��XA�?LOy����9y�>�iC�1W����1�'��ɪb���$5��O�ʓQ>�� �U�,a�!D��z�&�2�'�p�ak��qC��3C�R�xm�t�dX�p���4����<��Ǖ6��xgL��B|�\cW�Y�D���͓�?!��?�L>���%,=��$��b��rFԜ��2`����H��C�)��I6	���٢�J$4D����q����g��{Ҍ�$�O.�I3V�v�pL�4*�jҺ� g��aB�'��'@�	���?�dl�	!��@K�L[�v)�,cq԰�y��]!�Z��Q`�>�X�Z���c���'n�I :+T�	@��BǼ]EBиSM*]�`x��oU��?YM>�����$�	��O� H�����	t��M� j��Xi@�':`����D��x}��� .ˍ����o̅%:axr,L�?	�y���w*q�*8S�����Θ�y�;j�N�h�TY�!�g���?i�'��%�2t= R���j'���L>��f�<�����O �Ý�(*������0�J�j��O�D	.g|#<E�����~�F!��)��i3���D���d[�g��"|
b���Z��9A���#B�9�mD\~b�3�?Y���?Y����+�(M�06>t�E&z�ۗ�|�'naz�E��]ը-�c��#	>��R/6��O��D��JD�xB\�-�n�v1�4b�*0��6�'�R�'BT�U�O���'��P����S�^ҥ+w�4V�Ȩ� �&l���'�)�Ph����Ϙ'$*��0�T�|@�S&̝�=E�D�C�
5��D�&,@ �!����`�l�ʡ�t�J�)���3�<6��ͦ��	�p�0�Iw�gyR�'�B����ޓ|T0��@i��m�v�R�"O��9�kJ!�ܬk�hR+T9*=B�\�D���D��~RT��b�Ҭc��@AO��^h�#��&���2�4�?���?�+O��O�瓃n����c�L�.$�%K���;�2����JA���p 0j����A"Y/�aW싕G낔��	�j�qQaN��	��\Bo�_f�жH�O��o��M�����D�O��hyi>_|��Ӄ��"l�*X�Tƅp�<��I�_L�yv`��(���e��b�	0W���<�"&L�n��n�O:�dA�E�j�a��@$^$�`�3�����<����?Q�O }QӏS�s$�'����#�׃s>���ڣL)2܀Ó0��,�"0�������83�J���.#'4�H��	'U&��O4��O�	⃭���D̃# �06��15¿<q����(�X�#���UNf�I1�H�1�����'���%L�8��e(�2ib����[�)��o��;�j`��W��?mk��
=Y���T�.z�x�s��$���d�� ���P��	ҟ��O���w:��UnY r��%��Y�V�8��'�֝�1$�'M��K�X� �*׸^t%?�I��H�6��5 Ƙ`c�a���7?�Qk ܟP��:�M�����`eb��@���C`��Z����|B�'�az"ϓ��
�W�ˈ�P�&B	��O��n៌$�� ��,o�i
�P�T"e��Â�4	Q�N~������?I�O��J\�\�1bZ$m���!"O�Y+q�J4B$AE�1��4�"O�D�E��J"u��uX���"O*ٺb��Z�,���?��
b"O�Ȩ��#'(�DOT�'� �Y�`[���X�4�z�d��a�����^�j�b1x@��?)M>�}ZFAR*m{�#QBS_	�!P���e�<�Ç�N.rx&��o6�'&�l�<�"�3�<�����J������g�<��ER?����b��|�@���`�<���@.���pq�X��LL�3D\�'��OX-���O��7'�i��ƉK�e0�0���'c�'1���>�`d�-W	
c��!li*�P5+p�<aS��:L@����١jXAPS/n�<Q���'�,�Q!J��+�b�N�<Yr��n�����d�~`�;��I��d���mO�|��ǉ4.649z�?�H<D{�,͈���:�l�(�By9�n[�<��9����OF�$6�O "b�~q�둣A?T9��9�"OM;7��2�,��v�щ)Q�B�"OV}��m٭&�Թ����)�x��"O(����@tƴ0I�ܠ0�A����h�r����ݵ6��5jQ&N�i��٠�'�"����4�����O��aV�!�AEj�*rd ]�;��(�ȓD�đK��Zi<�%΄������%�� AQ���Q��Ѫ�އyzJ]��+3��;���Nx�Z�lȉ>؅ȓ��#e��s6t����;3.��'�0"=E��l��P-�[e�6h@"P��.���+~$��d�O@�Oq�l��p��.81 �Pg�`�&t�6"O� f,0�"�Q����+1"7>�z1"O��Q�O��F�v��f�S_PplS"O4�
��Ͽ��()�;X6"T��"O��w�ƦI���??'H1�|2:�l[f|��!6���B7!�ʰq7��`����t�Ο��O�|adF5v�ܨ�͙+"U�'"O��녀��
R&�օ��Fpp�B"O��KR�3�@�d������"O�K�!�)NJL�aB�ly��aU�'���D��7むC� ��]�<�ÅLў�*2�'q4�;&/�;nq��� cH-�0���?a�NJ: Q^"Xvi�GM��,��ȓS��l(rd�!
�D1j%{�x؆ȓdyx�J�'D�ND0V,����i��u�jD����8Wv������۞<F��4ڧH61�G��t���+0�> ��=�ɜP��"<ͧ�?�����ܨε(�G9˼�Ph�a{!�\�mV��[���{��1���!�d�[�N���A*�dA�%,��r�!�d�s��*�%��u�2r�6R�!��<��q��9_,� qD�^��ɝ�HOQ>�@6�۲n�0�Q��K7]���!ï<9è֬�?i���SܧTR��H�R+bi��Jrl	�ȓ[�L]�`)@�ʢ4��d�){�t�ȓ1�Հ�f�y�\h��\��H�ȓ��#�{0�#��H�X$�ȓi��D sD��5���߇�d`'��S���%����>�� ���!x	���d��C�|r�'���8H��F|I�tEDV XN>�ȓD~�xx�LU�W@�1a�3B4�ņȓ�:XZ$��Z1*�j�d��\��ȓdA�1�g<�Be�EՕH^&$����?�b�s,iPk+yn��k��Y_�'�^����B(<�3�����xg�Y�-�����O���ĝ)T��<�i\2![���$���{�!��Q �R�	g��mX�Y��x!��+#�T���ӛ_G(\CFI�7Y!!��U�Xf�����.3:-�B� �џ�b���W~75� =y�杋b a������O�)�O���*?!E��,�.�[EG!'�R����P�<�L�/~��r�̞a��%( ��O�<�&Z?Cl�3ɓ6���dVH�<y��֪m�H@�JϽi���ca��\�<��٨?�z�PƧ�� �r@�F�ZVyҭ&�S�O��X�_�m.Йf\�fP�i`*O�IB�H�OZ��+��i�!��
��["��i*��j.!�D�G�$:�b�����Y�!�d�[��B"�X�W���ŃT2�!��MH��^�h������0�!�_�(Sƍ�ҋ��M����G$j��'�#?q&��J?�7#Z:l���ԫ!�|�����'�x�	w�g�D�)�����Ȗ"����O�!�dI�K�|�a���)�`D�LԿK!�Θ	��諲m���p���D�m�!���8J�>��R'J�?��\��	�\��b'�O�)F�X�T&⤺�i��a�R��%�IU�t"~*�>M�n��B�L�.��c��?�?����0?y���J�xI��IےUL��e��V�<�ѣ�*��0�/؇F��$f�P�<����#4l�`����:��iw�d�<a��.[�$S�DX%\�L���TW�'D��}��@#r�*5p�Y���UO�Ο�� F-��|b���?�O���i�M��5"6g�TSD�r$"O�8Gœ� š���m;nU��"O� r���L�%W�!�祐\�je"O�|bOS*�� �Ue�����Ҥ"O
��Ǯ�&��*��GG��0��^�����pixa�aD�H]�ͨ�m��'��˓o�܈"���?�O>�}���fRlwΩAn �S���x�<A�$y�`R���0�� ��_�<�A�>������T�cPH �B�Z�<�P�Rׄ�-	`5���T&ҠB�I#��PW��t��%�6ԉ7$�O0�G~�1�~r�� C�$ˋ��r��ӧݬ�?�J>�������Ix�~�zA6q�P ���%��B�I�wLx���ĳd:����
8٤B�	��|��DfX/?��)G�~(�C䉷z6�ܢCȊ�9^���h�J��D[ȟ�r̚)0�T]���1
��YqB5ړ*zP�D�t�^�� m���0	��f�M���'}a~���(:��@�J��t�V�I!( �yR ��0��X��@�le�1˧/E��y�E��, �>/vD0K4���y��z2T(��y�$�JG�����O4G�t%O1^�d��@!��?�ڜ���ʐ�?�Ye���t�'R���3 �BZ�,y#M�O�����!D�4�AG�:^�輛��^�`c�5D�Pb����P@���0)�3�z���&D�0�P)/J�6|��]4�80�O9D�H���@�<�b��6)y��`�N�<���)�')���iwM�=��Ա�fQ̲Ĕ'��(D�'�|��t�E��,͡��:�\@ "m½�y��1*N�6��AM��q$�-�y��.h���mC3JFi��aΆ�y"E�FQ�b�v��c��~����':���+	�o�����'�2K>)��	�q����8!
t$�C��]��t8eƮ{t��D%�D�Ot�?�'D�U�K�'p�PA�BѾ'\�P��'�li�-�<a�h�@S�Q/"��}��'6��!S�P�S�l�O=)�H��'��9&B�/� ��uc֯8�����6�J�J���:�n  )^��Fܳ�hOU��S���#夜(c�T(�")��p����?��+W��ypD *f�����h�a"��ȓ[:�黑H�/t4�P��z�����Z7��@ĿKސ��C͐'g~�ل�1�r�Ϳy�%A.�a�AGb�#�'C���ġ��.���p�̒BҚ��I5��#<ͧ�?������"A�P�m�����"1�!��G���U�)�?�^�[K��du!�D�Q��-��a�j��]���O�!��A<�<;agN�^���p)B5v�!��K�n����L�/;�(�e���.��I��HOQ>5�Ɏ&�b4G	u��m;�/�<�3e��?I����S�'L�F��1�O6@�|�Ti�Jf���G*\JW��"X8(p���e|>��ȓkq�u��
�@X*�(�5�ԩ�ȓ>�%siظp���˃.
;�Pa��;<�aE�(;�`[�*�W}�h%�����dA���P�HbbpiU,�<{'�@��3(&"�|��'F��s.����rf����T<2p�ȓ<.��(-2�}hF[ 9�TX��.��!�D�5z�<�Zb��Ue,���zUL����A	T���§��+�$�����?�m�5��0��Ԩ__�7��T�'���`��)��8��U�K�"�<���O�5{,��$�O4��d#?ʐ�z�J�4��$���>o�!�$��f���� .������H�s5!�� ���FQ�kV��؁�ۊ�"O�-	�P�h>!dG	w��@���h���YV�� �^�q����<���'�rD���4����O��
�$���*��=@�%�ׁ:[Ј�ȓ&���AC�
��Þ�B���ȓK-���QH���Ä�&pRL�ȓ
��u2�� �h���cW�J�F�P�ȓ%A�Y�ł�;$B���n�(f�ԕ'n#=E�d,�[,y��� m�>%8r,���Z=m|����OΒOq�^�@%��)>���ȕ<8m2�"O�³���O*�-z�숃p!B���"O<�⊃/t��1B���Ky<��"O��ʗ�� /�>u�&�D\���"O�h�!��'y�.�2�$Q�C�`-��|�.�1O��V1t���^��XE����!�����n����P��O&�Irb\��e ��@.��"O��i���.La��%j{���"O�a�ѡ�%	���P�9RgĻ�"O���	�х�TO�R�G�?����O���	Ҁ��P.S�F���퉙��"~���V�4 ��ℵ{�5(F難�?a��0?��ׅW�M�p-��6z�j�	�f�<�Sc6<�1:���@�<r#M�d�<���.4�b�c�H�9gh��L�<���_�$��{���^��h��i�O�'�l�}R�O>;���w���~1�9˷�C̟�D�7��|R��?��O����8S-�r��U�6"O�EC���1'�0����B��(P�"OXl���8mqr��U �M+n-{�"O�i�f��0�D8e�]�2*�`��"O��y򋑶d�D�d��]���W�����S�m���;�K5^����K�&�H��f�E�L@���� 9M�|����uǫԂ++z7m�X�����O $�Ch@ͤ�h�g�X1J��<���?a��[2�c�AR;gF {s�T7Q�Ni��O�p3�Ɋ-�$՛  ҿc�D帎���Wɺ�X@㔬\z��[��3��t��$�X�K������*F��m�'��L����?9��k�(N���r�����H�$���Od��$�)~՞�2�d��]������<X��}+�<�f�T-
��9�F�Z,�.(��̄}yb���yBk	�l���	�O�-��f�9@��d�e-��O�x8�p��OF�zL��i��!.6Y��q���O?�2�`�"�dl�3�H�W�P��7�q��S�k��P<y$�	3M��EG�Dd@�l��eb��Rw��a�ĸ�y�X&�?�����������(��HɄPa����T)��#V,D�$Q��Ʈ �<�C���2n��1�d�+ړQ��?ݸ0"B�R�$R�i���Y��b�t��%�	���,�XQ�ݴ�����?�)Ob��`��M�d�BP��N�L.x��b���hm��1IX>���`ڶa`�g�'�
�H� {e��(�&R�z�d	9�(�#mb�u�uЄK����	���!��E��g��X@c�9��N����័�	x�����C�#�J5:�&_�#�CSk���y�H�46�r<�Ĉ��
�6P�r���?�D�i>Y��Vy�Z���Nd��{VO�q���e���M�tc�?1����D�O���`>���*�F��QY&��zNdys��]=h�|X:�$��u��MФc�۰<)F�=/��y��`��Qe���;k�d�(��	)��2� �(�ay"DD��?���ʕ{Q���G�\������?1���'��>M
T��m��A�4�3w2DȰk�<)7J���<�YSJ��p0��3T��gy2�rӎ���<!���4A�����HϧW�D�ȕ�ո�,{��A�K�p�'�b�'R�_=kX�{ĩ�m��`ԧ�$�"�̘��K�f��TcF��4��O$���C/��!���D�S�=
-@���c't=0w�w��">������	b̧C�B���v4���ȃ�¼x�'@a~�
�qܢ�@��ֱB%.�zWЧ��>��Y����M��Z��+e������(��@�`y�?I���?Aņ�	g|���oϻG� ��DF�?Q	�'�����N�H����<�va9	�'���qwEN2S�~h2"h�be:�h��� �)�I�.!&�q��ôf�dM��"O ��l�*Af� P�؞Oxx���	���*�)�e[�Lx�^Pn��F�#�O&�I�Ov��3�d��Oy����H���`"�*ƾOfC䉘2B��cR%�i$�@cc�ކYe`C�ɮ2�D�6N�F&��회P��B�	&)�a�@@��(ؔ���6G�C䉟�R6��minPQ��Q�
��5�HO?��!e���D�[t�
Y�����b럴P���� ��J�)�'J,���$Gw.�@G%_�r���6��'�ZT��2��V;P�ȓiM��i%&�U�0�rt B�u��L�"���&^��z󌗾	C�M��	���O�3|�!ʺ��ɗ'��c�Dx3�z����5�4l�>1OrH�V䘸8,��R�/����?Q��x�<dJ0�h��|���U�PU�s�� �L���z�'��T�r�v�OPB��m�[��Lp5o�,��*��$ʨWR�'��OTp\��JO _P\�q�R�~1J��'�R��+L>����$A�+c�e�ш̈3�0m��	7��QL��dh�5�X8\4���,O���O"��2��D~�E��o*����ǃ<D2�����׍�0<Y����'��x�fC3F�@�tG�<!p�H��i߉'�|�|�g(�u�����,T�(�̗x~�	���,(}*���>C�^A�hO�1�L�2'Ν[-(Eєm4?�e�>Y%\���H����`�C�V7��B"��0uMh���>���Ot�}�7;��J�e�:Ln1�� �n�x9�c�S��AR�d��j��>\\��S�*G�Z�����e6��D�>:��n�E��"�?�ҙr�+ZC�1�i�
n��.�����.���:R���'P�7�ͻMވ�PT'�'&=v�����ɟ	�f�'gn#���V
Lz���#�Di�!���4���)��S��'RX�q�OP@����2�L�h��H�� 0��˓"H,��'�	E�d�I%q�B9���	#�-�r!��?�N���h!/)?��y�C��~�J_�1�֌�f�'��u*� ��?1�/�O�}X�Ê8%�bMR��O�a���b�"O�Tש�	� Q���9��uB�i�r�' �	8��i�|�+��F���Z����(��8F �M+����2��3�i>7�̀6Jμ{֫��,(�5�d�9%�'Uўb?�Ӳ�A:��z���
�td��:D�j%船.lr`�'�W��D(�
$D�lDnJmR� �Ǝ�OH��ԉ7D��r7Ę&:�Q�
J�E�4	9D�,�qL�@\x`6�	E=��<D�R�g'�${���0���p�:D��1#�:"��	[���&��t`e+:D�@HG�W����!�D2� £�9D����8�b��q':�J�o7D�����G�k��e0�jɆ�d���3��?���?y��?Q�cK�^�$,�2h^�z�
�J�G9�f�'��'l2�'���'mr�'C�9I/q[� >h'h�CL�;i`�6�l6M�O@�D�Ot���OJ���O����O =Js��c�(M��@
�7�乙�&�Ц�����	�������t��ǟ�I��30a۷(8�I�&��<�<�0�ʹ�M{���?���?����?A��?����?q儆5Q��8��|Y괩���<J��')��'0�'Z��'���'��'ʻ}Tu£H;A"@Q�XO��6M�O����O��O����O0���O��$� MBBAs@rC�6��g� �l��@�	����ן@�	��d��蟔�	3hTά�ք�$�*��`����=�M����?a��?���?Q���?����?A���Th)��jp�!�P�H~���'���'�R�'���'P"�'`"�
�q��=i��N�����[@7��O���O���O ���O����O����;ϼ��ʟ*V�u��&q_T�mZ����I�`�I̟ �	��`�����ɳw�T1�	�e�8�ۢ'52�"۴�?)��?���?���?���?���>9�(�/Mg�vĈc%�x%P�U�i���՟��'�?���IP6e꠩��̓���E��%�i}]����Y�'eA�66O����?0dN-��F�#�X�p�';7Ohꓫ�'35���4�~b�*�~Ř�)vs������?��'���d[��hO��b�x���M-U��h����L�3�E�O����"�����D-� � D'G*k&�����C�L����V}B�'f�6O�ʧ0��}Q��n<�yiǧ̀`�r(�'o��31����O�)���?ٗiy�`r��X:�s��9fP�'��<�+O��<�g?�4FΨc�P�ѡ�"�N0L�ߟ0«O�ʓ-������b�ϟ78�Ը��K/]��	����O|�D�O��$[/Y��7�+?	�O���iݍ���D4ӗ`	$�A���!ړ�?	.O4b>" �%�V��5nB���i�G	�<	[��'��I�>F�%�E�a]$��c�dZ���'���'��.ҧk���q�j�-2XX�:ă5�������/Z��Y�'f�'ݟl�P�|�W��!p�S�SJ2!w)	?S�VI���Tޟ$�I֟���ҟ��Ieyr��>��Ho8�Qj�+)� �3�N�)L�0�i��6��h}b�}�&8l��?A�j��L�8���Q:j�\��ɋ/m�oo~r/�/hV���($�Os�#Z�n���W2  dq�KW�O��@�+N�Qs$�j�.֎D�`|�4U����1���<9"�i�1O(mpEMO����$씣Җ|��'���'��=y�i��i��q�GށM�^���R�Z����3�A�������"Y��9��)�]�g��je�?�T�(�'���?٨Pᙣ_�h�zČTE��$��E�<TZ�����0'��O`\xxՀ>8D��FC�_�%���fp���ڴ,:�	�?��Of�O���b�<�̭��cɲh���Y��?Y��'{�i���!v���K�g,�1����$Nʦ�?)�S���۴�Q�D�A�7�ĳҴ)0R��Ѧ	�ڴ#�4��Ę�VD�M��'Ҡ�|�	@ �J; ��x�㮑�OE^i�	Ay��'��'Eb�'^R�?u�a�'/L�SG\�R�y򗅜u}R�'���'��O�r�qӜ��p���xe��=B��� ��Ѩ�K�O`6��}�)�i �+>6���D�qn� D��Tnr`<)�F��O ����?Y�3�D�<�'�?�VJ߸.�J�(��Q��Z���N���?���?�����n}B�'��'a�k̘ap�dhP%I�RB�)c���v}�'��)�$֕3�Z �7#��4�*<��ߡ1J(�y�fh[0�M-�ب���!ڟ�QW1Of���;C�b`8�Ǝ)M!�%�'���'�r�'�>a�~_�Μ�G�7��#pl�I����<þi��O���U�?�>��R�W9t`nxa�ş0��K��%#�4\�v��: ���3O��${�l���'=������O�K:�Թ�EG�EM�!Ʃ#�d�<���?i��?i���?�1�@�}INu�f郕G�IJ%�����_w}��'-�'���y�]� �l)A�� 5u$X��)#&,���?�شH�ɧ�E7&�θ�fUk�h��\�L�+f ����'���"������|�]��pB L,BЬ��1(�T�:��aB؟��	�� �������}y"f�>!��za�qj!�Z�A�ha2a+c?H��	қ�Ąp}�'��1O�9���:r6��w���a� 5H�$�Q�F��4"�)s�Q>��;	��fFK�F�<�hE�hh:��I��IΟX��ڟ��T�O����e܏	� ��� �������	Ɵ��O�˧����$�/x��sa,��K�	{&��q��'��'�2�8OB�Z0H�(|�f��2k�2j�-4�* :�E���~b�|�[�������	��1-L=�~|3*@/j�8@���D��yBb�>����?����I��r���`GQ":���jg��Y������OV6�@Q�)���܇]�H�1C��#e0"�S��K�D���(3����r���OHYqL>Y��ʴC�u��'INA���@�?q���?i����4������h`�"/?��c��/��b��O@���O�1lZ~��v��ǟ 񁀁�S��pe^�+d!s���D�	�[<>yo�D~Zwl��xE՟ �\Q�@)�'��,��#�T�9"����Ty��'c��'l��'���?3i�TAv�N70�h���͓c}��'s��'��Oq`v�h�I(~��ě�f�8�� ���*5�����O֓O\���T`�lt�J�I�`j�l��nM�my �6÷M�$ɶ9��P��'�'d�i>��	�4��bgk^[�D<��⏤\2`�I����	Ɵt�'�N��?���?	�KR���m�c/D�uD@("k�:��'qD�=�f�~��%�l�B�^#x���ӱ�ڂݚ��[Ɵ��I(��)�Qo�q��L�'��4A��� �1O�y�V�/G8�S5�P�`$�Iq��'���'8��'�>M̓��$�fǡOTI��+��L��I(��d�<ٶ�i��O��i8#�8�0���% ����_�����O����Of�CW�n��{�f}�R�~��&N--V�4ハ��^�ѳ� t�	ry�'��'���'��
ڜB����3AL�|�#4Ɓ!O��I����O`���O4��d�D\�|�^�9`j�,�Z��HX�&@`��'[��'�ɧ�$�'���̿H ��A�A�$��=�p�ީ>����#�iH���z����w�O<�OL˓e�����u�Y3e�la&����?����?!���?�-O~��'0"� d̡��I�'NU�b(Ȉd Ƀ�'�6 �	4����OH�h�t;p	@�`*�%�NI���C�	�`6�5?q�Ϙ�!��|r�wWh`[R�<QL������v����?����?q��?�����x��0�?L�4yFgEW��'�r�'U���?��t���d��@��j�W�f0�ġ�_�L��'P�'�rcz �֖��[ %��~� �������@���,I���G�Ov�O���|z��?Q�[A������1'��8�+&E��0���?�(O@q�'.b�'+��?�/ƃk���I����,Z��<��V�\Qܴv����!�~2UC���SB�Q:3�,H��FL$'�L�QƁ"�3�O��Ɂ��?Ig�3��Bg��@ ���q(�ZS�@����O0�d�O���9�I�<!��''`A8!�ʙ{�$e&�S�@b���Dܦ��?qV�02�4���xqFN�C
ui4�N-EY�0�i'�6��vP6�"?!aE�I�i/�)D�s���r/�DW0U!'K%J��^�X��ҟ��������۟��O~h�dK�**y���*3��@�VS�X��ϟ��I}�ϟH!�4�yB� 	4L0q����9�E�4~��&�fӌ)%�p'?��&jUĦ���0�R���!HA���$�`��(HU�� ��'F*D&�����4�'��d9bċI�.dk�GX�\��* �'�'5�X����Ol�D�O����) ݪ:GS�K�0T#�$ڎr�H㟔[�Oj�D�O P'�T9�J�(sRީ�1��!):T,@b(Mly�bG�*�q�I���4�
\��C�`牅+��ykT�b8<�At(�'@+����O����O��d=�'�y�`ΩH�*� ��8d���P[�?��Y����Ɵ\�ش��'#���	�حr�j�} �u  #ϼvR�}�XHo��M��f��M�OZ,3`��2^wĎ��A�бfP�2��N�\�AO>.O����O��D�O��OP�3Eҋev���	9ge$[֮�<��V�X�'���ɔ�K��$ڵnʋ~�`� � `����'�b�'�ɧ�OZ�[�ϖ�ġ���V�B/��³V����<a1�s	t��_�	yy��\�6}����-j�`�3��R���'��'���'��ɂ��}�Pp%�G�1Һ8zU"�a[|��B��O�oW���Iڟ��	�<9'�݀*<��Q�WƶE��`�/CܸYn�o~��1��EG�d;���O�}܈�B&����(���'���'���'�b�S��N�(�����Dd\*3Nf�d�O����v}[�Dڴ��'�`����V,�a�t�3n@����x��'���O�`���ix��'Wj�`�钍/ry �,$Bl�nG��'�g�My�Ok"�'�G�)2���w�܍?��,��"U|���'{�� ���O��d�O\�'!�����ΣI�fd3��σ:��A�'���?ڴɧ�	ۆCUr,cR�9����jˈi�9�C79�P\��O*�	��?�6m=�$�zg8�
%�Un��9'
��tr����O����O$��#���<���'n}���>(T���)IG$����?������G}��b�"�j�I�IQp!N���$�rf �-�۴Z��P�4��ę�<Ei����'D:��խFR�j@�����ay"�'��'�R�'���?���!֗e&�|b'��+%�fd�bo�i}�'��'���yr a�B�	:"(��c�@�3/Z��^�U�M�OV�$/�D3�Ɉv��7-���Q�ĺ�h����7V��"��ON���ұ�~"�|rY�����D���R�=w2�IP�ߋQ|4:o�@��ҟ���oy��>����?��i��$�A�X����n��r;��ьm�>�S�i�7-�{≌1$�� a�BRĘ+N�-�'�
9JA��18�k��Ԣɟ�k�8O�Bu�"2,�٨� �#��4z�'�"�'�'v�>�͓1W������
��@!�-d0��	��Ŀ<�2�iW�O���J�2+�u���.!@�	�G�U�F���$�O8���OBꥉl��k�(�ql�~��#�%ވXw@A�;�z�TT�ky�'��'��'q2��w�u�V�[6;��	3#�-���e}"�'6b�'���y������H�����7kй'�듀?9����|2��?YtoH���cP3րU�V"��!��4��Ti�P��'M�'�	���]�wn�%c��:aFƣK��I����H���̖'����?��dl��"§ �l����?)�iF�O���'�R�'���r����eG8%�YcR�.�<D�!�i���o��%�'�S�Q��5��ճ��ɪ)Q<YAa�F�H������	ݟT�	ܟ�G�4D��)�Hl�Tm|$�Q�]��?����?�wS��'��6>�mb�{�@E�p��$zQC��P��O��D�O��Ȕ&A�6�"?Y���9��$��Ƈ�[C��jV��6
��|뒫���&�|���4�'<�'��ҥ��-y�4�BE�L�����'��\����O����O�� :d��U�v���W�LE
0�Qyrd�>���?aJ>����cW�+9jZ�!6"���ˑb�4v�.a���id�	�?!���OD�O���C��F����	��d)�@�O��$�OJ��O�� ʓ#
� TA�q�_�:��܀�/�59��rr�'D剱�M��"/�>9�).i���L�x?�|��O��#�������?�Q	��M��O<)B�ʟ��O��=@���/B��1�fѦ���������OB�D�O��D�O���%�t�ҧ[p"K/I���xC��,���<�����O�6s�0��nY�I�J�!%e5H�m�%��O���E\��W�S�f�m�l?W�Г7�ƕ��M��RE�}k�F�џ0y�j�Y��d�w�I|y�Ov��^�s�FLc�/�঴����W=��'��'��,��d�Ox���O"���ҽOKjmxG�3���	�E9��������U�شZΉ'��y�K�I���j�W�-aY�4(bJ�0t��4�%?�'n�:�d	��y"���a&���J\5���5��3�?����?I��?����p���EV:?����.�ahR�[� �O<��'���'{�63�4�@�	�7=�@�8"jDVY����;����O��d�O-���tӬ�	����/wd̧l��U��!e$�$ju��!J~�A%�4�'QB�'���'��'��0��E�<��ugM�`*�ʣS�Xz�O����O��6�9O|py����:P\Y�C� �Qކ��E,S}��'�r�|��d�"T<��يk�����p�l�:�@E���D�+T��p�����O��`��E�b�Őr�ܬ�e.DTPb���?����?���?�+Oz��'�2ŋ���f��{k"�+����I?�M����>����?I�'��{�/�`�)-Quqd��8R�o�x~r��
c0�'�䧴yw+X��Ҭ��D�+�zxX�.��?���?1���?Y��?)��IΤ�����9,c����YI��'G�ħ>i���?�þiI1O¤�Um����5���grH��$�|��'��'?4H`0�i��i�ҥ͞����i7�Òs� ���n9|^���䓯�d�O^���O��Dք.��9��'��'��i6˛#l���O\�z-������Iߟ`�OG��ɋ�Hf�c�A#o�R1H(OJ��'~Z7-UѦ%�L<��̔�eQ��Ӷ��5a��	ό (���QHY3�����lDs��cz��Ob��b��"�1B�b͝*���x�!�Oj�$�O����O����ʓq����:4v�y�G�*k�:(��?�+O��mZq�.k����P���2?㰹����PK4�z�D� �I*'�6�n�n~2�O!l�:��~2�-y��pC"��;A6,db�Fߟ̖'���'Z2�'���'�����;�Fal�	��U:Ud�t�'"�'�R���'��7�n���`R�^IB�h��x���٦+�O&��4�$,�iq��7M��Ѓ��7	s��CӧܚP��OHx�3g�?�~��|�_��Sş�hRL��p�Ԍ��a�� �
��%J�ԟ|��͟H�ILyRO�>����?���n���1��U6k��1�Ӯ}�A��̿>1бix7�Mk�1,�*�R ��(0��C�\	��c�<y�`�:�p�'h�f~�Oj���IM��dƍ3o4� e���7�p�C".S���'M2�'o���<�p�O�dp\pI��vD�д�I����O@���O�5l�{���zg�C���� "j�/�P�g�O�?���?Ѣ�i����C�i���O*�3@))��Xw�0C�M�:3!�p'��l,^�rN>A/O����O����O��d�O:�o�<g"tPal��s%ؙ�s'�<�aU����۟\��F�۟�sa�!;Z}�%��8����vN���W�;شu܉��Or����Z?AL ���*�<v|h8�����O�< r@���?�'�)���<a2 	{RbE�%/W<�����?Y���?����?����DG}�'�Z\�f 7~�(h�w攸1�����'^ 67������O��d˟x$���b7�B��8'QP�APL!D
7�2?Y�FJ�a��I9����ҌK-5�t��GG�	`��c��
����I����������,D�$��(Ff�KG��-O*��I� ��?y��?�V� �'�6�6�1w��SD��! y��y�FƟ7#6'���	ߦM�S�}R>ToZv~b�X�oV���гdrų��*5��8��ɟ�W�|�]�������X"��0
�xUp#@�'�\=@7i��`��MyRb�>�,O���!�⃄,V[�q�6�^�-�v�!��oy�B�>1��?�M>���I�����X��~$�3��t�"�i#�i+�i>��$�Ov�OR1��I6�H�#�y������O��D�O�D�O,��@�^� �*�}�qeH$Jf��ժ��?�*OV�mZn��Of����\;B�� �8���#h��)��Ė˟��	8b��uo��<	��vAbT	E2��'���X��Lx�5[�'B$֨�"�'s�Iߟ��	�����֟���A���nX�鵂��b���aNE�J����	͟��Z`�i��d��	lV�����D���!˻C��'��'�2�'��RI�v2O؜)��63���bu#�6���`��O�mCB�J��~Ҟ|RU��ӟ���錮j�А��Oǒ:�L�ڟ�	�@�	uy�ʳ>���?�@(Ρ����5:B�t%U;@�����B˺>���i�v6SU≕��s�V?*����Ѳu�<�����آ���,��yZ��7?���GZ6���/�y������a` rn)�� U��?���?Y�����<�  p��Sg�=��]�^����'������]�?������a�ҺB�:� ɯfh�R���?)��?�I8�M��O���+[�b_wE՛s��ZC�M�6�W��A�L>�.O"�D�O^�D�Oh��O�H��m� \�d�#vZU��k�<!�T���I����K�s�<ʱ ��1FL��c��'� �z�����dF��q�4V���O ��(3h!ɚV���H+��3�����Ձ�R�����O�_	H�Isy�ޤ=�! �d"i��gnI�`�2�'r�'�r�'T�I�����O���嚆Z��z��A
6׌�!���O�)lP��m��۟��I�<QD���4�V��rl��"Z���0!�o*m�b~��Ð|E��f�'�yg ��L>0Aˇ�]�~�.�1E���?����?���?i��?����{~v�q��X�%�Tܪ®W�!��'��.�>a(O�]o�z���@r�Z�I	�p8�n��_�,�'���������a�m|~Zw��|�F���2x���K�!�a�㊃�h6��2�d�<���?���?)��F'��[�K��[N���Q����?����ăC}��'"��'=��5!U"�T���ay^�@O�O�0���� ��d�)����;c�(!yb�C�D�`@�1���㦧ԛ�M#�X����=���0�d��r�L�q'f���00ذ˹+��D�O:�D�O(�$4�i�<Y��'�b���G��l�۳!W2VZ�)b����d�¦��?��Q�0�ܴMq���`J�*��1��#�67��]� �iH7M�1XN6m/?�@
�%�����6����`!����T�,�N�"3 ְ<Z"R�0�IџD�	ٟ��� �O+�I��K��@4q`+J"T`�kV����� �	Q�s��!ڴ�yr�הH�0Q@��FӨlJqK�F�Kp��$�����?i��{�h�m��<��'��5�n@b�)?���(�%�)�?yc�E�'��$Y������O�d��z̛4떷.vr�Z�V���d�O����O
˓(���ߟ�����a�7�fTXv�4O�4�rb��T��A^�	ş$o6��EZ�J�Z��xp3 /���	ɟ��5eL�`�\�AQ�=?9��g����Ż�yɖ5j��{�� W���SW)���?Q��?����?����e��X�F�!4����n>GZ�Y��Ov1�'��I��MÍ�O�.�j�-�J?��(���v�W�'[2�'���K+��8O~�Q�:i�˿~��\�E�@|,�)%7 �c&�\��iy�'���'���'hr��5I�PY1]��ꀽPB_��ةO��d�O��"�9Op�����W�T))�B7�a�@h}�diӤuo0��S�'\X=�3)j���x F;{���VԀ����'	�`s����W�|\�P��\�P�:Ռ��E� &˟����	���	iy�B�>��Qc���C�B�}�$�`�A��XHBl+��!T����Q}��c��(mZ��?y'+E�h70�ۡ��D��20퍴pHބnN~"�`�������O��jg�th-X�X^xp(��b�'���'�2�'qr�S�F�:�FV��aɀ��~����O���D}��'��d��c��ᶤy3�j2|��#3� �O�6��要�Ӧ/�(o�<���uP����H&Qwz����G�̈���7^<���V����4���$�O��D ���	��|N�@'��'ep���O�G��Cy"�'!�S�UR���fO�L�<�(�o�r�N˓'I��ޟ��	`�)�d�׾VF�a�R��D*dqi�(I��훆
R0�`�'��$,U�4���|rL)ꠔ`%ʗE "��'A� #R�'���'=��W�lI� V.	��P@�.m�A�M�%'n|�	П|����MÊ"e�>�� ��Uh'FɠR(��k��ǋ m�l���?�� �:�M{�O�� U)��SR�Ċ�S����g�(�xt`N�?-O����O��D�O�$�OB�'B�84RbM�^�a�R!�&Qz�O��$�O��7�i�ObQl��<�G�
/2��Ғg><���I'��p��a��i�S�n1lZ~?��+ߍf�.�;�� f Ɓ��/P��h��=#y�$5�$�<A���?�`
�.�@ي%���0�H�eˣ�?y��?i����m}��'���'
�<�H�l��T���*��̐"��S}�'_��|�E�U���Lθara�9DB�ɾ#8�!�H�ܦ�PJ~"Sı�͓c�ތ)6�-����fR�J/���ޟ����D��I�O>�$���0���9�j�S��)��'������@Ȧ-�?���ER4y��F4� �Hua �m~�$���?A��?�E�Ҟ�Mk�O�j���9k���$b,{��C����X�h�$�ԗ'&"�'��'�"�'��py�A�,�6,I�\?L��X�`R����O��$�O.�d8�	�OTa(�k
�g}\�bg�٢O�$�cƢB}��'��|���ѷZ48�s$�}X�!J�fل�����i���6���`5$��%���'GjqBI�>}G��� ��}����4�'��']��'�b\��Q�O�d" Yb��fD;.�P��DE�)L���Aߦ��?��V����ڟ�͓t0�1b�+ :*�)3�B Xj�%� �����'�` ��LZL~�w� d�����&�$�:l�2=�ɳ���?���?q���?Y���� 0 ����>O�4:І���x��'�2�'CN����Eަ�<	����jLhӂ���ʭWr��,���<���O즱�'�0i�K�+8� �!���s�2�����Q������4���d�O���Mfe氺��ܼ~JJ�)p� �1J�D�Of˓���Ly��'�S+�Z(��N��G�1ڄ���!k��2�	ϟ���I�)��)x� ҷi����Ŗ�q�����ͯ*��������6���0���y�t(pB�\�)�b4��aB�52����OH���O��4�ɮ<Q��'�>�� aP��d�� !>�i����@��?�]�����O�VH����*5Tdx�mLq(���I�X ��ܦ�'�&1c���L�' �4��r�˨1���`EΣV$�e��zy��'���'�r�'���?�S&� `x�����Of�+�c�b}�[�X�	P��5қ4Ov�:'jϘm0FEh��Ȋo:6\`��'"��|ғ�4�FuV���O�ٕ+�+1gv��Ͼ]�\�R�'��$D�j?H>!*O�)�O4�p�]$���ZE�ƃ1vjx�k�O����O��<ѧU�0���h�	�L�|ڇ)i��	�G��?�R�|�	ɟ$�|bf�.uf�4:4HQ�djũ�sy��P;E-��7�il���JJ�'��W�Me�bj����37��X���'���'�2���<ɇ�Pr��7*�h$�VI韌��O�˓L��������7Ǖ+��Ҧ��(��!��O0��O���U�>�:6m:?���<6�~�!x���@���L�L-�/IRX�8%�0�'O��'{B�'r�',�بD��P�|�`՗vy��Y�Z�Ta�O��d�O���/�9O�ȻDM<��j��_2/;t�&��x}R�'<�|�O�R�'�!q�GJ�c��5BJ��А�R�If�֚��+VFCJ��D,�D�<S���{KZ�Ys%L�Nߚ�iVf�!�?q���?���?�����e}b�'����D9?$�gdR'54ZT�'�l6�'�� ����O��d|��
���L�B���$.,V�
3�Ο��6m(?Aq��.��|w�&��u�OR[^���+����l���?����?���?y�������4,$޾Ly�%r�b��'Pr�'v����D�Ӧ��<�c��#*�6�2֣Z�@'d��EJ�Iڟt�����k	����'��@{�j�1,X�e�TOE���ҫ�!d�T�������4����Oz�$L�{.u��[=x?F�)�@B���O,�L_�	�L��ʟ��O�0��%Źh���0I�U8ġ�*Oʍ�'�B�'cɧ��?-*&���+�#�ā�%S<�4����J��6̈́By��O�]�����L=�D�X	�8#u	�f�P�����?a��?	������E��, `�,�N��`��)��S�(�O����O��n�@�=��I�
�Ƃ�T�*WჀ@:���� �ɛ.� �m�k~Zw�T�"wџ�;�����|r�3Em�7c�u��oy��'/��'�B�'�2�?��U�ǆ4�Dس�nݻJ�xrU�TK}�'�b�'���y��q��	�(�H42�a�tҮ��I�TRX���OX$�0&?��Φ���h�(��Ã_�g�8��ߌJ`�@���?f��jf�'���$�������'.f�(q��)�^��(�!5��e2��'�2�'�X��b�On���O�$�	GuE��},�kE)ƕl4�8�OT���O<�'�(�GAݒ�0-����[�,��T@Ywy��VjN�W����4�����j��I�(S6Ş)w����Y�D�:���Ol���O�)�'�y�.����7��48�d��5ȵ�?Ip^���	�l�ߴ��'o�4���r�N��dY@�!ˇ)�7�"�'��$x�
�1ffvӊ�%�$�c���Z��(n����Tp�r(���Oxʓ�?1���?����?���:��swI��&�H��ð	Z�xy.Of�'��'����'��|[@��1,M��2bY6i[����ͭ>i���?�J>�|�O[8�n��I����j�:*Ҋh��Q~�#�.uA��ɭ#��'@� |�eE&%<jE� Mf��IٟL��ʟ����' ���?���m�v�A��
Zǲ�@!�5�?)G�i4�O���'T�7�̦y[��C�\
��Xr�E!⑅��P��¦��'j�8ԍP�?��}*�w�X5r^�1B���W�|`QK���?���?1���?�������@�)ٶd~T���/��a�S�'�R�'2x��?��%���% ��bE_90�V�*�ʉ~��OB�l�;�M���w�z�P�4��$W�:28z��V�������!}�� TU#�?1Ŭ ���<ͧ�?����?�g�ͽE����6��Ҧa�?�����^T}2�'���'���l�N�*D�S��� `����W��UI�I៨�	I�)����2V?�(JHB�y�n����j�)kf���M�_���ӱ��D>�DX�pެq�m��8-%c=D�����O����O$�� ��<i��'St��2�K�\˕l�*?������?q�Bٛ��Vr}��'P��Mʤ��xV��k��8f�'�r�W<W��v:ON�S�������򄛄c��T�q��l�$h��=�F�$�<y���?���?)���?1ɟ� �M�!܇|�`P�4됆4��XS���>���?�����<!��iv�d�7�E�KW)Lh����c�"�'��'JR�'���Q2c�v6O�㑧S��(&{X�����O�0`2َ�~R�|�\����ߟ����V�y�t@Ӗ�R����s�Dɟ$�����	Ky2�>����?I� 2(���ɏ-C�Z�/���#�L!�����榙{ߴ��'��\!�eA3
�J側H�����_� *5R�mF`�|�SlB��<A��I��-�B�>W@\BD�B͟H�	͟��	�`D��0O������F�̀bŶ��Q��'��듑?���bE��$��`A�tf��T"�$�Я g�n�W��O���O�$6\��6�8?a�-\ ��'&ᬩ(��ɀs��	P�!��~�Y'� �'��'R��'���'{��E�
1q������7��`�[�l��O���O^�/�9O `	䃊�R����Y�;k���R}"�'��|���+%+���r$��B�x��(��%��Y��i��I�P��[r�O��O�˓#���CE 5ޮqʴnX������?����?��?�)O���'�R���n�V4�!�\�|˺�{$7�ybhg����Z�O�D�Oz�ɺ<�ĸe�J`jE@C�<vf��ړI|�,�򄙙�N/�'�ygjժe�́�M�.a��%�.�?���?���?���?���ؠ}2��َ�8�IӤP!R&��'�2�>!)O�uo�e̓tV5� #��#�LH�i�<]��'����䟼���t��n�a~�.�"���&�z=�3쌢Q�d��e!��D��@�(">��zE��Qք��
*�ZQB�-O�A� 	�4�K�PW�P �eNN����/�[ơ: ��c2>�@�T�*�f��5��	�fbAz�f@�e)�wZv�����wn �e��R.B�2�
�Ȩj�kS�s3�]�vE[�L�F���W:�u����"gC�Uk����)�u�`iV�g��҇)_�&����v�7A�Ќ?���a���Qs����bE
7٠@Q/R�� i���>t�R�+�J%��V�9��̒p��q�8u+�y�lE���-
϶H�W���Z�ZAx�MT�0��l�1�`���K�)�m��j��ّl���J�PU���$N)1U5�C���S�X��	GΔA��	7Sdf���E\�$�q9��M�rւ0�e�eH�u؀#�I�I���AB(i�GGY�ڑ�5��<~;^� ø".6���[��9td
;��<J!�^� �0]P�H�&JS��Т	Ȯv�5�C��O�����g��h��!H
	o���o�Xx�i!���,�BQy!�O����O����O��D�<�7䖭H�)�Mܱ`f��J�`��?���?Iƀ�~���i/$I q15&W�S�Zţ����BN9{E�O�����E�����It��OL����q�� R��X!ƜhTƇ5�?Q����'���o���ןл���5)L�A�"� *k�e9Pj_�����ߟ�I��x�'{"�'X�?Ol�`�-�"äP[��V+{$(�'�'��'a"���'",�ɟ'<2�',�탃���C��b�, �4͏B$B�'�£�>	)Oz��#��@� :B��9�`K���<R ʓ)钼
�o_�Γ�?����?ɟz|�g!I��\x�n�F�b��'ޔ���D�O��O.�d�O�᯺(T�xGFK�9�̱�oܩP��ٙ��Ji��?���?qO~�O���JSl�+�-�,ؿ ��a���?����?	K>���?Y����y2�
#���b1B�$��@
C�A�F�T���?Q��?�K~R*����A�1h���
Ƥ6B���̏3{���$�O �O���OH���4��8��焄�W��0Q�#�P�����O�DԬj��$�O̅�O���'q�bբ`�.���ԑs���s$i�/��'�2�'ގ����|>��2y
��D-�b@���OP�h�>O���Ħ�	˟����ORd�ԫ�.������ :b��x ��O��D�O��a*��c��!D��z��ŌI�8�k�c�,3�L �a�'�"�s����O�d�O4q�'�剺<�F�ɢmK� :f�WdZ�dC�Q��=A� �Io��]�D��.�yB�'P�t���ٺ7����)�cp� P��'���'��'��I��|�Iܟ,��^�Y��UR����/#:ޝ�?�aH�*�?�D���<���?9�7.h�" ,��ɀt㗭&m(�����?��,4�Iwy�'{�'B�Y��:=���pG%k;X�Ҵ[�4��ܟ��l�@�������N���V��=���!3���a�Z�?!ҙx"�'�r�|2R�y�/L�T)I�H��nNF���O����'vJ�	˟���֟�%?�a��b�b0�E�4#���i�?���'���'D�'��i>��IpC�2s*��^�0|V.˹^�LE���t���ӟ4��[��=����O u�k7$�t�; kA��u��O��$7�$�<ͧ�?�ϟ�1�@�@_Ⱃ����^�<�)��'M�'�Ĕ�Y�x�O�R�'I�.� 'i[��Bz F�S�(І��'!�X�X���*4����n�Z��>p��dq�.ģ)O����O��d�OV���<��F�D\��D!�?v�Y�EB.�?���Dɶ*G��S7I�d��S��t�Bӱ? ��զICy"�'���'��'�)RàL!�
P�"/©\뚰R��M	��dUwX��
���&H*�(�k�����ǶAȬ ����?)���?���?	�'6��*]�e�>�����gVu�o�'}��d��y"�'D��'�4)�s���)]
�+�	K#3�\���'U��'v�O�S]�U�? ���M_7$���+�R�2Ȩ4�!�|��'V�Q�O(�$�O��i`���C�;\�H �	4*�ybv$�O���?���'��?O��J!-k�`А焐&��Y�'�'-L�J��ٲ���O*�4��ʓ��T$Ƿl0��"P��?����&K+�?��?�2�'?�I]�@�⣃�}�����E3���	�#S�����������%?YK�����J2
���F��;^c"�����('��D�O(�O���|����i����i赁�\ڡ�G	Ǯ\���'RbN�%�y��'���?���y��:Dp�Qj�.�j�"ي�ۭ����D�OH��0�9OKd-�fܚ��D�X� n�sUf�O�1��<����?���?)����Ā�3�&���R�W�0�eo q�"�D�O*�z:�Dx�O��a�"�P�[�]+��>Q[(i���I i��'2�6��O���O��DT�?��Q�9�
 ˅
��
����q��O��$�OV��)�4��AP6OJ���J�:����4�����G�b��lmZ��	ӟ��	$��S�49Ot8;Rf����t����$�؁ˑ�'HB�|r�'�x�0��5�4�?y�2�6�xF��(J"@,� f��F�y���?���{a����>��ٟ'��ر�\/�-Z�7\Vd�O���ވ#���O`��O�F��0�P���ܲsQ��[Yx�	����<�����OD�$�O�!��S�^�&�X��[	V�,x�'H�W��7zм���O.�$�O$�ɻ|J%�O$�슗�D�A�~\�N:�J}������O���?���?YĨ�<��c '(�:�q��]@ji`g(�3y������?i��?a�'��I�P�t�'Sl�CR�_��Q`�L�9����b�'T"]�x����T�	-s�b�y�D�_Al�@��@ 6yơ���'�?Q���?�d���<I��+B���x�Iڟ�Z�������^��l�@�X|yB�'z��'���J���'��ɛ�t(�1�IͱBW���#8�Bn���y��'L�7��O���O��Vq}B�rB� b`ò^*�ʴ��!c�2�'�'���yB]>�IW����(C�ar�!H�&y։h#kMy��c�'"�}���$�ON�D�ON��'y�Ɉ<4�-���u9�U;7�4Ye(A�	�j|X�	u�	r����y��'��xa�lI)K<v|qs	�1�4Q+�n�:���O,�$�Op��'<�	����_�2 AێSN&Y��a1]��`�	�1�牟|�J�	럨�	� �5�T2@�2 q��3�.�US� �	ȟ@"�Ol˓�?,On�݉yZ�SժЍ}��Aؤ�	�u������Y'(L���?����?a��<i�D��k�h���C*lĎZ���?y�^�@�'B�S�D��ڟ�	�#���=��2d�˽9��P#u/c� 8����8���ؗO����"ti�/=���W`���[����ܖ'@�^���	џ��G|�	-���I�R*� G$L;F�U(v�a�p�Iȟ|��z�S���i�O��r�D�>�t)*��� �+�?)�����O����O2�20>O��z�pbS
� O�5Ҧ�S>B���j�O����O�أ1Ob��f���'��'@z��']�bH�3Bk�8�fT��X�(�I�(�IK�"<A�O `���E� �Q#�1��^Γ�?��ivB�'���'�F�7%;�jD�h���+�MH0Wxz����?��{
�������O�'B���0T��u,U�sÃ�s�z��eEA��?���k4���'���'s��&��O$�P�hF�"�DP�5eA h�E�OX@XF�L���X��y��'n�r�'��֕Ya�ƥ���i��f�f���O`��O��$���I��&����T�9�y��o�J@���IQ�	�(���I.5D���柜��ҟm#�428|Bo�=),��FB�ߟL�����ʋ}��'��'�ڼ[S��V2�$1�'� M��7\��c�|����K`� �����Id���G2���*˚<d�`ReCS&�?�$���O�OV���O�{�*M�S���9�`8�Ri �) =���$&L���OJ��O�����K�m�C`�3.��R�`ӷS����?���䓏?���,��9���q���r��OG�p��c4<��� ��<Y���?����8����<j���2&y�Y�GmĶf�2��F��ޟ���a�ޟ���'~/v�]~r��5��p��C��3D��?����?ѧ��<��A�������	Ο�A5��Qb���DR�qִ�v��I�	ӟ�I�gD��	_�?��Qb��`	Ńŧ\��o�O����1OT�D�Q��ݟ��ҟh8,O<	�G�Z`M2���g��L\����'���'%ze:�'��'~��0�TJ�`oN��T QV�t�������	�M���?����?�7�x��' �a��̠f1`! 3��K�\��4O�5�4�'a�'��'!���ҟ��:{����S�"5C�j�WY���'�r�'�rE+�I�͓4�@`��5V"�L�Kͧ����I@�	2aVp�	�Y���I�x�Iܟp�W�W���a`�l�p6̊˟���ӟx�N<����?yL>����W�-�O�=���u���L�!y�d	*1��$�O���Oj�?V<��h	.E�!Ԉ٨E �������?�����?��]��X��	�e�n�Q�޴9T��*��<� ��<���?!���f:�� 8s,d��l Eˀ,�C\ ���?IK>���?Ap#���?�	� �It�� J'�e�͈O�If%�.�y"�'�b�'��O8���?�6,����k�=Z��r�����?�����<q�����ڔA`�U����q#�f1I�'J �y��'�꧀?A��y��4␱�V��u��XHD���'��Iӟ��?Is`R�0p���M[�D������?G�ܸ�?����?����?����?���?�F	� �@��%��k:��2(�?����k���S4K������bĦm�W�?h�$�X��
ɟ,����M���?A���?1�_���O�Lh�_���p�IS����
�:�<ء���O'OL�y��'�N�� �E�h�b%��ꎣr�����'���'�2�'��v�$�'�D�*����$��t��N� Z
LP��D��ށ��5O*���Ov�$B*q�%��ˍ�|���T�\�%U���O�$�O��$�|z����b�v�qR�s�5
֧�8b���H>�!HR�NP��?����?)Ο\(s⇐=Ä$�w�ͥU��)ct�'�듀?����?����'�61*�mE�R,���ӁK�إ32O�q���-�y��'�2�'��U>���28�2lY���(4Z4��B�z�@9��ן��	۟$���I[y�s_�Ő�O,�� `Q��N3�����E��8h,�
k;����>=~D�!Hц������4 �`\��E��d�@�#��٦E�5�	ןx�I�D&���O����d����kN�eȎ4p�ƉF ъ'��O����O��O���i��Q�Q�}����+͛I�S���-Lz�e�;!U�l���>+E��z�'��m}��dΑa����ʉz�`�!=̘SB��qP!�Eq$��rU��~E��+��~0���$A�X�I�J��R�P���Uk �;')HB:fⲍ�/"�T��p��n݆��r��N�F��r�V.��K�E�c�J��5�5���R�v���zȖ���]�C<Ȥз,�0y�މX�bڢC�ĘOsߪ]�T	�0YH���FtU �q� �M1!�ET�^d@��% C1��A����^<1�2��( 1�,O�d�Ob��P���'F_\H#7�ߟ�9f�.����N�fH1;�!E��#?9���% *�r����N ܑ��Ov��cY�/�I��#N�p����X�R�'v�O7L����+��qr����IXL�(����t�2k��<��@����3Z���Si?A�8�ڈ�S��P��2Ԩt��Ʉ\�dU�O2��:���O@7-.z�R�D�iO�����U#9~�a��,M#�e��\�Ʊ��Q�ʧ�ħ$��a��I�i/bq:@�qVh��'��2�Mމ�n���%#��h���ڽX�DD���I��n�V��'��O���6?%?�' ��B�	9f�t��p����
�'� �z'	��K��J y.\���MQ�O�����OZ�o�j�����~lv��'�R�'wj	��+xӲ�d�O���<A޴;��)��I�Zhyv��ҜBq�� ��>5v9�$ 	2'ǉ��'<0y��+U hQ��r���$Oݬ�F�߯^Ў��	�?���/���g��ؑI%�<��0&۩Zfn��OΕ`�'�2���H-8�,̦>� ��5(����V"O��0�"М\���%�I���#��OEzʟ`�ZP����]<���u ɮ>%����&V!<�v�'�"�'/��ޟ4��؟����1�J	1��6Xˈ�r�)M�LC����>�ì�c`X eg�7v�i�@;�5H)��`Vx�q���`)(t���
Hq<6��jt��;���&[���`�صF�\d�	�M����d�O����·#� �"�*�Q��$�5�qO��=%?�� ��]iXaz!	˴VXpiP�8}�uӒ�$�<���'J.���'<�i~��r)].B8	�a��Ȉ0��� /�	������� 5c��h���'��.��aV5isEWM+z��c2W����A�EՆ�"����*�@i��{��X�ˡ4��9�䏋8�t�F~b�Ƃ�?�V{�v�'��	8dՓ���_��5��Ι ����O�⟢}r��p�m8����������{?Ɉ��i�Yk����H�� F� CB�(�oȻ�P�'^(쀀�|�����O8˧����M+�A�#�l9����5ĴS�g�b "��	9�0hH�"�T>A$>�0�� -֥���AtD����l�>�2Ș�G-��I>E�d,L"<Hr���OP�x���������b�'��'��>-I�g�y%6e���݉27Z8XO=}B�'{a{��M�>��� h�q��ax�fK��O&)E�܈	:HՀ�S�o�ެ�-��Q�V��I۟0��;zK,Eݴ�?!���?�/OG�~�̈����4o�2�1�"�6��J�T���	.Q��̳O�-zo�����2u�OP�v�'4�`	5"�'|H�����<�D2N<Y��������	�2���uj�0B���a���K�C�I� J�\�$�d�!��HNs`����HO>�!��3���+7̈+8Ēd`F�C�-�.h8�4�?����?I-O����OF��{�6�PLI�"m�@��["�,�a����M� �Ժ�&�r����#g�R��1��'�x`��4P���VG t�.�P @ץ-�,� �O@iɔm4�<��3/�"!p"O��iq�Z]04"�E��h�S�>��d�9pF���'��i���( K�(rgA
�o�*�� �<���?��x�������A�Ao� ����K'�Tx�W!��� BÇ�p0"?�#�)/�J��FL,R�A�`G矴��EW�.{�l�qD��g  A;p�ɞ�~��'p�O۪u�r��M�#�O�j�D�H���ɽZ�ތ: ˾	�6 q�5����J?iBg���qFA g�LCv&ʸ&3�	�F=�-+�4�?y�����2޴�M[�២l�V;��@H���  ��-��>������|BM\���MO�~�<�A@�BZ��^r�<E��
<Y����%vI��uhJ*���V��'\��Jb?��ԋA�p���Y����a7}��' a{j�]"t�3�AB�=f�oW��Oh4F��I�O��z�M�}�@�5�Y�����O���"\xmZ؟���ޟ������'�� ��6��=5yX�Z� �a�IL:��r'�uR��P��\;��D�7�'Z��ۓl�r�ᔃ�$��완 
�E�N)$���3��O���Ӱ:�,(ei)f�v�Hr��V!�ĖHW�B��i��C�u�J@�'c�#=E�t��mvȘ�N����ܢtA8&:�u0�Fg�����OJ�D�<9��?)�O��Pش�d���$�I���Z�͑��F���	Hq�7-O�R�`u�Qm+�ܮP��u��-��m�q����?֖���N�m��i�'X�H���1��,����� ����'J��+���5eO�Y��悴��M�@H�}�� �6��O��`�j����P%5�9�cjؑ	hͻ�VIyR�'M2�'5��Z�'D1O뮛�cӸ���o��V�R]��^�}�� ��8ҧt��$R����=�����h�F~���?Y����.���5�%ogri2S���y�(�M:8���Eea5�1@D �p?���Odp�Q�S1Jr�aĨ�0-�H`��>�'�֡3a���'���'�Fo�=:l��Gݖ=�V���gԦ�F��^�D5�|&���A ��r�T$��ˍ56��R��>qU��m��H�  �C�9�a���#S�rt��P��!��O.c�"}�`�. ��@�m�:G0|/�B�<�cN�"�0�;Pa��Q>��`,�|�'��~BTH��m��X� �q��QR���8D���'GB̗�}�~7��O����O���MC�D�/q69��X_Zq�e&Rw�I Fv��D@7�b�ؗ�
7xuX��B<f�'�4���X��[d"S�8�-���z�&�l(Ѕ�O��dS�uBuᓡP{��Ъ:z�!� �l���iw$��Oc�- 3�	�}����D����p���AZ��t��@�a��D(�l��TJ�m�П���џ�'H��'&�1o�v���%������ �g���K`���?�h�򦹉��H!����_�	[�b] ����� 7�6ˑ�~�>���/E$JU�i0����*C��;nc��E2J���v	܄4p,B�I�J礝#Ҭ�Y�	d��3F ��'L���d n%H7瘺��|��eդ\�!���c��k�(S�x�tE.��xO� KZ^xX��c�;PF���q3�L�PƆT�j?�BQ��Em���� $ԂW�}����ȓ ���D�3T���.���5��dj����C`JI`�eԹ,kRɄ�%jD��ȠH���&��x���ȓ{@��%#
/����4�ʨ ON���.�J]ڱ�W6&^����8n*��ȓ����G%V�"i����P��ȓ[0��0���]��8:2I�o4��ȓr�6�X�!�3^�L �3ʉ1ye���T�|#�K>"��J֨Gdm��c�L����z24ēף^�x�D���S�? �KPDL1qU��iGJ�fl���5"O�����t
�ᅌJ�sU⸱�"Ox��Ɔ�9BQ����\-xJ�@��"OT�z��?���?3!&�Q&"O6���a�='j@QR�K�G$�h"O�0�hR	ݰ�k���4`T�v"O�`�W����&p��mء0�V�" "O��
��C.<h���k����U"O�TNG�	7�h�D� r�Z�C"OR)x���(Y�t�:q#�/���"O$qqsD�/�1���	���Mؤ"O�(Ҋ�l\HI��b�0���J�"O`��uB�K�T[�l*O@��	D"O@M���%rC��+�뎼rKnX�2"OP�����PgL�Rdk�0r!�C"ORQ�5$�Zk�""�O�6&�Ҧ"O�pH1�P�!jvt	��K�.ڍ�"O.��b�/�&` �ϞMl69�!"O�I��f;::�Y�0:�v!��C�h�&m��4�\�if�՟
_!�dԵK�Be`4��n�ZdB1���t�!򄔤Kn =�P��)��
f H�!�@TI�)O�Y0�L0M�b"O�dd��6/�!��K�	�P,Q�"O��Si��oZ昪宆�,�{�"O"@�ǒQ$�z��;h���"O(�����6ö��"�6S���Q"Ot���Z�P���"႘h����u"O�0`A&Mv�m,%𐹄Y��y2���X{0�2�΁.,"��Қ�yڤOu�D�fl��P����h�#�!�/2~�� �&D< ��3�Gͬr�!�d�_�@��l@8�d���p7!�De���*���(z��T@�3�!�-�]�2�R<E�	j����E!��/&�Z���/�0|.�QpU.�`�!���~�ʌ0A�.l| "c˺]�!�D��`���4� 	/
��s�[�w�!��r�"U�7�ߙ�@u���.�!��d�L�zӊP"-��:���!���LIا�ZțR�5 !�)ʼ�Ic�Ӧ���o���JC�ɗq��Qץ�i����W�!_6C�	q~|��P
��5��cd��j��C�	,4��l �lb<yG��yEB��2yH$�ӶBR>0�|�y�kߜ�4C�I >o�M�!g�,�@�aWK19��B�6�xEu�$�2fE�"q��B�		P�D3�G�+�&$p�|�B�	�o�0=Q�&��"��J�fB��_��<k�oE�C�I �f
�S��B�	�M2`�p�l��S��Y�*�R�"C�I2/d4u�^ξ��&(Y�c6(C�I�xi�}�QgԿ]h��2�Y�N� C�	�>B�0v�L,^:de)��״W""B�I�Rp ����]���ՃoMB��9{CB�c �_�a�H�2�R�@�C�	+���Z�iO�i2A�նa=�C�:q��ة��7$�T��S��I�C�I?u����I���a�4�g�C�I`EA�OFk�a#RbLx�|���"1�8R�{"@Cl�u�G��`�,�[����y��+ww���aI�^��J%���ׄ'�p���
5��S+N�<P5	��9�b2���W��D�6Nq��+L>� ��ҡ���|ѻg��yɾ�)�!^@1�ꗽz��١�۬#��3X���0#�2x~��؄G�0F�!�O�@[�ϧc���O��0G{�5��ɍ�;p �fF˅.�؈���br��s�ob�H����H��faJwܽ���P�M�B����a�D�"�:4�M3�"��i��Q�j��(@����d�aكnfٰE�Ch� ���`�Aq#�E%}~]�v��?2�a��02xNd��V�j���C��]�{C4)sgD&yz�?��$m�ig�e3��G�)2)C�0<)��;���X��fh��ƌ�$S�8�PA�^�tLR��	iƲM
B����e���Rh��s���Vc��V(�A	G��a�'̱ "̓���O���
����$��x��L�oj%Y�M�yuX�A!e/ش�v��'��{��c�x����׬�['G��Y�'�nT��/�"lc�A�=Y.���M��l��I�! ���5�e8!��M�ƅ�j��� �D?�O�5�(;ۈ�Su�:����`�V�f���<SgH-q#[

��A�nG�zی�35�UP�'y�4�9�(3�Q�'LD3>��s�ɦ1��Y�aڢi�(�ٓX�sd��+%I8,2�c\��N�(T�^�K�Сj�D�#s?ʹsP)ĊC7�q�D���?)"��d�w��tk+SX�y��N�)���;L�2�b�@�e��0��M�$�*R���N+�`� T�g�F)�Ԉ@��N�*�+3&�.��L�Dʐ�'�� {t��]	<�PWb��I���y��O��r�i�9��m�N�VD�5��d���h�CQئq��4�;�4�HţR�_�X\��E��x�M��I�>�2Y�qA�ϐb��	�w�ʼ596lq&��Dq��'������B �E¥P*�U� U,n���"��)h�#>���o����-�<y�mˣR$��K�]ڲ�HT�N3X�����.^����dC�Ъu�,f���YVdsP�d �Y/��2FɌ���$��r�@�kY&��''b�	@�O!v�Ev<�Ą�}Vxz�gF�?Zr���/�Mԧkp�����m��A�<�;=PJ�)���ć�{Z�+pʁ
Lp8�b��D:,t�~�N���U(��@Ϩ�+�a�MS4	�
�b?�I�	��@r�[x�џ�Z�_\������v�nP�Uh#�6������%}B(C�vj��P��<N�����E.���u�	f��ɇ��6'�|l�tg�S�:XJu��#��?��E�+OD��D+�	.��j̎�������y��ì0�ȕc1�
w�8}��/ ��D�?�Ny�{��	!Y)����!��?���7쁣�!�dL�{}H��bȐ l~�Ks���!�DB�2�uiq��!D���̔�n�!�$�=�lq2�H�.스աĨ�!��Ԩ`���Q�GE�g=PK7.�fA��0R*԰DO�,D��Ǚ@�!�7��ض� ��
�yb��9� ��!��Uq)c-<^I������6��H���Y u6F}*O|�ɒ
���P�ڇlL�J:y����䀃a�XQ�Q�?A�&��k?��p��/�������<��㞀	�0���	L���<iF�ӏU���f�W9m� ����@Y̓m����M@�d�:�H긟`�f(Ek�c�iǨ
�� @dΓ�%���c&JA1Ѱ��ƓO-6,��鄡O���'���< `I҄>�D��ʑʟ\�c��I!.�C	Ġ���Ҟ�,��1��$i�m�P���%�T?!�C�/U��@RN�"p2L�Ï�]�e�B�!�2<y�ä2;��ϓ.Q��p2��!v>X:K>!p犟o����?]^���aX������:y������@�Pᣂ' �ޙ���N8qȼ𥊂�6+2O]��������]��yBKX�o(<Xw��( %�Ȼ7D,��PBh�o]�]J|-+��B������z�ҩ���e�P����6��as� �i4r`��D54�0�e�*m@���wV�#�DY-����Oֹ{W =P_\,�Q+nD��'�M�'Jʼ{��A�2�,ybυ("��@P��J(<�� ۱Mu���&(�7!rF����A?R��	��H�i�@]k�gU�+��+��N}���樔�$xT����S��Q�~�xI��-c�AR�/�!n��x2�V6�-2��<���$�/����3�`8uDB�3z(�{ :OJ�!���RE&�)�'R=��%��O����
Ω;�
 ���4B��Q�O�   � m�
��Ư�0X�R�5GA�'a�^�[��I�-(cOD�,�;�<f�Tu�L�\��Y���q�D�o�\D�@�!4@�G�XzT �v�D&,�u� �C�̚�>}$��`���3^����1aO>�@d"v��Qar"G)uW�  ӓ6����9�ʠzŦ]�oC 	)�		�M�B��/)Rf�%�f�R��'d�9��S�]&r�/������ˀi�T(h��R"�p<i�⃒,�!�,O��AJr��:��ϊ�L�Mpu(\Nj�ɈyR��)YBtؙ��@�Od�u�/�4Y[�Ũ����I�H<y.@"j����͹j3�q��f+���M_\a��)!pM��l989>��4E5�Ԙ�OvhD��O� �8�Qi��l�QRj��1l��`���6���� �$�T��ցx���'�z���� }�9h"�[�I��T��4V�r�R��"I ���ڒ{�0�� P ���P���9F�!�Ǭ0K	��+W�
c��VU7A�Xa��'ꀔidJ�%V��&��Dy:��ϓ'P��v��F|0���n�F �|N|ˣ�N�,��#(ç��' u�Īĵ%�?�����c�����L�x���J�M3�	���v�<����[�c�Q>-��@��q`�i���/P�!���Z0���s�t�����,���k5.�rp���7I8|��B��y̓I9~��r���t�a��5b��$W/	NJ�D�BF&D��g�1���SS
ǆ�(�N�0!xN�:�M}��I����n��!M|�	�g|��ۄ!2o@tl���7�B䉔7I����oB�s6���҂�(��.�*��;/(�܅�ɇQKP�{T�M�&��/����#?�O����*�j�"��DN��iY�7^+#�?�HH��'�<�S���� ����!�TC��D�i�I
gnڳ7�\�?�A�v��`Ƶ"�u���I�y�Df��lDlنXԳ��^yJ1KȕFȂqp�P�"~Γ?
�(���N�R���>*�R��ȓ{|���	�^'&��F)�!b�-�)������+h�2ϓ^\�m���4Z;�
vO��ilP��d�<g�����x�HP�&�
����S'�&(��ʤ�$4�P����tr��!+Y�7f0(P�o&h�՘�oY�'%����D��6R�d��Hǩ+c�u ��'�y�o@��T�6j��^'��B���p�� q��j���M�"~���(��[���)E�T�� k�C�I�5�rt��*0<̀���D-��Wk�H��)����=�6�Y�[Oh9cCC�A�4��d7D�p��Ι><�Z$�'t���	 �6D� s[^���C��đg��I��J5D�p(���t�QҴ^��9�v+-D��Y��o\��B��h�ץ/D���F��h�<�����t�r���!D�4��N�`:�v��D� ;`�?D��+��(�qf]=o�X� ��0D��1�'�2ͼ}ZG�,k�:�!�(5D��!��%Ect�S�^�7<��.4D�8CEC�(����j��a�T�1D�� A�}R(�sG�]D�����)D���ݢ)rq�P��!�I�gG(D�`��'j��)4�7C����a$D�$*G�Q�V�ܝ��b��$+`q[� D��P�)��x ����+5�L9��0D�P��'U~z`@J��>��)���1D����<&H��b��B2S�q��l,D��,�	a�US�Eڳnl��&7D�d�p���e���ee[�h,���$#D�<�Rj�'�"�3��_�0 �a�� D��2�j��B{\5��S1J�*�e�?D���2n�Y���gP:<\Q��.D�<�D$�8A�B��v/O�H�
HbGB*D����/if��D��.q\�i(D���'R�	�$E�f�1j�A��	&D�<�����}-�<bR�ʲ~�0�;D��y��&�ux��J�Q}����9D�<���� D�2KͿf���F#D�0�b�ٱX�Ψ�v�
�?V�a
��:O|�BS��-��d�w�l���	��O�^+ ���'�5S����Ղ�+�yR�Y�R0��$0���yB�Ȭo"h���n�1'���4Aʟ�y2�	�{���rG��T*d4{T�.�y���`琑Q���MU�(3����yB�ܼ0 �B`�]�F}L��ւߢ�y��)A�l�#�+[#CC�)����y"�]�<�<�j�h�j t�H�e۫�y
� ���`E��p��RnU�nP<�'"O��i1���M]��O<>�*8"O��).�6PJx��.�4?�^���"O�BT/K	u�mY5��y"�"O� � o�U��*�͚�A���v"O��� Ce
���L�w���H�"O4� �V!�:h(�S�r�����"O���� Jc��mr��Ǽ!�xq"O� ��ŀ:1�l�+��|���
�"O��s�n���k$��H����"On9�P�@%{� @�Qɚ�-��\
T"O`	������5IY&Y�Z��s"O��C��Q"D���f�D#C��dc�"O�l1%�ܹm�T�4G��j%�u"O�$��lˆY����F|c25)�"O#�7F�̔7�D�b��e�e"O����D�f�S!�G���i( "O<ݙ�lïi[V�ȴ	N2���3"O�0��ܪ@M�U�!�ų`���v"Oj�Xg�֠~zP��͞���"Ol�H3 �)�$�0@_$29P"O�\+@-����iH��Ԋ+��(��"On|��/^Ү@� ��$���"Otq#�)Ў�%��h�dM g�"�y�&�h� `����t��1v�d��'Pl0qw�N�^�Ge�MI@��ʓ��Kш�THuk�����1j��7�Xc(�Ri�6�n0�ȓDpZ����o� ��/�(C%�-�ȓ7�e��Uf��q�N�	<KjM��/~^|�'���,�����2���|ˀ�p��� r�:)+� ĝ�ȓ|8<��V���Y���N��vq���ȜE�d$iˡ��t�8d����q൉���Pȡƌ2\5�ȓs ���WZ���D%Y������Q8��Zhғ@�8J�i��iP������,�%g:,ؤ}2�:D�pV�F3Y����.Ф^3L�ළ3D�$A0Ɯ5D���`D��
T�co2D����W&�<쉳��f&�%P�.0D�;�O��I���`OK�&��]х+D�@����{�N��`L�窹B�E/D�| t���r�61#rOLRֲ�S�-,D�(x���7b��@�JIukȁ�n*D���%�W�t]yW�ф��	�)(D�P(���^�p�Y� Ši��IA�&O�����@�a��0@J�3c�����_�je�� ����d׿���R�A��T�(y�'�% �H�S�OЈ�ّ�B�و�
�H�f���'�nT;A�B4/t.������(�\�q�y2���,�L��%�r�����3�	��JC��!�b!QtI�'�����+ُEލP� A����Pi�y#&AêP-S�M�2��xb��	�Z�@x��*<���ė+xB,x��:D���T�Δ}5�	���Mv^Tk��7D������*D�F,�jg4D�D���ܖJz��k�� #j�(�sCD0D��ZW�2��Ʌɀ�(���$"D�<H�Ӓh���nTc:���+D�4��\�(�P����43��M*D��:A%B )��;5&�@�����'D�����%Q�UB��u���'&D�X9vA(l�6�I���KBָ�3�!D�� �iʷ�:}����£��h���rR"O�)���7|�с0�N�%�@�"O���b�I<Q�*`C��*ZJ΍���O��:�O����e�'dp�b#�!#5Ջ��O�<Gzʟ9�Š�>Y�dK�v�T�jh�W`N����Xi�<�f�X�3�l�����#d�ݐ�^���s&$��B�DS<������͕���Y�%�S]Ұ����3��1� �bĂ~x���7��qF �`̒M�XIwdK/��Axb���C�<�G qO��2�%��?9Pأ=�� sl[O2�L+�I�--�e��͍"�J���/Kr4O6�x��O�r��i갭�lr���U���,OX�	��:$�\��CZ ��mIԉŻ)��I;]�%%�#�0=Q�@�L���r3��;@6�j��%��Ȁg�w��	���`�<R�ʟNأ��E�X�f�jg�f�v8w
O��p��׈9t������79�ݳ�
���0=�HȻ\X��h�_�f?F��G���-2d�^�J�
��eRf8�|�����;e*�(��K�	|%��4� K%��TzJ|3�N�x�1OJ} 7�^�8/�;E����aJ��$@�e>䙓JY7�H�y!H�!3.�X�Ɛ��J���\�ė3rB(�?�%X�����o�\t��{�lY���D��'O�|��A��[����`I�)��L;��� ����*N�i�f�ܔ�萄�I,2�Z�\$:������W�0C�	�-�H���!,wܵ2#�[�V���'-̉�%bA��B'i�}:�CD�Z:=`�V;��H#D�0O(]I��2z�!�'� 5{t%�#n�R�d�3�Q�l	�U'F����'��T
#N��Kb�p*�Gs�Dˊy��� q�m���<<"��_(��	�{�xy
@F����,ޒmZ�h@ �T�	ɮT�Ra�Eth;���&DBL���Z%m�F�kU�'�n9Ta:��-�`�U�a��}����F�q�!�"MV�zZc�6u!�N��D�t=���,�J�	�'�K'oS�
u���K嶝*f�_j8�()�a×o�|��r���?)���P+�O��覈E��p�
\�@p�x�>�T�6�
0Q����гl�d��$\��r��r�j�Xa�'b��
�MT~�����l:��ɋ��K2LH���4'o.���GQm��)��]��˟�hZ�pK������?�R�9_80�D���R$�)�A�� T��������*k��6e����qu��%G�����<!�F�ztf=,O��]z� `c�Ȋ�`��9�E�8N�|B�	�䘻6�N�M��P�&s2X��t��D��M�i���(z�6h�Fኜ���bu��	yf�6ƙ�am̭)�eA�.iLp�jV��p<1��@�E!��3Ł_��֍s�mH�x��	��ğCK�5s��R~����L��Xf��1ro��ץBn�=�G��j�>30o�A� u�e�V�d�V@���my�I1RE�'"��'q�iqİ:f �{s"C�c��*u�^�:�@�g��0?�R)��1 E{��	�N鳢���iMJ@�G
�2�k*�ș��u�d9�O����(�JDdÏg� k�H+=`4sU
OD$ ��J���X7�K6t��e��0+�UKt�'��D�8Ol��'ά���-�a��,OBQ����$>~�(��J9Y!`���'������jed���O���!��aL=X_�<KW"����	�œ�o��Օ'�R���/7�ax�� (i����h�<3�4��c9��9�hx��2�P!e��4��c���7�L��i�:<� nװ$� ��r�� ;r�da��3$��J������Ѣʺn4#� �9*ĩx�ǘ+^�����JY#R���B���M�OM�1�w�J<�P�F�{@�M�"��{̡8�'��UH�BO,�P��0,_b��:��V�dnt6��M�S	��>{�,�S)�+}���A��P�3=~좄��Z�f������{I���	�bf������;ɘ3��מ��D���:9�(����$�����T~�����0���'�"�Y!/_-�'� h;�_5�4�3�/H� ���RL>1�'X�`O��P���3��T'E�	>5	� �%<�i81ǅ�*�tH��:cW�݈�#2=�\��z��9��GF���*co�N��V͘1gP%(�o׈rv�Q�pț U�p IX�b���)ec�.�<���j@gƪ6�� U.5�B�Yb ��e��պ��$D��0��\�|,�u���J�Ҹ�f^sLu��FQ�I/�p����f�ra�M�8��t���'
��I/��L20�!4����J�#Sj�!;��7<O���B��ēB��fE�1�����,�f-١-:�$�Y�mŒ^�Nm��d��<�`I�Q�F�<I�MB�e����Pe^�Q�>�(T��s�I�>�*PZ�,)��ͧJ3����^�r��� -C/��Q�]��L�F��*fXpA���o��h���"f�'g�h�B��~F���#�H��T�wN���1ƨ�x�ES7�R�S��l	'H@C��h�]wT��7��8�Ũ!�~�@GI_��t��O@9S@i^3v�~�Ѵhvɱ˒1�)�6��i�Bh[6�K�E�"
s����#��3����*?�7��`>�9K �F�K����f�C8��j�$�[U.��bK��'�����\�-�a�I�@��i��N-�N����qZ���᏶�`�1��$�S�? �@'�0!�*�׏T�s��>	@�N�.���bѳBh�`"H@� 4z0�&��DO�n�x0�26�*�!"	�E9�O���UKZ�~��thЏL>Z�>�P� ��5�ꓢ\�f=H���%O@��'����C��]���<e�d���J9���W�_B�Cቒ,2,� ��@&H����;%,�� S��b�O�(G��%_�j��)b���r��>���8~l�]�v�?]�M#q�w8���rʅ[|du�3�ԉG^<�0�N�İ��h�#�FΔgc\X��D�j�q�d��8&��l9��'�	
Q	�)�ʐ�耑"^��bM<!��!cż��b�* 3AHH)rA�'�R�Z�d�%~�|����!!R��e�CvC�	�l*�p�	M�d���aFg��h*�ʢ�N)�EHң�?��2Y�8�&C�ZU�S弃g	J<5�0����{�M��� YH<��T.�Li �BN[�������7<=�'>f`I�! /�z�ȡ��	MdTɋdc�P�F2��D٩7�,ȘwC��q�����I3%'���$k�-yz���B��L� ��'䉎L�\�!�(�]�35B�8��@�8"�0�E�2�p<Ib�^7
S�}�L�;#�>!D'C�$��7�V|@&�^F�,��Bi��1O�t����b��R�j�`h2LT��y2B���њ'�*U��!i"�M1����Dh	�y�r�P��O��}*��� �������i�6��9>���y2�\�Rl���O���\H�m� 	��������~jA)ۥZ����J/~����G�Vџ�"v�:�|I�	܎�Z��r�4O�m!�-�0�Z9hQ+ہ�y"D<:�j�htBуwܸ������M���Z��^:p�x���i��L�4�N�Os��C��F�~��N<���4��G匹������Va�^S�E"��$ng�q�U���R/;96Q{��'6h����١A�s����	�H~�C���;�ظ�r�Qs���烀}k��R$�,4��2��;8|`�C��r��J�>ғ�\9�:8��?�hvB�8��Kg �4>α&�=D�0��nT�V|B��R0+*�U���OV�+E'2(e0%'�"~�GB�=7bE��l8h<�5(���yB��H�X=��gQ4_sR\y�ٔ�y"�ǜ }�8C� Wd0��tE���yb�U�B���qE��R�E��
L��y�#Z"3�3Q�_�U����aT*�y���IY�Lځ�_B!L+U��y"��N;:xa�@��CН�c+���y���!�J����sٜ �"�2�y®��-����;1�� -�y�e�z:���tƛ�0��܉�b��y�`O�R����>��$7�E��y�)ܐ�V\���P$ e�}Cv���y?:��)B�gS$#j���J�?�y�⎞l& 5�օ;���p����y�&L�m��ՙP␄c��]�p�<�yR��J�F$��n<T Мh�g��y��OdC��Qφ�#�
�ZS��y�ʔ �d��é
�@íG��y"��o��� ����1��L��G��y�@�POԍ�b�%mBYEf��y��ڨ٠�y�I� ���w�@&�yR��%�f*�> ���Qh���y�E��'R�����u/B�0�`��y�Āg"E�2f��m��#�D���yRX�h��mDt9���ا�y�*��q�	� �:d�w���y��̆*Іmq��Ϊ,������y�N�-���B�5d�ي����y"�	1��t�,*�d26ͫ�y�!�$w��e�G? _��I����y���piʝS���)������'�yR$�32B�どȧ+1ZhÅ����y�L�+�`!qO�0*(�Dk%����y��̥eX�D����k� 4�W��y��Ӱl�r�I���^T���`�L=�y�,�8%(�գ2��4i����[,�y
� ���C �-%4Ĳ�̍����r"OP�Z��GL�1�f�Z��f�k�"O6�����n�́zcj�#��U3"O��[wN$H#�RԆ�c�"OLSc��=�h�WeV�%#&"OD�Y�*��!�f��Lu�H��2"O^�UGV�0�ٰ�΅��P��"O���"����m��_-bؚ`"Ol,G&4G�V�ٲb�2OKX�hD"O�Ǆ(;��`B�ጭE���"O�t��	5}�d� �(�dZu"O����J�4x�Lc�߇@k����"OX����1}T������.6gT ��"O5��N1j�3c��H5as"O���/�*Lؘ��Cđ|����"O$]�p$W:r��M���ԠD�^��"O)�	s��p����9�����"OИ���#R�81x��@�$�2��"OZ�ك,��2)�@I�+*�"O2Y���Y2m�Ɖ�f��p|� "O�!�4��6��뱎ڡDL���"OPwрbP.p�k'*��w�F��ȓ�,QX�K�zTł�M��$.���ȓSE�U0V�_.G�0�����&E^,�ȓ#6��A&M/nd� U�MFΩ�ʓp��D:F"D��mk��نS��B��g�F�2ȋ g % �ט-�B�IUN,��3�wo4e>B�I�q\�0[ү��ތS�o1�fB�	:v�H(�GB�Q��;���;ԜB�IE�&��F��6o~h���%pB�.h����1˒�#�,x���ԍ;�PB�	3?��сM
�h�e��C6BB�ɋs����>e��H5)�?nDB�	�P�|���LY$+y�})¢�2y�0B�I�z� `�p�-̚	x����B�.7�D�q��UfH�A��l�2(��B�ɘML�|���#O���c͛u��B䉠�<�#c*��;��Q��_w�B�	�w��i1a�/�|YR�F�B�4V��S%&o����s�B+a��B�46� 4Cr�Щe��TKT�[?PB䉚,Kp�h��4W~D�R(��NB�	 vsh�7jݶ|���"ֺVc`C�"F&Px����l���a!S�"�4C�I�c>V�ha�K�-�d�)�"�H��C䉓+�H"2N9H>�p��*XjC�I3<܆`H��ۙ,$Xѥ/Ȑ8g�B��nek��֠�` �u�o�zC�ɖZ.�0�ԥ\qX��&Ş>�C�Ie�� ��/Tz@�B�
~3�B�-z&�����M�j�p���o�B�I*j}����
�l�"W ��m�.B��+z�	�����H��!_��B�	�s�I �K�7P���У@ �B�I�j帲$�y�J�ZEmO�9�~B��I���CY0P�*�@Ц9wB䉛
�} ����,�R�1�#r/�C�I,�� �2�U�s*��Q��3rC�?U������O;@�DAb�[���B�I{L��"U�.��}J0�W0`��B�ɝ<zn�0���Sgn��B�I��Y��@�-�T��0'�C�I!I��ԣFZ�N0xi���&��B�)� �U��i�턡a�H��HѰ"O�\�0D[��"W�޾&:���"OL��SoȦbciG�#:��i�"OZ�z�炉uKL ��Aץx���"O|�#��oF��&�ws�+�"O>��gGX��Gd� R���"O��X��̞hd(J@�;.`�E"O6](�P�<8���Wh��&X�*"O8�6`Y8�Ωq�f�%��"OT��'Ü9NaQ`�NӲ�a�"Ojiy2��6( ��1����"OPDåŒ�zl`,9P�C�C�I��"OH���"}`�q4�\GL���"O"�5%�H��j�FI	�f}8""O^X2��F�c?��ef��Dm,�2�"O��XQe�6ZL"�H��8b&0�q"O�͢�j�^?�J�9�r��1"O �sT`K.�j]�����좝�B"OlT��j��P���u+���xݫ�"O�(��Ɔ1���*0Nl�(�R�"O���_�4�%s'K%M��1�"OY�#�i �ĹG
��.J�݀�"O�����f@D�fI'fR<Yӓ"O:4I���c��6B��RC ٺ�"O��B������@�F\��"O^�+�#�u⽣��E9C찙d"O8T:�e�'��d"��'X 2$"O�z�K���pNԇ/�N���"OV����
��m��-,�b�"O	3���w����9&�3"O^$9�oV)0��r��6A�lE�"O<HPmءq7)�@��'����"O:9{1�\-il�e�eIV��!���:D�@B�
�&��K�9D`�:D�X32⍄q�FP�VI՞WbXR'7D��7Ή�b�؄nȏfd�Ջ�f4D�\��E1Ʉe���S�'�^�c�1D�2`��.5y^8{� M�>T0Ļ1D��b0��3MPH����7�!g�3D���VI:2�252��\�kbB����5D����&�d�f)�1%�h���8D���Sǐ�a�z{�"�<x���`C6D��2l���d�I�+�QB�M�p�5D�L�ADE������R=t	z��'D���Y5
 &U�&L >C.�x��"D��+��E'ƹ+���9B��� D��)F�?"��QgР=��(5�=D��"�M�������>8����d=D��(%�i�v<�3���df���K!D��`���"4�*�m�v	f�>D����A�i��4&�cN�u�?D�8�/� ��h;4b��(�v�:D�,�+�%X��ઃ�ι#�,P4#D��+�/���)�O�w�V#�� D�8")������M��!$D����L?_P�Õ$/
.��*,D�h��
M�jŒtA��׵d&�t�@`$D�(��D2@x|�����9T��-��#D���aR"�t����8��e���"D���I7p��"E�Y��i�##D� rV.
�=�52��	��9��l5D��E̜�j(Vh�Ц�1y0�Š2�?D�p��쁐{�BI��J+���r��>D��yA���"��|�g���1��Ybk0��0|� ��Q�K= ;�و�g�O�N$�"O|�q���!DO a2fE�5F�H� "OF�i'	T�`�y�Q�����R"O�$A�Z�8���T����"OL�aa��9M�aɦ$�<y|�""Op4C��ү�������S��:�"O���T���q���%#{|T�&"O8`*5·r-�5��;x��"OfͱpO�&(Ӳ�	#��� Y�`#"Of���83�
���T e���q"Oh�;�,O��6�R"	�,Jʞ�j#"OL��Gl�;��BA�ׂl�����"O�	�(�8��z�/kML{A"O�ĒDէ�L�k1*ӴpDq�2"OС+�O8-\�I���\6�X�$"O�}r%S�bߖ5:�F�U \�r�"O��4��}�L�J������"O��%.�C.Ԑ��L�'`�L��"O����I�e��paM�̀��"O��:�c�gՁ�I ~Ĩ�pu"O�}b�Ԙh�@��R썍L�:u�7"O(��$��d�N� E���DX�"O��K�n-Wx�H�'��>�D�B�"OTU��Ta����˾+}���4"O���7"��F��r���?']P��"O杂W���"բ�r�CL6FР�"OH]J�/�,�Ρ��]�!/>� �"OZ��a/��P�6(���0� ��"O�8��ޜ;��01P�.2��k4"O�i�cC9���
S��7W�e�2"O2=���)$�����mD-)�U�@"O>U���z���5��0Q&`h�"O^UBc�9/:���:��(��"O��qԆW ';0\��D˂@����G"O����p�ʱ��2�(�#"O��x���3oLl�:��ԓI~QB�"O�q0W	�L�����ՏbC<"O��i�HX7�^{@kQ>���C�"O���,�`����ͮK��$1u"O��HS�LN�J�2�$�7�=�C"ON�8Q�7.ҝ f��0	E���"OҨD߄AX:0p���IS��p!"O�ā;&�ZW
3'��}q�"O ��V���x���
./���e"O�ɻ� %��!4nJ.B��0�"O�y���L-���L�9["�H��"OJ|�u�߱}��N�n��X"O�H�2�F��(D��ᜰM��0"O�h�ⓡ��d��*,�8`�"OFI�`��-Y�~�s'OK�ƑX"OT3�1�Ru�e��IE0,��"Oz��O\[��5s#���"|1w"O*�%@�*���ä��$h"İ��"O����86�����*:*���"OVAq��L�:���30M�-cU$��"On�D�^1p�
��lE�I�`�0"O@T�����$��e�ɾ{5��f"O�z1��>:�&e�t�� 5 E9�"Oljm^�!���t�Ґ?�!�U"O"5�Z��Y�pe��r2|E��"O��:a͜4�t���[3��H�"O@I���05UΈ.4�؛q�&{�!�D��+cP,�J�e��#�Õ$�!�ď9����#�u���1G+œ�!�� �93��co��⧇��s��1��"O��hX�3���h���"O�څ�O"y�$��C���I(�:f"O�D S�"R�Ճ�`
�Pݨ\d"O&3�gD,l�"ݐנS���Cd"O�=*1%���U��4;���'"O0pya��4cxH����C�z%� "O���I�w��Ȩ0^�V��94"Or�R��%4j���6+O4;�t��"O&P�NY�x�P�J�,�\D�Q"O�@�G�I�Q>D���F�ckn�Z`"O�m��LP�u�j���S4)W��3�"O�&�DQ��a�2�`+^� ��'M����e��svX�d�@��'2R�0��D2^���3�kPZ�C�'���P��1_44��J�=^�I�'T8UcY�vi I�4B@�I�����'��̒�ս �6���in�H��'pB �q�̤_@>H��V�j��qX�'�b�⎔  z%ǭ\���y
�'E��Ԇ�(����A���H�'c����H��v	~ !r�Ǚ1^@�p	�'�����/2����OV�'V�#�'��--i\��jİ�|IB�'&�r��o��F9s����'������ȎcKl��ÆerV]��'$�DKpρ=X�F����%c�n�{�'�R=�v�_Dh�hH@��7_�(��'�x��`�oD���Ao�B��'� �(��Z�Q�f��q�Ǒp����'A*q���s�
�AE�kI���'�kؘi�&� H�2x����'j�Q���H�Q���"&��B�'���vi�9[���#t�=j�'����4��:q�ajB������'
F�Ũ�9�jH�a-��ayЕ�ʓi-C�ғw��p�",�H��ȓM����!M�b�B�8V��%D��X��N~�h1�� وY�wO)}sp������#o�3�LPdM�q�6Іȓ;�2�ӄ�܊��,�q�WH���>E�i�"ϋJ�Τ� (��_q.�ȓ6?H))��Z�t@�J��[0���B��"�/n3�P�Ä;C�0��+D�Ȱ�7�1:J|��k�5�y��Ji�)��P�g��0sg��y�D٘|Ҍ����T�d�i�B,�y��ŀX�ج:�J��W��� !E�<�y⦟&I&D��ȢNѺ�±�D-�y�h�Tq��"�W'@#�y���yR�SO<�|�f�<p���ȱ�y"+ˠ>�8���a	9��-��yB@"�ڌ����Cj02���yr+�j=�9Ѕ�<�NP��O˖�yB�܋q�⴫S,ӕ	V̪�"��0=	��8gpۣ-�)0/�y��>0�X ���`��Hfi�*�yRO��f~�:c�S�W��b��y§�" ��|�-�w���#!�S�ynW
,a1�BP�8-މ�J��y���)�����]6��=�%�A��ybe��d�0 ����)q⍑�%��y�,�	&芝#7e�0�Τ���@��y�c�c���K��\����a�k���y
� 
�QB��r��E1db�"s�lkv"O��{��P
ucd���A.SL��"OZi�$��+�d1��!L��QQ"OƑzV�j�>�"w�Ȝ��]�U"O@�X6 �U���ic��3Uxtxg"OJ�A5
߈>uzU� iR�t.\*�"Ox%p���2(��� ��$aص8&"Oz��%kؾfX��YB�� Wn�%A�"Of��Bc��0�ڭ�B $Yg���"O�P�@��΀J�o�FB�:�"O��q!�̱g�6�Sr�G*w��QC@"O��!@/l����T.ʢt����"O�{떄v��9+��פ_	�A6"O� ����b�N��gP#g���"O:y�"�YF�F�C��8s���"OFeA�$��̴ ��ݹ]�بq�44��)��-<8�PǨ�Y� ��@6D�D#A��"xi&�)y�� ��:D�@k�[#U�Z(b�!úK�R����9D�T3b�L5��8�!&c�(�f�8D�ģp	�;�����D�C��7D��KAD�|2���A@�*;���J%F!D� ��a�=�m�T`�<G�	�
,D�x[�T�,|��`��\�a�qp�.D�d� �@�S�X���,�;)��B�/D�dz���,��9C�Ò�
�ؤ�(D�t� �;U�%$.,/d]�4�'D�dpP��53���G���p`�#8��p<!Ec�7xt��xs�Q�&ڱHaf�s�<�jH>^qғ�����S�r�<�cK�Q��
�8?���)�ɋq�<���J��x��߽7�(���X�<	��
7����(�:Zo� �a�U�<�'NN�$�*Do�:[@��T��P�<)0G2*y0,J��8v�\|�DOS�<!0H�~ D	�gm�,SB0���d����'��X����sdHq�É� �朙�'�T#��I<e�8�B�N%d����?��T�&���+�'A��G��r���ȓD� �r#J�&�@*�Ƈ?�a��}?:�D+�]B�P�僜8���'d���F2�d ���!E��`�O����L�f�D��,���4:�煛n�!�DY�gr@ZP�K3P-h�"�d]��!�D��Vbx}�'�b�*���;�!�ϵSQ�A��]�U�b\�U��8
�!�$�:9� -8@4W/� ��ȓl3X�L^�u%H����F��@�����E  4b�@�a	�J�X ��k2 ��
O�
�؄bs�
,JX0��b��,P�k�?&lt
1����ȓ3�2 PvdR;X�n]JƵS�Xфȓ%|���$��G��!'!G4<$Ʉȓ*bd=��k��f�i(�:1X���ݔ0{"��+���y�cW���-�ȓlP:��3J�\���BvYx,��E�l1��gwꜪ`@_r�h���-���q"��9K��FDQ�cF����?�@E�*�	��S��� �PY��g��1"Ӭ��������|�B���5`���`.ܤ
9�Xi���PZą��S\b�s��Ȧ2�R��e�,���`ĸ	�����e�&/�$��ȓ-e>��-N@�d�3��Z�\���S�? �͒W�Q�5".J�xT���V"O�Q*g��v�"��L�",�yB��'���2�H�(1"�?Y���JD��&QT!���5qF��bL��7��t.y=����'6A�pHX�C�NtT�!kL�PX�'�5b�Aѡ?,Л#��j�1(OZ�=E�4�2����c)&4�2 C����y��0k��0/��*����uaŕ�y"�Ȉ:L#1쁶W	�-K%Ȋ��y�F�U�&��m��'^��S`��y�c_1r��Ј7�.߈�"�h��HOƢ=�O�6$Y�kߔ����*86���'�Zy��/4)tU��y�������#�6�tB�GpR��f��:2����	W�3�Tȅ���$�T�k3j@=�>lEz��~�Ŏ��H����tX\�g�XW�'#�'��'?\
�Q4a�|y�32`��TI����'S��Ȱ���l|a^�� �"
�'l��p��ӒW�l@����njy�'�<4�P��Rd<ðC�8_��!��'�4�
��
�SOVTk�?O��i��'ŞU`҆��T���~d�x�'�D��3���
g�ڡx~xP��'6t%�P뚄�t}�!'q�x{�'"�=07�E�0��0�M�42����'H�|���W�*��5,��x�n1;�'ߪ|�S"�?#l��lʘi�E�'�Du��]�.��fF���"}�
�'%���4�Ϸw��(Q��EUz�
�'�̰��a��E��eӐ�E�>�>���'�D�`�j��LhD��kOm��l��'Q>�� :j�$��-�j[�� 
�'�N<�3��
�����F22D,��	�'Ѷ�G�F�c��i�Ȗ*{r�I	�'������N(L�{f�O�A���'jRxP��DC�:��RaֳJ��'� �*2c�s�\)7|���P�'�v�2�&��� �j�
t��u��'��d;A�J+�r�	' �^�ts�'[`	#0#R�jѲ��0�8(2j@�
�'��� Ŏ>��!їIU����'�rh�$lO�@�,,�\��4P�'/�ĉ5�V4.��A�Tc���a2�'��`�`#P�VDE���q�h
�'�Tq�a(s�Z��Ϊ�\��	�'ԦqK��=*k��C�h�}�T�Q	�'�PE��lE+j���fO6��'���gĎd�&!y3� c����'v�l�������sr��)\���1D����ӭ>��sU.-M=yAb,D�<;��|�6�yv"�.{J�AbU�<D����^�#�|0��Jf��ڶ�<D�<�P�_"=:>�	��Ah����H:D���Ua�l����D�ߟ]��@���"D���=/��3r���rx�)�n<D�TtO}�D�"*>"�	�Gd;D�`�e��(�H%����aJQ:1j:D��0��]�z�T�w�����4�,D�,k0���It���2����A.D��S�hI�*$�)� _�
��SP�!�]���4�A����<	���.{!�C
P���;g��v�J�ʷ�W*. !�d�uEFH�����+KT�#u�!�D��CH�q���Z豰S���J�!�� (�*U�����/7�($�V"ONZL@~�"P$���n�b�"O<�@�'�5��D��C^�v����F"O����k޿ G� 2ТN3�j��"Or͊��Ԙ����QD/M��Xq"OЙqg���� ۅ�]�V��rF"Ob��q&��*��A��'MP�6"O@�$ޚ1�Erv\�ZAN59R"O����-_X&y
�
�[@��"�"Ol!Ȧj�<sBi�� ЏK݂�"�"O�c�Y/h���w�%(�f��!"O�钔�ƭxj�X��	�R]vH("O�`T�R�0��Ʌ�?���+"O���ٹY[d�k�ȍ'��mh�"O�y�U� ���&�y��b�"O�4� ԗ!)�]�垽C�^iʀ"O �	�F��=��˞|���{"O>t�un�?@��� �!����"O�� �][�<�x���)��h��"OB`�Uˊ�H�f�sW��l�j�"O�ٓ�i{�h��UQX�%"O֔Ӓ&%&��sB$ˣ]��85"O��`��<0 �!4i��x��"O����
��+GNE0�j��|kT%R"O��+��[�Q�0��H@M8�q"O�pP��Aʔ��V�' �aw"Oܐ��T�n ��ҝ)��\��"O@���M��Z9�@�m�&��"O:�X�D;d8J'!����"O���BA�S
~���#B�)_T�w"Oxu!��$(p\����I�'I>!"OL�BBn��BK��� �Q�QX��Iv"O��Q�$�%-,X��n3���"Oj�8%��Y��P;g%5X�2���"O�œ�������jG�b�0"O~��ԣ݁|5"!�Cj 9�x�Ce"O�D�	��o�t�IIfE �"O(mQ ��] p�N�p�:�"O�$H?-� �`GT�z�H)Rq"Oj�	�Owi��ۓ��<.��8#"O)�C���]�� ��b�U"O���#�7'FZě"�A5~��q�"O��8��#��)�Usr��"Or��tH�&9%�����l� p"ODM�w�F�2�yf�ږ3�0�x�"OƘKE�A4J����`h�99���"O�(�#I�'���A�����Sp"O�]+a�#�����J{��"Ov��ïF
A�n����Zv�"O>Y8ĊJ=��*lWq7D�a"O����ƥEj�EŅ�.�ʘ��'��i˛x�� ��!��a��ȓ���3��YZU@F�B/ܭ�ȓk+e�'�Ø}��"fK�?�<���=�1��cG:e���PاI�M�ȓ49���B�y.ipg��:����� ~.���ɻ~�X��H�T�����y�HŀVI�Mt����a; e�ȓO�",j�o��8��ܳ!FԞ$���ȓ[�N�C3�S�:�: �R��2'<̅�XRjl�UE�	�Va�6L�. 4�@�ȓf\�E��.�7�|��h�L
��ȓd�byB2� N�La�G��w>$��#�ꐒ�ęt����6��
�����S�? A3��%��pC�g��v'hĲ�"O44O�CI,��#d�')B��V"OЍ+�*3�;�b�	#p�b�"O\##�I9?̱�q�ܧh8�I2"Ofx��/�-!δcgB�g�^��u"O�5Iu��b���J�!*f��<Y!"O�9sF�b
����m�B�v"O�xH�E� a,�2d��Wz��С"O�q�DSQ�\r5b�26f
A�"O��%�O�EX� �co[�aX�"O��� J�/-ʖ�H�B�7M� U"OZ`���κN�,�'�`���"OR��6��I��y��n�.X"��"O��"C��j����׮N�PϠ1�"O8A��J&_Oq�"$ւ|�h�"O�	4�W:`.�4�'�W�X�h�h�"O��R�I?`h@��@�`xK�"OLD�s,�Vt�#썴f�v��F"O��!�C³G�Z�d��I�((#u"ODE�U,�#$u��3C�>0͔Xs "O(�I��V0�H�F�Ł ��)�u"OԘ�@��<,Y���/��\�q"O�4����[�x�����Uw�	i�"O<�0�)l�)�q��C_�t�6"Ot�:qd
n (+��1�b��"OVq�Ԋ�@}nY��0�lS!"OzȈ��ն_X�u.U�.Ǧ�U"O�YPԅ�y�%	�l�c�콂"O�5�� ƌ����ɚ1N��Dx�"O�k��J�n@	pFY�lxvڂ"ODD 0�вQ����AE�Yn�@w"O:�eI��8X��Aϕ>�����"O޵"���"6����cf�3<(1i�"OBP�%�U�m��8�f������"Ob���07� 1P��4g���B"O��b��9.ƾa��݅' �HG"O�u���>"��B ��58��R"O.��-	��v�i�mE(ln�B0"OJ���	�72����f�צn� �9u"O
u����^���8&"�/���+"O�3��>*>=(EF�<j(�kw"O�d��JH(��;dD7<�x@U"O�c�dQ�)�Q���F2��v"O�!�I���!�E@$.�k "O6�pWO���I�D�d>Lr�"O ���,$�\�s�-�4"OlkD�M�b)Y�ʒ*Ԗi "Oڡ�g1QHn̆Zt�$ �h&D�(ᗬ�=6x��Yň��m@� �$D��cNo�a��h�,vu� ��D"D��� ؠ1�|eK�!�+\$'`?D��ѳ(&�![�mE�<����#�<D��*S��KPpuj �B?K\����9D��
5H�.8n��a���m���`�b$D�(��)̮���� ĪN�հ�.$D��!���M��<(�@��x?9���-D�А�.(�>��"@\<�\B�',D�ع��u-��QA�Z<0��$s!�)D��(`挑k�Jtz�o�fFA	�"'D����ܠB(��@*L JL9��%D���ސs��+q+ɍg6
��@,$D��!�Sm����ȝ0{ ��B�#��?��i�!.m"	c*�!��M��@�-8!�dĖoI�bv��@�$5BP�۾V#!�� �
�HC� M��g��JYd�b"OR���/�X�z� ���>�ɨw"O$�{��J�u�<tɕ��
2���"OБ��M��+R��1`g�w_�M��"O�����=�@��Ĩ��tW�P�6"O�<����K��RC�[�R�(`�'Kў��֫���HsSDκ6fD\(s0D���a�Cv���F8B����"D��0�鄑CY(��rKP�Jf*� � D�D�bM=�T�	�M�"��!L=D��(a�:N�,�p��̜*�b,p��;D������5G8�J
�$�x�q�l.D��b���	����D�Z�3= �5N+O��=��+E��D�1�(�yWFQ�C�h~��|��i>Q1`�~��E�J�7S�����>D�R0L��B�@xk�n�,�x��+<D���$�N���#7�2j@*�hւ&D������%Ϻ��H�n���6`&D��!��A�����I�V��Ӂ&*D����-Ih%e����5�Bg"⓻?q��)\�%��[!apT��ӢpV��xyҚ|�	�1=sF��@c�P8����X�s!�$M%E<�2$%ח(3��+��6!��f�Bm���"n(j����@�7�!�$)��Xia�L��!��{!�d��rn#Q��0Wr����'8a!�Fw<^�`�<)�\dATk�az��dO�h�����^G*�H�4G9�1O�=�|��f���ȡ��G��h��ju�<Y���WC�E�@�	�$�	
i�<�Q�נ_�De��i�9�l� �I�<���ь9���RF�R��L� jL�<y���?m%��3V�"WGȵ���I>R�z-��7D�,{tO�|�ZT97싔_�x�� �:D�< �!Ϫ;B���!K�'8I�d�9D�dc�+B��^ijGKH�lx)�O%D�4E��>q!�X�!��=��h/D�Z ��>�fi	��>NsB|�M+D�@�"��g��E*pO*�Sd'D���cN�j�	�񈏗m�lp@�%D�Xr����T��Ɍ��1�6D���
�7�����e��U"��9���	��I!��)VTv� ���
�zC�	�*tZ���M�r�p��'+֊DLC�I�x.*���^�,�p  �%R�C�	 
",��6�A'��A���"!�#>���J&����B�2�������z!�R��4q
"�+q�A a~�R�����E�A�\*��\�����*���I����+� p�&i�@�ĆƓ.�rU��I"�j@�ii�(��/���F�O��D����`�*���B�S�G��A�nx9�{RX]��-#İ�T�E�D�Ё���^�vP�ȓ^8,�E=8�M��6!W蝅�	B�,������)��F�S#1�B䉥�<(RLѺt1��&�nu�ƓoF95�&Tt��Ԡ��-5�!�ȓH(A��ɞ$3�@�X<!v���ȓe�(si��:�/Z�)�c-D�Da��@#Z<N�#ORu"jԂ�-D���hN�K3B�?a��ԓw�6LO\��2��]��e�4��5P��2v��L�!�d:5���C�P�B�|R���!�� ������ =ob�	�F�M�J�JV"Or�
��M4�,��놤ӎ\�3"OR����6��i�*P ��=ȗ"O���&�(��y*c��9��ܐ�"O�\���P��D(� Q, ~D��"O
I�U��"�b��֣֝��"O�i�F!��^���� �b�;��	Wx�����6#$�dQ���Z��o)D�ȲQ![6�,����1_�����&D�T���//h� �.�,a_t�f�%�O��6{�(;��G-[����%�n���OyR�(+v4!`�	vC��yͯ H���� �
1{�,V4�yH�]��Ӗ�ʹt�m�q!��yro�0b^x��"��gd\)!�O��yr�� ��n�KA����5�y�[�]BT�1�[�EbF��S�M��0>1*Oh�d�#y�"���-�Z��eDAn!���O���5�˺���7Z=:�94��)�eU!o&L�q�A��|Q"�?D�܀0������C%N|���4"=D�,���J1^9�4M;Y�| �Ph;D����m�1k�8t�Љ	�#�J����;D�8C��ˀ$ d����� v�2���i'D��!
�V+#���[��$D�0k�`ֶ{SN��� ֈU��а�5�hO��.]2�E�-�*\n�Q#�&C�I'+&, ��I��A�F�y0 H8T��B�I[�b�2��(;�,0�Q@ʝOH�B�	��"!�2���-�Dl��@�B�c|����I�/�&d���ܾm��B�ə����T*�'c�@�&&:��C䉊e9æ3M��(�%�E�C�C�I�m��09�'�B���W2��d�9?Q��ᓷ4��|��#�`0�#f��0۬B��2:�xVɈu92���~[�U��'��f
�?RܘA+��y� {�'1B�U-ĩR�v ��Q�j 1*�' 2]hv�V'E���1aK��gT�����'E`d�G �.�pT� f��1�i1�yR�)�S��.!Q!b#:D�@�K�]PB�-6fmi�"ʮT1Ny`%"��Q�B�I�T� ���Q�#|	񢉉4)� B�		da@Qkc��b�<q�.T�"NB䉽3"Ua�쀄C3�Xb&��+Y�*C�	�WzP��O���|0GdA�Y"����2ړ& &��*�ZY�� �*���ȓ
�����oͷwl�['A�`G���ȓ?���Q$*ʬ@������Оjpf��Gm��2tD�kR,\���55/���kڜ�¬\�y�R�f4�ćȓ&w����B -*.�	��zʆ�ȓx�����m�M��$"#a] 4�Vфȓ!|F��`�6_��в�P�`�̄�'ԉ��l���P�� �˞B�b`�ȓ0�x�@1ΓC����M�l ��'�ў"| �W�k�P� ���&q���B+K`�<i�dU�=Yp�_�Y�d�V��\�<1V��q�$���v
�%bGL�D�<Q�*�8����P&�D*u��mMZ�<A7E��1O  ��4rm�x p��|�<��@õP�1$ Z�?��x��v�<�OB6���@a�(ӌ�;ɉ;��d%��s���,�^`�<S1�Ѥjy�5��*<D�� ��
���&5|
����*	d@A"O�ٰ�%ܫ�bhRCHUv���"O8(і%��w�L�$B@<��-��l"4�H ��4c�B�Eƶ�K��6D���aK�*)��8��ݓ�x�a'*D��AG�R��GA��"(�H�S@'D�d2p+v���聃U�"v��D#D��"�Eł��	���0�^�m.D���A������!"[! �*�n�F{��9O�|��ӠL�2�: f�t|]`"O y�D��S��y ��_�P\��"O��ed�#��|x��L4FX6�b"O,%3 �H��t5���6D]h"O� �!@$#�l4�0�ݶ0��"O�ѓjHa`t8V���O��Ƞ"O
����M�Y�Qaf�2C���;f$8��|����'�.��P�[�	TJ�S'�6�@q �'{R��%�X��xE�Q��>vt��'=�����RH�B`��ނ/c&-�Ó�hO��j�C7t<�8�A��mX���6"O�iW  C�pm�RW��)k�"O��B�E�$���Eǁ��Z"O��Ц�2�X����W�T�VDk�D?�IV��2��͙�e&~�����0RS�9��/��A��͒�jVMR�S+D�����s��亣h,�!�h'��hO�S�>���� GH�U�H13I��#�nB�*Zh`�D�lvR��A�� ��B�I�8�p���M��s�Y�`S�zu�B�	�T�� ��]�	u�2��Ь#�,C�I#GRU�/�?2���6+����ȓY[$���'˫d�p@3ũJ/R�L��ȓP�n�BW��"4<F�:��K�`�E|b�� 956T�u�Б$�T5����Y7�C�	�	\��+WIж{W<��5$#�vC�ii�dF� R)����
�$� �
7D�HC��P�9b`𣓘+�hq�K(D���'�(B�Д�Q�}RX���(D��Y0�ݺf�H&�\�%�l���2D�@���#�UZ��X�*����e/D�&�2�T��%�� Ҫ���#*D��P�'\>�����Ѣd�����k,D��P����,�TaQ�-�r�e�.D�� C�O�.c|��B O$}Q�C� +D� !�+�2< �=�֩N"2Q�N)D�|����h�:QR��92��*D��y�P�q&`�C����)��L2��'D�,�b�G=�5Y��T�4Ϧ�xc�:D��"I_�V��գ@��c��q�%D��c Bg��]r%L&,P���cl"D�L�q�y=f�tK�,!��-S@"D�P�Fm��'~@X�dIVВP��$K!�լ|hh��1������mQk�!�DM&h�@��Ka���p�&�2~!�$�W�*����|{��:�LK^!�d�� X'@�{b��7%uj!�D	�)S���cG�U�Gc�Yf!�$Ơt��p�ԃ1K�I��/�!�/aP���g��`?�� "� c�!���igv���nS�S'Q�"h�!��3l#6�I5�4%�e+��!�DO�&��uc�K�nxƌ۾(!�DU�i�~��ˆLA
����&,!������ ؊MH��."!�� �<�G��8���	0cR<GP�1"O����@ŭ(_NQׁ�<�,�� "O��x�'��.[�X�
��h�Le*$"O�̺��@_�2e��o��-�Y��'��I:,$�8�e�(.�=P0I̟�*C�I4 ���SO��8KZ�wˎ ��B�	 o(x��'8�,y���6�B�	�0w
H�%�̿0����+��,oHC���ղ����[��� �R�C�ɋ-kl�v�؏&i���3�d"C��.b�:8xB���p�t(2:���)�����,E���#'��D�N�w!�$E(���Eح?��3qD�jv!�\0���h_�����bN��^!�d�ybX�@�\�
�3�Jw�!�D�u��rG I�@�N�&�.�!�D�O�~�u�V�x���i'e�
?�!�d��=��i��"n�zfK�2�A��IKy�̝�J�8�0f F/Q���Ǔ�y�϶c���rAjU�K/dq����y�*���͓F��%<&�;��;�y�߃_@0�8��ƺe�9 �g� �y��S ����*�(j�*08!铄�yb#Z�tv����G�6d浈����y��A�n���s�,�)	�ͱe�����:�S�O�PI�䍃��ء�T"Ҭ���'�6Ezt%�X�VxC�zv��'j�H���/2P�6�S)�����'�(��.!e/�1k�`Б#�����'O�����
&��eγ����')��2C�,c�D]�uߘ�Vp3
�'�بŵ�g ,1�5B@?m�F$��'&��Ċl>� o�..צmx�'�"� ����8<8��$ϟ#�P��'}�mv��L\��aW�1ެ���'������/N���6!M�|.�%��'�АzD²o'xxꕁB	u$ԩ8�'��ᎂI�}9 ���<m��'�Z�&I�"D�d+E9�m��'3�i�`o��t��b�'��sX�{�'�l��==��-S2���[PH�	�'P*�!�" ��D���@H�'J��;�*�=(����2{�J���'G�A���I�ṴCfQ�4	�'Kl�ن�މ���"��]Bh��'b[y�ډrZ�� d	�}�!��'��Li��	�2��+�N�A~���'}��cΜ�f�lq{��:��IC�'����sdի7��;��J6�N]��'�HA� H"v�<ત)�z��4��'�`p��CP5ed��1TÐmϬ�S
�'��ĸ4��,��Z!�r�d5��'al����t���[��'X�x���'t�����D�)�\Z�h#%!����']d(���Ts�Ң&M� ^�5
	�'5"���nø<_���Qb
L؂j�'Bt�� ���|B ����ǰ�b̺�'�B�(�cUp�4�kj�z�'~�ze�Ϋ�H��c�\$�'n4��oR�V^b �l�<���'��M��E�h`z�qt�*�dQ0�'֠8��D#k����̢'8����'<*$i6l�oN,`����J���J�'��hj���;����ǩ�6������� ��p��D�sT	���4��`�"Ot$��g�pP�i���j��$z�"OR1`&	?Ge�͡��)eN�H�w"OЍ�!)��-�qr���~�*u@S1Of����j��X�RW�R���V�g%!�C"D�XA��-��_����$
��B�	��.��u	�*�r���R5BW�B�
I�a��%iR:�x�`��zB�6Uj���Nۮ/�کѦژ�fB�Il�(����/(��]�tHV�1JLB�7{�,E���Hǆ͡���M����6��� C
�0@�$ܑ��ki!�dE�6�C�aץ i���O2B�!�ċ�1!
Y)���<L��wm̧@�!��!-���;bC��A^�x�w�C�B!�DϺZ-�vKR%Y�Ͳ�у`A!�Dݦ��b�nP(*<�<1Ɏ�e9!�D��A��d�@��o7�e���W9!�d�,}*L�P�؛[-��#�P�!���}�`Z5��6G��I{F�[&+�!��%����!����4@�V�ӟcu!�䁒Q��KBAE�L�d�:Vg!���؉y��Ç5�Ftq@�/S�!�D�4d�̸�'Ȝ@�@q[��׬y�!��X����ÍX��~=�Ҁ��x!���t�c�`����4�H�!	�!���ڌ�D�� 4� $��(5h!���_����4��nB�A�#,V!���g|؋�נQ�&�ꧦ�&Fu!�Ď�hW �΄$���;�[�6!��
0 �*�`��:沰�'#�I!�R�s��\*3�����B@6!�d)W���BY�x ��`�@N3 %!��l��5q#��C�B�(6/٣z!��|�H�T�b��ճv-��h!�D]���@���Lb̕�!W?X^!򤅴�T��ݎ�M1�k�g|!�dҰ;�(A��$}Bt�8K!�F��s��ɢ{M���JT�[�!�D@�e�.i��A]	�2�� �&C�!�d�,��p�D@,v�MzB�^�N�!�7�D�KV�F,e�"Ӧ-�!�D�%q��qQr����l�D%��%!�dK�z���S��	�J	{�#\P"!��F� F�����k�\�� ��c�!�DŻ$�;�������g*�=Y�!�d�=�~PS����pL;�ɛ�p�!�$ݗWUR�&E<;��W��&E�!�䒟U7�șuA`��d�8\���`"O
�V�ұl7�1R�fD�y��6"O&%J�J����p@�.Zl�V"O�H�A����v!̧CN<{D"O��)�&
�>�9����[I�mj7"O���kSv|m7�]�{xq"O�ذ�.̤S��+�څ
�Z��6"OZ\Z�!Ēd�x��`���H�"OVK3v���q1�	Og� u"O(W�-[?M���ƥ���a�Y�<�#�ݽo��JDD� k,�q���U�<�a��u�zP�ˋ�Ϭ�9v�S�<�Ea�e�&�P�P��y�%�[�<Ձʎ7ib�x�*K����mLa�<IƆc:��BfO�1]_��� �]�<Y���,<�C�#ժs���AG�U�<� ��)���\���s7$A�.Ѡ��R"O�8�����:�%B#^ƴ}�"O�(� m��AjI�ք�z�V�aq"OJ0I��.3B�*V(Lj ��f"Oh=H��N(o0�i�ɘk��C"OjS���/
�b�ae�9����"O��c��F�`��7tP���"O0��t
W3����,����"O:�)Y�&4���0Fz�� r��]�<�s�M�I  �����7g��$K�d�<)CoA�]��Ȼ�Ȝ�`B����' G�<��%��<�B��ʵ5 ��f&�F�<I�-pRB2m�e�n�	�IF�<��M�6�@9��>�2�]~�<iR�E�t$Z��㬓/eQ��a�EE�<��/4J���2B�ҩ)����7�P@�<�FF٘K�d�geZ�v�4I��_�<�O>�-O1��IQ6��,�.�Y��)
��1["OP���F��fy�U��cm�h��"O ��EΙLg�['茷?UF��"Oļ�X�!xg�C�Ĥ3�"Oʘ¤P�nx:�P�A*Kߞ`a"O@u�%D?[r@�R�%�\�
X`�"OJx�d��+n�ۣŇ�O�(�S�"OnE �,��W�d���P%��M��"O԰��%�O�8G- �B�T�ٷ"Odez��Z"y�A��жQD���u"O����-�4|��{�(M�����R"O������G��%1HL�ۚ(H"O�;�-֣rKƄ���8�>���"Ob��fG�0=��	�n��` �"O�&��/�i����'\\Q3"O��p(�*UV����Cޝ
�"O $�ٳj�����_����"O
�2��� =,���\�"���X"O$	�T�ԡ��R�x�P5"O��$�/&[*P HE�Z��Y�"O�(p�Y�݊���)�XB"O聓LY�m>��pi��p��5"O����C7��U&y������]�Ph	&$�����.�U���ȓp̾('/�\�d�ڢ������pVGM����Pa�P'�ȓ;��%�/��0����T��;����/u�)a4�"x|c�o@T_�̄�ch0 SOJ����"U�>��d��8�N�	��.n�b���jٔX��ȓ*;�4��ʂ1�V�@�L����,�����;��#2M"/�ȓ)��Zt��&JQ�!�Dx<��B�'SԐ�hG.Ͱ��`��*9��a�'ֈ�`�pkV`Am!&��k�'0��TfCC��x�PǓ��R�'�t�t�!BĐY�㓝C���'a���AK�;3�t	iԍZ�>���''pS1HHS���:�O�m�bȳ�'J�p���-��9��jA%kR �8�O\�=E�	!Y����=^1"&"����'`ўb>����ň H��b%����,`u�0D�{�o4W��r�K�*�h�T�/D����银f	x�H�ǉ^���5C-D��Ae�5]/�"䇣(SrB��)D��)��/[i�`A�@-�Xa��,(D�d��� z*Lp�b �ͩ��1��hO�3� >1�c'L����r��%B���:6�1|Or��토{�.P��,�D�:�@"O��AwL6P�<�	����g�>��"Oh�&�sޮ�+Ê�'P��`�e"O�	b��d�r��#�X�3sLIj�"O����n�RXw�M�s�cA"O�����^�K-��Zq�LlB69 㗟�E{���0�t�!��>y:u��H�V⟤�)�g~b�L�I��ei��E*�l�Z�E�7�y2�]�ST|�1.ֹ%�^,�'�ѯ�y	�$$��-ZQș%>��)w��y�ЇY�Z�c���v �C�I��y��Z�<� ��B!D4���3b���y�c��J؅�'�Ѯ����,Q��y�+�P��M�-&=�5�P�؟&�ў"~� ������vUde��@�g�=�ȓo���"�H�]ĆuKE��2:q 0��j-��l��@��Mb��B` �X��'�|����9$R��0h�M41��'�~DR������S�*�J.T%Q�'*�QC�cB4��A�R��4E��H
�'��-k���;�Q+K ����O��?�,O�d��	�!�5�;V��i�נѽw�!�B,"��2*Br��p��A�!�ē�/����bJsАQRb��Iu!���B�Ltb�ۯ5aȵS� ��a�!��"����Q��T�
�9EmVN�!��J���آH�,{�dhD��g��<D�tf�q��P�WB�`�Ȍ�`*Y&���,�O��G�(�q{F���J�d��"O�t�����6���ھp�D�'"O|UKuë*�(ễ	�'	:H��g"O�t�����^lz��^6^CViS"O
���-*QrECC������p"O<�1���e�I�B`ڪKUh���'�ўD��!Y����L^p�*��M'D��hc�L#2P�#�(]3Z�ƌJ!J'��h����Cݜ&x�����n��3tc D�0Pg
ш��m��
ـx��eJU�0D��#�i[�X�(f�w	��b�.D�̡'DI�@M0'��Jb�;e !D�������5���>�8U���2D�,S�e�>�B��`����'r��G{���V�2.8aV�W	N\�	��!�d+c�9p̩[0�5!��D�$g!�ؔd���R�J�{�p  ��',�!��7b�ȸz�"����ŀ!�IP!�X:G�p�f�R	t��9`1ő:.�!�H�XY��5�M�t~P��eT��!�ȓ;�ƈqU�+)��#�M5}axB�'��O0T�ģG"�1+3��<}R��r"OV k��ɼ���1�?tB)�"O��B$�G5E��q�@A�&;cV�@'"O��ۅg����6��/qF���C"O�;A�/4��q�2NUf�i� "O�$��n�b��t��L��gL�ȓ"O�L���'�$�ya.h�4��<i��I�%cҶ8�R�W�p�:,�EI�
<!��.N�D)����'D�N�x6��J$!�]$�䱀D
�'�lꑉ�4W�!��c�}�W�_!s��#�Ǒ�B!�D�?v���Ȓ$g��5����-a|�|�a]�(�Pd�j%�x�.�5�y��J�?�  ��/�9�&L���� �$3�g�? ��#e��$K�ε��`�eG@d�e"O��jQ�02�����"�7)Rd1"O���LS�6�p7!�_HjQ"OD���J /WP�F
1�X��"O �� $��FXUH�;TP�_�<��E [� �\�J"	U���B�@���ba]� ���%g�]|xE{��9O�%���ܧ��-�!d�V2�"O�[�̝#a�|�Gj-#�"O�5�&F�� ���q��9$�rU"O�q�b���l^�Б��0��4�"O�(� ��UfRUI����{�"OY�h��I�F�\�Ȭ�vF�O���� ������Γ �(�A�nf!��y	�5��_|ri�VG�o4!���S` ���D2hb:t��+{'!�D ��,ZӊG2rҭ��F�- (!򤟘B*Ё�F	!i��!�ֶ7!�^"o�2t1��6S�k� ��!�dG�{>��F7><pY���P�1O����<q.O�O(|�F���Pz�9Cc�Y%~J"9�䘟��ɧ%�zH�Sj	g��ZE�?��B�I�,*i���Ťp�Y D+	��B�\����[��Su�Dg�B�(�@I�Cϵz��􃦠.#J�C䉍e�gF�\�����!"�C�	�j<��������/Ȇ����&���^��P�#�	*��1���9a�C�pG�𩲠u��(s�U�qu�B�	*�T;A��x2���"��N�B�I�qH�d�E�K/�ҡ�Q�ðR0�B�	�N���ՠ��|)�W�D�B䉉1�@����M�o�N��O�jYfC�	�E0�D-�m�-"V�D�T�B�	"a��[g��7'��;�"�l��C�I�:�.TC6 �m��}h��uc�C�I�`��rT�A8t��)BV�U�F��C�:^���g	}���!�B�	�rj�$��-�/dʺ�Y�/Ч(� B�	4i�h�j�
�1`�1;��Cy��C��#RQ����TȘ�9%��)^N�C�	*)����N	il��a�uP"B䉑bƢ�E�͝spː ӓ)�B�	�8=A�b�5c�� S�+��C�ɣ\�>U+�C�-uL���%��)�C�	�`1�l�6U�*F u�'fۉd�B�I9a���;�ۮP��ܩ�NX�T)�B�I?|�5ZSAƈN=�h���_��B��04^H�A	�
Pb���mAs�B�I/�&���G8N0D�{�c��t]6B䉖~������#D^�����s�C�?RQLy���6Y����l�4*2C�I�T�0�q�b�#Y��]�`�^a�>B��8C @"��R�P�t�Z@5�B�0aO\ zK�&?�f��ĉ�=LB�I �,d*P
�1�Z���A�qNC�ɘG�<}�����ؒ�@�?h�VC�I�{"ؐ�:@۔d��C䉧O/�d�7n�_Q:�Pp晧)a�B�	�J��(��&.,8sm�p)rB�ɷZ��b�΀�2�`y��S+<3PB�6g*Ix�j�,�삶�=,�vL�?���|ʌ��'�n�)�M���Ha�j���'��u@3�ۗ[@h� J&>�M�	��� �MK�)�&���a�c̣K4]ѡ"O���S	�3�@DZ��L�g�;�"O�t!�J�;,�0�J��[o�l�K"O���� ��N�D�� D�I�&,{C"O��5��*�L(�#�ͬE��͉S�'��|BĐs�:�)֡c"Hj��_�y"�ۂ.���T'��R���o���y��äY�X�#��
��@�#�>�y��	���6"����� DE��yR�؏>�q�CN�*w�$�K@,P�y" ѹ�D�)��E�B�B���yRaU�d�<�rl�.|
���"^��y�Я87���Ü  Vn��qbܦ�y�B"JAS�D�+�$!0�y��cX 1�l/v�2]��$N��yRF.-�ق��V�u�� �o��y�a��wԼu �� !"�-�D^�y"씳P���iU"�� �!.[�y�&X�.=AA�'lR��q1�y���p�p�{��<�&�1Pb��yb��56	�b��0� p0p�B��y2lݫ)�R��3�61 ����?�yR����D��Y#*�Ӥ�[��yҀ�P���ڲ��UT���Z �yB�n+�α��a�HJ i!�'X��y2��T�*�J7EH�;����a��y2퀢7�t!�b���͒$��yr�X�ּ���H@���ܘ�� �y�@L�/���)�'�,�%�.���yR���s���s��5WUn�y�A>�y���X�+��˾?�� ���ل�y���'v|�hA=9�иK��y��
>}	��7f֋F�9Fϐ�y�*��y�L�yB��u�:E4�y�%�:�8m`��[������k���y��?$���Z��n����y��Я�X����
��`���6�y"G���2X�!еJϨ��`�V��y��Q�,kt�4c�$��F���y�nC`�� �&�T8 t�ۡ�y"^.��x���4�L\*�y�=S����EF�|��)iـ�y�,J�-��*�/	"�f9�1�M�y,�t��[V�;ƨ��f-��y�i_�bf��1�",>��@b,��y�OUX�u��c0�J}��n	��y�(�"���8��L2P�3.�yr�N�ǲ��鞜D�4$Jӆ���y򣜊E]#U��ZL@c���y��N�Sg�D��d������R<�yRc�Q�S��/^�����y���9g�������~��qv�@�y�@��5ݬI(ड़�?�������y�#B�	���Ċ��1$�6+���y���0���y�χ�X�����1�y��킡�B� F�h���ޏ�y"��8�H| �hR 7'�|jUc���y�O9Z¶�P*�-[��{gX�y���fc�r�J7U���"�'
%�y£Ҍ%�Ti��k�G�$���Ι�yR��S2�Qq�kR�4l� �/��yҢ�5R�N�h၍�Au!K���4�y�#\�`Ny1$Ո3�mJ�$��yB�Lmg� ��F��0��=B&o�2�y
� ������*Y!eC�#���E"OD��a%r�Ą���E�, tj�"O(H9W�bP����ݓ�� ��*Ofl�pB��$��q��� R�<`B�y7��a  
E��)�T!�X�<���W�6|���h��U#���M�<`E(�Č1@N�#Y e�'�L�<y��G�i�8P �;�!	"� M�<᠍�n|p�f�12\8W��p�<��N�Z����D��}�����b�<y�� .��K��ڡD�
�;u��I�<�v�PSu�����K��g	WF�<q�URh�r4��#�(q�E.B�<Aԓtp��\Xu��� M��P�ȓfnH���f8w����W�m�A��)�,�AP�U�p�x�Sc�pNҌ�ȓm�	�ԯl�~E�$M�H����ʭQפ�#�X);�k��u��M�ȓr��uP� �87��SSL�#^
N���]�����׬[�4d���
rh�m�ȓ|_�@��AF]��dQ��� �P��ȓD"U��NܮG<�
�aĆ0�v �ȓi���k�� �x}�t�W�s4��)������\@F��#G�8v86Ȇ�}$��l��|	�8�2)���h(;5W�`���ޱ=n8х��Đ�7�"U�@1#�R�|��(�ȓj�@|��W�|qҰHX3SEv$��Ks���"�"��SmR�P�̄�;�����K��6a6\zB�g������tX5D�{I�U���y�����Tuz���
:x�9��Z�QS���NĈQ��(�6sR�,�a膀�%N'D�4�vHQ�WA�$rը��B���R�i&D�dH �߆=��e��!CͶ����1D�4���v�(��J��4)�0Y��0D��sHPSb2U�fA׏ox��C�(D��#Cc҆;��'���ի�9D�p�t��� �X�ßk�y��8D��dM��I����W���z^E@�O7D����"J�0� %�P�TH ���*Oֹ��i�*��Z��݅<�����"O�$
Ņ>1�\W��=�����"O�!���ԑw��S�UO;���3"O,t ��$W�  9��rF"O���_(o>dx�`������"O����n�?1��ԡ�d2{��}�R"O"��va�;e��yPр�'��7"O�(k�+�C�La�΁(>���"OJ9+�E]8xG��x��Mh~̘�"OR���N�,x�r`��X{�11D"O<���L�b��R'�B�=yz�R�"O�PHe�E�V��G<6p�G"O� ��b�Ruh�u�InI:���"O�Y�a�Q�j���J�"-6�r"Oꍨv��#��QKWL�]�N4As"O2��2!�2#�r�
�)%�ta*W"O�� �%���Ġ��Q�i��݂1"O@��F��^�8�Kfΐ����"O�����!]X�"�L0{��DBd"O�QR��d?j�#jՀ/ˈ�i�"O�Y�'���Y�k���6�\��"O���J��I}������?�H��"Oة�F�1y���q�(O?��!p"O� �4a�&LljL�F�.l@|G"O��!s��T#�E� Mu��q�"O�1�G��B1P����1t�82s"O"e3���$!�0�oE�I��|��"O2��Ū2�����R�	���R�"O�����4$��5P�Ε&��D@"O 	2�i����#.��|`�"O��d�Py8}2уG��A�"O��rR�D[h(�C�gǟ�|�)"O�#�@I<I�:���J�lq�W"O�0�����R׈�����Dh|�Q!"O�qJ��Y���3���\Q�q"O�8[��XG(��д@�nB����"Ob Cb�Q�U�e�_" HXb��y���$P�(G�׫fׄ�ڱ$���y��-	2d�εZ'<y��\��yB���+%�X���e}*�)�E�?�y¡�,�V!Zd� �Q�J ʇ�=�y�"�)��q��C��|)�*L�yb�я�0ѐf	.S��㵧��y"��B�d�Q#�47�D��bA��y�Cݼ_�!Y4�
�/~Z|��Ơ�yr�^�A�� �w�� �t�	e ��yB[.Y4�9��W*kʰ��@\�y�D
�{�V�:�a%a� x@���yB� O��da�Wf%�#�o�+�y��W2,�Fm�4��H$�Ͷ�y��72��iÈ�!��S�Q��y2
�0Y�D�&��$��Yȃ���y�F��c�`I[�+V�Z�:�&��y�f��x/L�i�Ŝ��dT�����ybL�$,�إ��W��)�L���y"ǘ���E���G#Q$,�*����y�&��7#��'#Ès
P�[wD\6�y��V3��T���,|��#k�y����J0�׭�G��}�Rg�y�Ì&g8��1���M�)�*��y�o�!�<��V�L�Ba"i�bᄉ�y2kĸS-� �E��'LT��C���y��Ք5�&U��b�M��483슰�y�O@�.���r�ƱJ�l ��C�"�yf.U��C��Ob:���ˎ%�y��J�b\�ijcB�rފm���<�y"�:���	��H�"�Q�cN;�y���y̲��f'��mx��� ��yr�������0$Z�H�B��y���>l���чȘ�1zZ��A䜖�y2��L��SB��Xa�
@jL�y�ŝ!.g.��5�J�V���3F��yr��-T2e8ѦB4�M#�.)�yr�& �\js�̷$�,9a�Y��yr���dJ��"��6�H:��G+�y��֧�̊��������y�&[1���Y���֙�#!���ybǀ(NȐpJ� 'o�����G�yB��.� 11DCƜ<�A�R��yB.�4t�A��M�#|��A�5�y�� M�|����)/f����'�y"#�g�N�;Əߤ�����Ы�y�I@-}��M��!w{*i�%%��y"b�4$��&�3xLL�Iu�X<�y¤͵H��2�g�h��I�M�y�;a\�y�U��eFz�A2���yr	A6c�b8�/��(?�(��#��y
� ,YH�m�_�]���=4��"O �`EA%T�ni�e[/)����"O�q�Ǥ�lN|�"O��y��P�"O(�p��R�b&@��7.����"O��Z�G�.;�ԅpUO�z���"O[C�
<_�x�;58J�|I"�"O�}#��J�x�T3|nqP"O�ɸ �N�mj^Q��k�af� ��"O�$��)�?m�~��5h$��"Ov �6&]�g��Ңnӣ6PibV"Of�%�|��;��A�;��#%"O��yE�*V�ʕ9��|�� s�"O�*���B��B-�P�u�"O�8����I�́�����)�"O��kE
�%���`$�^���"O��2�w�plj�f�:/���p"O� �b��"i�P�p�-f~�PPU"OD�Ȑ�0��PF�#\f��w"O
�y�	�L�l���W�J����"O�鵂J�?u��Y�8<>��("O*	y'��!:M�.0B�E"OHDi��� ��<K��UeJ��"O���B1%4��T�ʪ&�]��"OPm�&ޯ:Vf}�D�N ąz�"OX� �[:ġBԺP���9�"O��Z ���-��@�#7�h"�"O d�E�j� �ò*@p���"O�|��h�.��L9�n�9A5(<[�"O2-"�LK2��$�� . M-�d"O��2��$�t`#�]2L=i�"O�q	��S��$�* ��8L�qP�"O,��,_*V^z��y��E�f!�$\���sG!X�
ڴU���3B�!�$��/�zg�[\�5pb�|}����
�R��."�4M	 #��0ib��ȓ,J�-!d�\�":|��c�
	$Zln�u(<y$`�v9d�Z(n�pӁ?O��zr��F�B]���W�
(�ׂ�!Cu!�ͫKֶ|+��,7���ġƫEY!�D�;=tE1s�X9R������-"!���4T4�sF���kS��!��H�(!��1��Y�N��]��!�D�h��h5��GX������p!����s	��˖��-���s=wh�z��,�I>
\�Z��e�6�7(1�B�	���:@`R3G-�	2�A��� 㞸F{J~:`H^� X��A��x�Ab�<�(��|a�7�ƋW����5��<�	�.���qo�T�|=h�*8��1�ʓY��1��0�O>TuB�ɤx�@Ca���֩CB�Σg��#<9���?�����NվPi��5R����-;D����
��S�l%��K�5���gX��yb���O�|�ŤܡGP�sҊф_R�T�&"O����&��|���jI��_GtU��7O����:9J������kpő�
|a}�>�P���vC4u��zsf�jJ�Y�<сO^9X����U�o�\���Xܓ�~FGG�O�j���b�#A�$�(r U/��r	�'�U��,���଄'�9`�'ܲ"=E�$�W?v=��R�S�����j��ybI��3>�@3"�H-4�Q�V��y�b+j�,�5�H����p?��O�ɛG�J����f燯 ��Ĩa"O� �p8`�˾������S4w�]�U��w�O���2S�ܧfe��x¯C0R$M	
�'d`�xd���`�a��GZ!<�¡��OD�"���S�P9�K­[en��l�b�C�	6Q��5���Q�L2�Q�쌶��C䉫��x�$)6xN��BʜJEC��<{���d$Y&Eڭꆡ�%��B�+,= ���>��ˑ�}���D�/?Z���k��1k����
@&�!�D�+� H�R-�n` ����'"!�D�` P��T�JnR�ђ���!�V�u�ʽB�'�&K,��7�דl�!��ع݀퉆�T�'0&��<�!�<w���q�;"�a����=�!�D<�8<@3��$<�c�>�!�	j5鵡T�x�Q1�ʒ2v!��)v��)h&H� �����\� �!�d؃
`"�#y�� Z���u!�d�!E����_W���r"'|�!�dгi���a��0K�QߨC�!�}�x���Q/�8l*�h�g!�dՇU�$�D��]�P���D��XEaR�O�Q3���\3�1�%���@=B�U"O����T#< �s�S�h �`1��IM�OJX���!O�$���A��Bn���'!恊�MH�J���6_y��+�O(�=E��N̦%��!\����VgL�y��)�*	�bMS� &����و�y�!�0p���@Ċx��\	F��y"�A�c)���J�X�XًmM��yBJ�#�҅�pE<e����GI��~Ҙx½i�a�T�B16ED�	D��%K4j5��%�?�y� 	�B�h��(s����ƶ"�6Mo���'3�x��E�REv�󆈍5�
���[���>��4�~.P.y����lO$(D��i�?ܴ�p?��g�`�ϟ]'�LC��ʍAn"��ȓ^�H�C���.-�^��k��1��ȅ�R��b�(
�l��TJ�j�E|��+y :e)aFP 0x 	 ���&O��B�#
%T�êa�j!V �B�I�u��Q�@	5$B��5�1�BB�I��"�i��[2:qA 	s�XC�I�I�꜉�	*_�D��ȯ%QPC�	�NF�!P�F�5�F	��E@"pC�	9M10��'d u �H�jC�I� ��x�f �k�$��ۯr�BC䉓!�����ѩk����fW�\pB�I�I�����ت�p̒w-W1/~B�		x��Y�`�[�~�jc���=(PB�	4z�z!0H�V��$gZ�jT8B�"Co:i �H�	�����T�B�ɝ{Dԃ��Z�e�$g�F�L��C䉪	�pt↊�";��4CT���B�56D����,��H  ��k@? ��C� l�����Rg���$mZ�C��>	����7M�  � �K�$^�u��C��?�
��U��+e�Њ�-�AøC�ɰ(��7!�jg�9��74	�C�	)OK^� �Տ|�,a�Q�Q"OVyH#m[#>���¡��C��t"O"�"��UH�,Yr`�A��	3"O`�p�Oς����LEH��IB�"OLu
l��L:UA
o�~(�"O�`��o�������*)p��Z�"O� ���B�R�+���a�,�HX�P�"O<׊9��}`�"�G��LZT"O�I���g<���V�P0=��B�"O����,�0[m���V�#_͠)7"OR@�r�Ed8��HASĊ���"O��y�ƀ�f�~ez���!Rօ�#"O����'�5"��ǀI!9=I"O�5#`�W�;��kDO�j�PZR"O� ������Lz���nP0���"O���7�(~�p(Ê�*@*��u"O���i�4(�AHp����Y2�"O:)�`����|�v��&���y�+F�[� �Z3��+&���MA�yB �<*�
�ȁ*�dٕ�V��yOՖM̒Ȋ�	@�:� �Cʋ�y�KK�֘���� ��b��y�8ix �qRǓ}XtA	���y�/��mh�P ��i�4A��-O1�yB`O:��R@�d�d�BRdB�yB���n@��P�0[�-��ԍ�y�φ+�@ 
F?_�$�ZP���y�@�3i�	�틷%��(��Ǎ�y2MI�S�����$mP^P�S�y�f"@_���R�a�Ջ�ڶ�yHl�FM�ƅC����&kR��y�3e�ë�=q���.�y��^�#�k@a�5b��P6���y�`["� h�0��&�ʵI <�y���6{�!A�$Y!Q,�c"�B��y��Ħkdʓ	D,Z�ʑ`�7�y����L��H����!���y����^(�FD���ȹ�!S��y�
�L�
�;7�ˈv
���0�U��y2/X"jg�#�%Q	W���[@���y��,}�̐���I|�	�w��y�@�%cm��A� 9��pC��y�"%f1�r)׳@�5rD���y��Յ|�x� �	Ο��u����y2�U;�F�(����ֽ�����y�L�� �@�3w�,���CK��y��#�}cg�ڒ@K��2E��y�i�$N�0Z0�7�ya�* �y¢�2�x�f��Ӂl��yB+��\�6�B���z�HA�P�y�oF�F�쌛aB�:��� ���y��
7 Gz��% �M���ZceL�y�
$l�(���Cd�X���Q5�y�.^�R�Rs!C�=��Xuo̭�y2�[?'ƀ�Q�o:�~y�R��y���S��|�B��=~ ��+ �y�d�n�T�8�hVtnU���-�y�I�tIb���hK�����3���y��:)<��V*�Rb�jC�ب�yB��*2|e#p�[���X$����y���C�0�@E�0K�H�8�E��y��9�0)ꅨΩ>_Zu9�2�y�,�e,��h��Ċ1B��c����$$�O1�a�S6`�.<��\�B/�h��"O�
�`"�6Q��Y�5 FͲ��G8��r�E4��eR �ǿ,}�%�B�,D��:�O�e}��r�hE}a��E	~�
Cቾd 	sae�qN4�d+�/?vC�I%/�`� �M�-FL�܆PUtC䉸S$�%���Ҩ��U^ C�)� ��CG���,97�g�X���"O��4e�"y2�qSb�S�d���ȥ"On�Q��.�h@���0���G"O�=�b��*���Ҥ)s����iRB��	aSļ�*�(s������-ih���$��`수#�KW2ȉʵ�#Cr$C�	����ȧ�ɹO���"p���"��OL�����X�W�[�46�X8%eU-zay��	]\��g��S�D\����c�"=!�Bqd�{�ȝ�!ծ챴�
	0w2X�ȓ �t,�:F܍1��� 0��;�rls4��:_�J઀�/On���k<��Q*����W�(N�N`p3(�kH<�J�|ܝ;u���|8�cKN�e�!򤍮	)���S�.}���K-|y!��S����

:&��{lU�o!�D4#4zIg�\�Z�A!+ޏ*U!��5|�H����ڪO�x�0tI�h!�$Q,%���2Bg�E{DL��g�
BW!�d<}V����R�r@�&Z�6U!�X4%��=Y�	@K�:�Ұ
�dM�s��(�Vx��/�"'��I�������"O(mS��Ǯr��u��oЩM�D5a�"O�Dc��)9dYz6�n�r�;
O�6���<@��l��,�8�B���!M/�|x��/u���2�#�qM�MP�@ϙ�p<A��$L�060��b皲|��� [Q��D{*���Չ�|3DY�e�e�F葆"O�DJ/g)�tM��&���+�7D������
�0����b�~ �V@;D� Q�N�mo� �Q�Zv>��0�I&D���E�_�Uþ49� ����u��.%D����T�]VZ�Qf�9�xmq*#D��b��Gv�Bra�;|��c4D��@���wM�U	U�ы�:���h-��&�S�[��}��BT� Q���k���ȓV�� �q�:#�"|pb��J"I�ȓ*; � ��O(�	@�b�> ��N��U�B-%��T��\�	.�Ѕ�^+<e0��%���S T =��	������@�IВi%�'�m��`B��h<�.�0@͡ۮ�&�<E{��� ҩlw����#@��Mӓ�W��y��?s[T �c��(Ed`�Q#]"�y����8� " �7-�~����'O�V�~��'"⹐�A��p���@�C<���*O���K�oc`��9y�8Ԁyo!� uO|A�d^�pSb����[$P]1O��Ez��D���pl����m�T;�DS<ט'�ўb>}x�τ>#��d��Ϙ�M��y�2��66ay�)H�*,P�	BΡ~~�v����yℋ%Y@����Jl��V���Ms�{2�'d�9딋��x��,ȃ!�c��8q�'2 ���?->����`ņc�� ;��Ip���I��f�<8��bJf��� �;{��DE3&e�Qḿl)22w!�|�|��Qf5�S��?�&�0{�5؃c��ZƁ
Ax��Ex�#A� ��԰�)�5z��L�B<�yR���dR�!2�֓ �$hF)����$8ʓAT#<���Ǽ1H�e�r��h�@,#0�I8��O`��NI�2���'�J���΋C.���?	���~�V�X�}�m��6z��!)�hMV�<�6e�O�<=����1���@[�<i"��i���R(�JUP�I\p�<� ���ӯBQ�O��.��D��"O$m#D�-&���bD2p�X���"O���D*�$J��Y#�Ǔ_�b���"Oʝz���q��G�ʣ~/�<�U"O�H�oο8b	p�N4X�s"OV���%ѽs��I���Χu�B��"OL��;i�Zj�^2vR���!��ēBO�X
3S�#���0I��F@��ȓi�x��S,�	���C:eDɇ�'��Qď��@�h��q��5�'^�}���E����`!bl�0F%�y�NQ���� i$-,�p�C��y��a	6|���I�%��)xd�V�ybn�*p���dN�K&��T"�+�y�ꗖ>rС�&]�A ,��#O*�y��7�$����cE�|j��7�yr���H�%�0�'e^�b����y��R ;�`�ആ��K���:�+�6�~���v��h��u�aL_��]��J�>Vx�X��"Oz��tO7\���zՉ�5
�4�BU��D{��i��#��ɠ��2�~�z���7bK!��]�$N�d1G�P����ԫ�DE�'}�|Ö����$](7Ϻ�+�j���y2��*zcp���(�4������y����eaR�Jy����C.��I��ў�>%aD�6�lPPD��V��鈴�9D��Ҧa�)b�X�f�K�:��U�P�7ғ�hO�Ӝ-�$A�BP�]�r��Pa]�I�4B�Ɇ#R<�Qqe�A�ZẤ�#E�(B�I-��,k����\�P�1f�5NB�+2� 8���@xN�뇎�.�C䉃jj����.mox8۲�˓s%��s�u���32�W)jA`���G�8�.-�D'�|�'=�O�`�R�
��3{�U��H���~�H����OB��	K�e��A���(Bu�%�w�ܭYUQ�$�=��yr�Hv���T�խ/'�d��iA��y	:�V̙Tj#D��n�'"��p�OD����_��X�[H�|�:���'Nx�[�A��v���ɦm`��aÓ�hO^x���ZF�I�BOG"?`�t�'JQ��a��F{P�aP�݌8J�n�<����S�X�dDRrH��I��]{�I��z9O�=�~�o�8�>��a�:X����B���=�`�~S,1�Ȏ
P_�]�
Iz�<1`j��~J��"�M(+DQ30F�~�<!�Έe6P���,bGN!{Ň\c�<�W.҈W�,	(f`�%cT�͚2��v�'ў�'O�ЕӔgԀ3�}��Ʌ$:��i���Pt�#��.�\�טa�Ȇȓn�de��'�#��M�K�/Q�ȓs5�%����!�&�ږ���C�ĨD|"���2= ��	7AJ�#�F�&q�BB䉸n$�ơ	rE:%��(�8=�,�	&,�Q��}"�"S<V�0S$���4��C�<	P/X7h@���UD ����0cG�|�<iWAD/���7 B'�\:��@�<����T0�	k�a�Bh ��t�S�<Y�h[�v�R��![� h�5���JN�<���:zZR42g����	I�<�\�_s�]Z-(j����{�<�j�.$DhɊ"j�(~X��2�r�<����$�8KF��9���2��l�<QL Mj~Y�����"���.�i�<Y�q���"9��h��AJ�<� �y��6@�y�Slݚ7f����"OhӬ�*<�4��d�N<�+f"OD���*	�q
R����"O�� ӟaS�h�F
P}4Qd"O�����PS��	�f��
o�l"W"O�)��^�G�$���_$9.��"Oz�y���� ��KOB�*"O��3��*Rw%!���8/>�ȣ�"O"��o�Z����)�<L�%Ps"Ormc�<�����Z6`�,H�A"O(��R���k��d:���F�h��e"O��04O�!�9J���Ѡ���"O�40r� 0�t��\�i�j(��"OH�����&��0Q%
�OzRXc"O,D���@�$rg�X�oq��c�"O�ᤢO6D3R���F�sk$t��"O�!�╅n�dDJ	2���"E"OԊ�`�=j��g�!}�h�"Or͠aûuR�*MG1p �v"O��⬄�	������[]Z�XC"O�!YR�I �H��2f��^���"O��p�	Y�d��"%�1<8��ʰ"Ov���K�*at̙�D�	?�!A�"O&Y�Q
վ ����P�\0hL��"OJ5�T�?!򝀵��v+�iU"O�	�g��+�`�~n�ڒ"O.e;��@�-��
�.T;"O�xQq-޽6*�$��f���+��'�� ��Q�}���bN�;QJ`k& ��q��Ē=Y&�\
���O�<)�*�۬H�d��a��D�<Y���?�>�;`�E>\��=�aȍZ�<)@��q�jDx`A�9'�5�2,Mi�<qG��$~���j�
�#�|�!�g�<����d*B�9Cj� K�#u�a�<���)d��-aQ�PZ~q�CX�<�&fF.f̤�@��küt��J�o�<�v��4g�>����Uےe����i�<)
;��yr�҈M�p�(q�g�<QĢ�&DրA�$�/#sh��e��u�<�V�Af�pxdBG�0��V��<b��946%��,W:8�9C�ϞN�<Y�a�	b�Y� �8Ӵ����WK�<F�*Tp�!'�&A��Ur�H�B�<awbѽ.i������|	z��~�<qDn��6��eiR+�=t��KNa�<����%P���N�S�<q��&�E�<��üp�=)c��81�>�����T�<�q.F��9C�*K3��lat�J�<I�Ɋ$:Z$t�a��]���\I�<��޲k���p"3w�	�N�B�<w�O#q&�eD
�!�8H�"�y�<i3.Ĵ[9B��BJ&Qe ���Fh�<)Ei[-C�N� �g��|��$iu�FH�<q@�[�U]!d�6Mt�rE��K�<�5H��E�I�,�2~�����Sz�<��O01�܁��,ʔ ���I3�t�<�� $z7�Ċ`�/�q���p�<��C*%\�R�EM$~u�`�"�7D��qdϔejDX0�8QNB�A��3D�X�r犫m�b=���C�Z�I�1�3D��7nP�9@r�9 &�-����*O�\q�$J�d���BF.d���@"O:��ӂ��QI@t�!㉶��"O�A�N�(X�4�6��?ނ��!"O� vT 1�x��B��nϦ��3"O�Qh�oY�U�a��ż�+�"O�I1�p�ڸ���<��$AG"O&�Yd O�!�p�;����	�����"O����i�m:P#���;g(1@�"O�5�(ٛBŰ)� cX�	��웗"O.��7ɐ�s�����
��a�"OFp�t��([z����8B<lt�"OBX:#ΐp��Ѳ�W,&'N$�4"O�a���N�[\�D�Ej�**"�c�"OH0��+9����IҼ+��ș�"O^���E�Q|�"�Q6��"O��L��q���Y��\� P��Q"O��H�-�o�pܻC�2R/��"OPh���$D��iǇ�&�i�"Oh�+�i�R@�)˒HX=[��0�"Oh����Ư vՉň��|��-��"Ozi�	�-��L���W��J|��"O�	Jƅ�$�^C���S���#"O�`*taZ�-(Hm��"V�4�ܭ�e"OFt�G�e��Lu�>t1"O��Z���fnn�A�O�;u"O�UpPIH�V�T��d�8릉b"Oθb!HU�x4�p��?[��H#"O�)(��M2^�f�� �G�|�s"O�������A��}0C��.�jm9�"O�9^m�Ȭ��JҊN�R��OB�<�6��0����� zuV)����P�<�w�N�.k���U-�fI@%@�gZ�<���]3Pg i.�%1PJ\��B�<a��s;�����A4��Aé�y�<!�*E�:�L��N �^�|�I`�w�<� bݥ�*�+�� �z����/w�<��(U��]�L�(�zհ���p�<���1g~M��ᏎH�B�P��FI�<�)�&5�)eA��:8kD+QY�<Yu�U�p����iԁf�q@�o����N�qOBU���И[ɾh�en9g(P�(�"O�9��9>� �]�m�* �Y��*p��6t1��&��|�E� �Y+ԍ�'�<<X\�RN�dX���a�[x�'�ld�Tj:9�^���O��O6���6N�¤�����I�X��4�� ���I�_3*�k"�V2#C,�r��(!��'G�H��V P9ɧ��($����.,K����p�0=�C*{;@��Ҥ�^E��!�)3�O�9�T�қ�<��阞T0v<�����1<�l�@6�?$��D*��8�*�gW��>;�(x`hk��y��B+�C��>9�t���2 28�����jJZ=����k%�(c"a�<�Y��U�j�8t�b�3"�Ni���_�(8�1�ў6zaꔆD@��"5�Ȍ���Ә>)4ƎZ8�W�L�R%��lS*Ai�(�� ��z�҄I��މ�8��O/��?Y�� �:�CF���V�@8���G|~�,��f��� �SO�T?�X)�'T8S�kVp��ڦퟐV��"G@��F�Iu'.j��AE�'�1A��;�	�qNz���q�Sy2,F�?�s�N�-@@�QV%�z�h��s@^2�t��®Y�lH8p�s��^}8����A2��54I�h@��ӜU���Pfd�$۔y#�č1.�qm]g@eBM�62M�`��f�G
�9�Q�!y�P��k�,������>@�$rF���	#����U(
(s�@�#G��I�4tچK]��l+p���N�yq��R�⟈d�F�:���Y���]f;��y���s�Z� >���F1�~r�iĲ�y���d�ٹB�n��r��$cT\`21l�4�|�ڢ��OH@eE'�����V��Y`2�W�hb8��80�*�I�@�t�(��/N̉)T!�+O�(4ċ1<��Bфܘ�yg!O�$
��Bó+{|<2����0?A3	v�T��F2�F![�O��G�R$"p��*m �8Bi1���:�����?x�����<	6$�����n�xڗBN�&��Q�4X���:�*��i�:T�&�7%�
o��҇��	}�����8(b�9P�ɗ:v�BL۰��^?���H���kT"�<	W��5e.�j�.1���	{5
�j�wk�EZ� J�!�� ��&�ܠ���C��F�`3X���׈�׎ (BG�XyZw������� v�ɪ또��@�-�:,�@I�
���¿@�\�Ci�$1�N(���w����	��@���8���!�,�&�?a �3t�"�F�6m�:���Ka�'���� �Pq�d���$-[E�R�x���3��4'cj��n�"V�&����Gn�D�0Ħ�c���D�.85�v ���I��[&�$�\5~e��"3a�9(�!���B�4���ǝ�=w��I�C�%��;Xy�4����>G �����=o��+g�܃?��B�	�^~P�#CG5�td�3�hdB�	0J.FՀFjȿ�P�c;&�XB䉦2��9A�<�X�6C=�$B��#5��1j�1O0�0,i-��P��ɒ��8bd��h�O��RW�L�H�$��'H��XD���
�'�A�E�jb��"�$�-%;��2K��lTĹf�̩��韢��SmL����<��@P�ge$�z7�\�u�L���.lO��[�P����q��KD�sa[0~���w�̇nLV��0���
@9y��t�ϓ5�f�kD�B�c����Z*\l8e�<�����]h0uy�ֹG�,�	��B�2ciJk���k���DP���F\��o�xh<��g	�^����P)ZB	�2*�mz����(.L��ɰ-�
��6��T�ꪟ�e%@g޹����2C��l��k	��d%"J%4��X#
F��r�0q��M�f�2�U:5�f�PN֋���T�<Ac���|� �
���U$*��)��l=@��e��	6dP�3��~�>��&a¶��t�&_^}:8��K�q�B�qf�'b�y�'��f��x3�'e��9�&G')I�=�����}�YL<i4�Y $�0�S�29@���e韒B2O��,�3��$b��E�|$Av.��R��B�	�״�n�]��3Aԁg���X�-�N�&p�u��:vFXFO�к�D.��|:�4��Q�;:��P����Ĉ!�+� 1��s�^@0e��=b��
��XΒ³�W�Z���FI,'2^�������?�EA88n��R�EZɞ ڣ�OT�v��,\�����M*p`���'�`�N�L,��AJQ����bJ�/0�	Q��քYO��h�)��,��DhE��D
�g��]�2
�o�)�b	#INB�-.u��	��3j¨�O���C�'
l̼)���!LFLԑ��.��#m�|!��N�����ʕ#:l,�v ��P�O
�D��O੃U�"b�q�a#ѡ<��8�'e��^�Zz6�ئ2�)L�}Xq�O�h�!�#K��u$�1���!��iZ(�8�I�J�L��ɶ,&T�w�K�6�8�J�������S��~�������@`cp��I̓�NH�;�(�d�,�81a��� ��A�̔��x�ĕ��J���ֲVXn�cR뇫�8}Ӄi��BC����6�����2�.=�qj�6�h���0f8B���R�K�W�P����x�Ś&�`� �'�<�b9*��^�'P�֑c��_" ����G A9E�7�@u�M����Y������;���
�/N��[�D�;������9����4�Ƚ'NXb?Oj)�!J^���Ѳ�
	84���Űix(\�a��6\�\��I�ZA�Ȧ&_��W�d�0@K [E���Ɵ�b��XE(�I�A7\	��@�/�n�$��0,d�c��:m�B�X�Ց%�yr��l�H�p���'D4ӂŀ4$���mY�(EHx����O\tr�AC�kJ"~R�h�.C��R��:���1A�Y̓:��)hG� ��"+�'Q��a����r6`�
�:U�I0�7��"~�zW���n����@t�0��G�Јn��y�yRŐn�ړ�2��;$@�R��6/�dA�rc�S�(��ȓ,~���Κ+Q��x�֒S������天25!_I��O5�]{5��~��O: �ی9�T����Y)%B袗"OڭIv���5��+�>a����:O*0s�L�9A��;�+-<O4۰�ԸR�D�څ/ǆB��(���';>J4�I�ux�,�#Ҍ���Ƞjr��:�m��Bɡ�āmgƤ�0�	�P�X��A�`u���c� )�ּG��S�'&X2�C���'�vy��ؘvَ��ȓÖ�Sv#W�"C����(��Xx�a�:c8j�K�D�����s��J���-8�Н��@�%[	D!���(N]�3l��L�rr���0j>�˱@����T�Ƣ4<����>!=Y2�e���K�"M�7a|B��+c攙PM��, 2˛/]�P�s���	���`�OȄ8�%Y�VX���7.ȷ82��%�	&�ȍ1���#����:��Z_N�{dC�;�5�A��{�<������B���,Q 0#I���|��𯍮i�-�O?�� ��v��T�6�����
(�dP�"O�tႢuj`�J�g�y;XL/O֡��j	�l�����޻9'��JuEVoPֱ ����!�˷1Lu�d�"l*T�01��0,�!�F��p˴.�*}x���(g!�ΐE+����Q ���W�^N=!򤁎,q��x�
ʲ�!,ۂ�!�Ć�	k��xuhǘriD�!nłi�!��X�ܡx���"&Ͷ5��-�>�!��7=��h�!��^�L�Q�,�6Q�!��:="�#�dЛZ�2�W	�/b�!���,1����ι��e��;�!��Ԉ[����m�*��E`��N�W�!��D�6K���v�Y���F�[�!��;�3�ѩU�2]���n�!��͐%�d�Q� �v|i eHn�!���5��(�� AUВ)yP�B-�!�DM�]�0zd�N���ivj�2�!���3��S��*��h)>q�!���%_�L�ն���Jȸ,�"�X "O�Сd�!S���g�&h� d:u"O�\h�)]�)�hbV�~�Hw"O�h�/�n��8�nA�W<q�""OCi�t\�#G�J<5�>��V"O��R*��np���߅�@ ѵ"Op��âF"ENԨ�f�O��(��"O�L�� _��:�"��'Q�9"O�P�F��2fG�U%E�T��7"O��f+�#/r����A�n��U��"O0����H� z��X�T"O ��%S7#��g(�ظ�"O�����ֿ�0�B�èfM���q"O��3C�-�� iB���~�> R�"O@T	�͋�c���	KWvݎ�0"O�Qx�d�m���t�R�~�(s"O���!��S�`H#�I؃%�Tm[�"O����AL4ź��i�����"O:L���:E�D+��+"��+�"O������"-@���Nζg.�Æ"O@	򢈄�(����Ȋwf��e"O>d:�/��(���!kV�Rdb�"Op8h�.�A�� 	�I2�`G"O������`�AB�^69��;�"O���R'3Lk���~��K"O�P���p��[�M@��i�G"On�����F�'�yӵi�( #!���1V#R`C�fP�vs�= �I�X !�1"���{��C�_{�m�Wm4?=!�d��d��I��c�\a�1��F�^�!�$�r�u!�CY"jFF}#����f�!�dI�'�t�7&);H,�A�M�3�!�B�K����r'� 5Oh0 $���;���DƁecN��v�A�EMP��Ќ�y""�$k̍*`I ���A��쉇�y�L�F�z��6�>!l�H�o�4�y�Ó�<���f(�_�͓$k]��yb#��_\��ٮ輸hԮZ*�yr���f���2F�·:=�sْ�yRO]��* �aQ���a�"�
��y�Oے=�6<�׈�,����MҌ�y��
h���j��][e���y��	)3`�$��8w+��A�Ͽ�yR�˭Ua�!� DP�m��h���yb�=<zdɦ��f���o�5�y
� .(ѡJZDl�Ќ� ���*O"�AC���i���^�z���Q	�'9X����/���ː�L~ �'�� aD�>Cj��H��eS搐�'���ă4H��\���-C���	�'	�lj�fؙO�LMca"�^4p
�'��݃נUy�iTN	2�਩	�'��0(&�)o;��ˢC���$��	�'�@\�Bӑ��+h�Y���'����(��l���0�����l�'Aİ˒D�.U52 JE@�&}:B�K�'@��9b��68��,�e虡jX��k�'`j�G�Y4-���A3{r2y��'6.�ڧk�U+�Y����{�t���'��Q�RiR�x� ���h�p���'��P��V.u�ƙ1&g_ � !�'0��9̑�1�:Vc��l���'<X���G�8h��~�43
�'�	R�m�Z
t� �K\�����{U 8�ƪV	?�b$*�Ϳ<O�ŅȓM7�)��ǁ!g:��E��_�8���zH:5�u�ك5���sg'���;�r�QҩF�q�Ҽ���*@����6��*_(}�UaC�EԹB'�Lr�<iT`[�!'�`X��݀wu���,�n�<1v�S4:���j�V�͹QDe�<���ݒ'��iC����ݱ@��O�<a�D�x�(��� 2]����ăF�<���8��TJdɁ�I��hQ![J�<� @�ETf��fʔ@4���V��J�<A��-����#nϗ_V���oy�<I�����������G _n�<�D凡N�2� �
C1S^�C$-�h�<!��D%o�q��!��V�)�$�M�<���~q~M�!���[�Ҥ)�m�R�<y�/��T��J/8Q�`A���U�<aVg�B�j��Ǵ��	I6F�W�<�sm"1O���Q���i����W�<q�*�S�o��X���=G2!�Dí44��wgL47�T�#C�}!�� 0�́9f�\/U�|4Z(� YaxrNL1R�~��=q�g�3H�4��I�>�*��*�}�<1�o�-k����jR*oPQ��M�ByjZ)KT��QU�|��ɢzh�2v�	*Fx�Ȁ�SPayr��#V��$��c��z	�%�@�ͫT�( I���:14�(�����ިzeng�n�g�'�:����g5�D���H�L��qM�t��o�v��%��'N��Ye��D��h����?��!��	��-��1�Eo'\d�Ѓ���0>Y�c�^R�� 4d\�s )14�1g:��'�
b�L`�|�ñ�����6n��%��T ��w��B�Ԧps,H�EټRĴ�'�	��,𰨢��v���,iΎ S�xTD��+�!+eTԢf��20�x��5��. ��c,S�j3�㒤Y@Ȁ��b��}���'�D�'���фCN�D���ꡯ�T6�=:�ʍK4�@H�����0*��"���#��'꺍�!l�1p�F��Fŏ�M_X��Oܙ*5K��� M��'���P��ܵt:�Ͳ"�^�`{�0�f��h*����.(��jF玱l����D��'@b�)`���2��G�0+�z\j*O0x��J�?̰��i�^t�ȡ��&��ɣa��>��cq�ڐ'�&e���͠V�B�cԦ�\����e'��hK|���Qzm�" �>$���ņƊn���X���+�S�,_f|��Vo����O��)�}������8�:�*�g=�3�(���"WU2�2�`�<������!�=i�(��T�Ο9�NŲ���`X)�ڷI>4���'ΰR� ��Ӕ��O
آC����Ks�W2>QP���8O��РY�1�t1�SE�m?��4 ��[c�OPT�ʴ�,0���$	&�
�cd煳#>�D���'��qIR�:Gwa|B���4���V Jp���g"��Q�e� �E<֌)`I	�~m]�ː��P��C�Ѽsgۏmq�ᣦ�H&?A��9��z��R&K��\�j�+0dL.Tp�9T�(o�����> A�ɥ9��]��j+y�џ� �h�%�ې[����'��=X�k �	���M{��X�4U�ɃK} �rVa��^i�m��7o�Ơ�ʏ�Uõ�'�@	`D��(X����5%<Y"�'�&(x!��hF�P�' �  	!�	%?�+Ch��N��< &��eGnMxk-D��s�IU�O��k�a2hs��Z2��>�@.^!цu��,T����=����5:�F˓T��l��nS�/��R�mʩZJZ��ɒWxXu"��/\i��d$�?5��5c����_�n��'hj�+fb�#���Fr#ܴ4#�9z�N�=@�|�%�@���O��	�Q���	�e2�Qs�"U'+;̝�T��=?j�`�嘸e)^a���'��O8^��9	��éi�"�J���<g�r%+�0�!��)�bM�8����l8B�	?$<�Ig��,!���"�Y�ކ�Y@��e�;�)§`���֬y���@��|Ըц�U�Qi���?'*|㤥�A����?���p���5�P!2�T,t��ȓ-�n`+"(t5\�[���<ָ��ȓ: (ڄ��'��i�P���mJ��Fz2D՝e���S�'avA0��5{�Mz ,R� >C�	P�(�"jZ�E�Heş ���!�ȓ*���y��4}���'��X���4x~ �@�b����'������f_�-��^aj�3�'̊[��LR�,��'\����J6(�Q��&�!Q�R��7��7��2+ނ�0��.��p���فm��#��F,��x��x�$��+#x�
�Q,�O�5�%�V.�28�u6�$�*���"]���QE�Z��C��0R�h� ŷ,Xh��mؠ=��`��&LL��%Ay��9O��`d'�&Q��EKR�ճ�J̘d"O�`ɶݲGF���,݂t�b�0E4O�9C��N��p�h&<O��[1��&嬽Z2�¼udB`/�0>�p��Ҥ�`Ʈŭhv�e�b��$�FL���M�2J�0��'��1) "�2�x��JMh����$�{��["�ĽXg��?��(�;[M�wI1*�����L=D��� U�l{��RBH��`�*�i�:Z���' �)'�ҧ�'d�Ju`����Ѥӟt}&)��)<?He�6�+D�*����2a��%)@<2ͩ>A� 	B�*q@�YkK�U�|J?Q���t{��k�*ʏq�ZdQpb3D�y�=:�f �hJB���$�͓C*�@��]E���D�&3dJq�p ��;YꑄN�e!��'؝����0x
-P2��t/��D��}�XfO�a����'ET#c�\ �C��n��H8k$lO�aXp��l� ��x(e���h�l��h@�J�d��ȓr��yvH ��� H鐒k ��>)���@z���9�'a<b�Y��l�=X���(��ȓ6��Յ."\'�[�9 ��L/WW�d�J�0[��Y�������"��D���	�
�!�X�\�L�"�l%p��Y.h��˝oT�a�Bm����l	�w�laѳ��,�x�g� lOT�k�aE��&h��<���!�:����Gca�R@�'�tm�fřv�x�֬ƍk漼3�b��u���6�>l���#O�l����r Y;��C�(9�����×Q�N�[d�֋}܍��*ڱI�qO?�I�e���CՋ��:q�6��t�#=)��A2Jn���I
 r� �Ѵ�Q�.uZ��VbY<b�!���:�,3�į
�Ȭ3D�HD��l�࣋��J��>E��E%���bQ�:S�0���R�w::�ȓ{VX8`Ƌ6i��P�'�t�
9�#l�P��&|8Iϓ%JNU�AK�A&<P���h 0��	�'��hs��H!����T���a���fH��Hh<���*E9Ta@g��!;�Ȋ��Y@�'S� [�C�$R�f�����;3��ؕ�M91r���aW�!�$5yx�a9妕��!+��R�.�&E�'�ߕUaB� (�<E��'��� DiĢI�Հ�a�u���K
�'�^0��f]�iD�=�I��`�%�'n�Ȇ�� w�t"f�'���Q@NT;h��C�K+l� ��	�;[VA���iX�� ����a�\�J����
�>)x@-4�(wm)b�^݊�&��a��8D�*��Mit�Q������(mu�q[V�-2��xҐ ��ybLG!GW ���x�x����Ҙh�vR$� l�4�O�"~�I8�rس�LĂF��J�\11ŪC�I�N<�}����;�q�6�Ӵ�<���i��7�p=Y'f܆8�`�;�)���%��Ɠm�<)�!:�@Y2#3M�|0���V�<�CZXj�٠�_�rc��f�_�<1�k�E:WH� QX$j���u�<�Ԃ�$%m={í�'zTn-JD�q�<i��<2Y���6����c �q�<I_#���ѯ� 5��dx7��g�<S�ѥE��u�-X?y>�a(�`�<��I
!h�T�!8���lY�<)��A.�@�{��7j���d@B�<�1�G�\8�giL�c�Z큥G�~�<�7�ë-�
�0�M��B53r�Wy�<�SM�6Ǧ�h�D�x�tU8 dAa�<	�h�-���cbL�+�hH2CH�t�<1�)�)ɥe�{�=��d�]�<P��O7N����F�����,MU�<1'�Q�:	BP8�ㆌP�ܬ���u�<) k֡}t���@W�l��أT�@Y�<Qcʎ�
;� PFG�]�#�
U�<�%bY�04dA8dF�	 p8��}�<1��_�1��gI[�v<cAc�<��ʷDs�ػVE�V@���w��f�<�U��c��8�"B�K��Z�m@D�<ɖ��V���H���F���q��F�<q��U��"A'+\��DG�<)�F��6�������	\)�h��C�<�IY��4e�穝-D�Đ����e�<����wZh#%I̫6��Y�a�a�<���/�h��,��8&�ID�F`�<���& ��7�+���ʣ��d8��kVC7	�v����N%4��Ui@�{s,�:NxF���W/�!�,] ,D���:m��X��؃R�!�DV �`�cP �:-�"]�dn�6�!�ZH�lS ��+N"�J�,�� �!��O�԰�E�H�|q��F�O�!���0i���� 6z�R�C�!򤁞K�^�h����%$�횕��-L�!���|���#�8�$�%h�qO�hFz�D��ME	G	I��c���	�Qr���Cu��a�1$K��q�p����O\�@@��#�M.KJh]s����)��+$��9��d�2A�\��O8��QK���$}ʌA`L�^�t��j�>��a��Т$��0|B%��J8D��j�/.9<�q+T䟸���ĹL�.���Cӏ���S7����E+leAq`M�$ފ�� M��P��F��$ح�0|ʵ#�;;B�@.g��,�f�F�p�����l�#i(U��#o�`�(Ǌ-��+��hBD0q�z�Z���jB�e����V�DS88�,=�.dz�/*���+T +48�[��ݮeFlRY�@Z�b� ��7���zf��'�MG�4G.kz�
ӤP��`]�eFބw�!��&Ǩ2I�ꀉ֔Xb�]�	ç/���fn��ސ�q��S�on��B�
l�z��	e.65;�fFO>eie��	h-�d�5!9|���DF�TrV� ��M�L3�C�*YMl����F�(�t��w�,T3�e�B�J�	�!O�pYwOB4qX�A�g�O]L��mT�c�>j���\b�EĈ�N��k�t��-���$�0|�@@ء��-�'��:Eg��	 �:��܃xf1��'p�I��S����po٦m�l
cB8+<� �^���3�Ќ��'�dz�B�*a	�=B�eE.+��!��'�Pu�%�0@`5{a��$w�|(�',�U��o)� z��� p��{
�'K�%�Ri���Ժ���!oζu�	�',&!�۝�:�&I�d4�	��� �A��I�/fL�q� lŁj��L�'"Od��A�~}�]�tm��'?���"O�x���?3�����a��8�"O�9��Ҽ*J�@)��QD�j�"O��֯�\� "�Y�T�6"O0aZ�Ό_��0ȁ��svpU�A"O@L��[-�AA���Ndtx�B"O��G+S���#h˱k����"Oh8��+	�y�#g�#.`�Ђ2"O����� YB��%Q�,z�s�"Ot�J3��[�R�f��
$[�TY�"O��҆4c�b��F
�	�zՒ"OHja�й{�����Tnĸ
�"O�u)�-�RP�b�Ƀ�7�HɃ"O����7!��XAt���k~h("O.`k����FE���b���L0��r"O\��nߓf��R-X�F�
�"O(`�L֍����G�k��8zs"O��3m�;o�^|�e���f���Y�"O����ZO
��Ιg�<���"OX�[�fr�
A��M�L<q�"O8P��H����rqJ�>��Zv"O>h�`F��<��3���K(b�{�"O�����ǚ6/�D�'!Ҹn�"`;�"O6�3�L�Cd\��K�4���"O�|�Q�G"|74���RFRe�1"O�U�$� e��-`��2l�R!1�"O��"P��/_,��� 1P�
�Q!"O�)�J 2P��S�F�˒�"O8DK��@�m�"�@�,^��A"O�)�V�@���K�0GY�Ur�"O4(
0*�! $!y�;`�U""On|����Y7�����G�����"O�܈Ǌ�%}�:�0���D��p*�"OH9ч݀~`��C����\�h��"O
���E�J{dD�rLA�_0$��"O �i�c1��$N���)""O��C�O4Q�$���X�xT\	�*OB�{E���n⒍!���3mtxi�'�P˗ETXRp(Bk1�&���'&�Y�"�]�Z�Cm�u?�yc�'��e�����S�zE�O_�r�\�' �e��0#T��F��9!Hن�
���AL�����C�[��ȓ<���Y�� JI�[@�ޔSg}�ȓq���׈�)0<Jᩊ�Y��ȓA��������N׏]�J��ȓA*��֣Ĉ;t�)a�-Y�9fj��ȓW�������$M�8�)��	�^��h�DT��/��r���	���.��ȓ�B)��Ŧ{���U@�=t4��ȓ.�=��g�
S� �&e�7Z?Ʊ�ȓ/`�	c�
	RQ�a��S�A�ȓؘuQtG�B�����͕���X�ȓZ^����ky�24��Y��!򤃘D� ݊6����*�h�!�dL��i֥��zs�$$I�/�!��k� �ۗ�(I[�I�mE =w!��M�P�Vt�bLW�V�@)` �!��:��Ǉ2�B�KB�Z�!�d41�B$:q�T32.~!�iº(�!��R�k1(P�����Ui���H�!��|<�!f О�>p�e˕
�!�d�QK�IڗZ1�d(���k�!�� ����e��r��b�2O;~j�"O����c��F���3Ԡۦc9��"O�$�3���y��u0�-8,��"O�p$�����*�In~u�S"O��F����<2T���)_(��"OV��G��_��`2g��SYx��"OLt�'����51Ɯ�^�vI��"O<$a�K�{�҈@�'
s��@ʕ"OJ=ha��*>�X��v���~q�Ē�"O���0��H�$)���e��y�'"O8MP�m� 0}q�dQ�,p�R"O�����@�P\�QC&K�h�xX�"Oj`�V�HR�\Ds�DK�I�iS"O̰��hۆRE�����A9ވ�"O,�(Q��wJj���U�,&]�0"Od}��K�A �Ԙ���7�@p��"O�=k��
�=CL�9�oV�JT�1��"O�8&$V-7��=2%��'7Ef�)�"O��:��E�0XR��g���>�,re"O5����j{�ɂB�=�`E�E"OԘ�1k��
���@�u[T
�"O^�
  >l	`@#�n�eZ$"O�PI�,ғN�������	���"O���gH?~��-�fg�6.'r"O��矎w	*�jAHے,Y�"O��85���<��8��&�
bf�C�"Od��6��t8�xP@��#�v�P�"O@ِ�%Y�� ����/�M� "O� @$�,�@�0#��2M�"O<3�.ON�"��OPXqr�"O��2�OՙqE��X���i5Xuг"OZْ��J�\��Q!�I�1�y"OX��B�qQ�5�a�̚)�c�"O�Уt`
�>)��S ������"O�#1���cKNܳ�֑��=��"OJ�Kf)������jR#ԲG"Of���A�\��A��ӃC/�q3�"Ob�CsD�,f(&
O�;�9��"OܽQF ��y䦥��ǉ9<+r}�"O`Y�%�٣xc�H���]�,���*�"O�M����@{B��s�Ñ5�D�r"O굂A,F�ذ�i
Jn��z�"O:p�d��qӠ6�P񘁚Q�<D��*�b�"�h|���ˉ`$���<D��2F_S�I�6H�"�~e b`;D�4�v�M�s�Ɛ���Ŭ%:B�X�E:D��+dDK��U�Q	� p�(C�A<D�(���\�F��ĭJ�6K 9<�!򄖎߆�+��4e?��G�7C�!�$S ?%����|=h�`�DʁA.!�$��Y�0���l�#1$켪�C��0!�䞠{]�]۲%��8��B#Η
Z!�dݽv6Xih�"������^1R!�D��8�P(׭��?�Z|j�I?!�$�,F�Y� �K�F�Z�!ȤB !�$�kr��2E����d!�(}!��[l�����-��ep���%A)_[!��F[f���j�f��s�X!�ď0�dԠ`ؒo���)��X`!��O;N�,9`��1���c6��U!�$� mʅ��s�l$:S�	*O7!��(>x��-D�?M8!�Śi!򄛫��1W�TVLl��@#�.P!�d��-D�Q�e�9M�����A;�!�� ����̐m�
j3�U�.�&%"e"ONY��X�7F2&�Y�R�R�C�"O��z�kU�' f둭��&�}A�"O���I�^V<<�6�
u�X @�"ODԓ�J>���Y�*�.��4�s"O����� �pr@c�gl��2"O�02�l���� vbD�7z���"O 0�`&ܿjw]�e�4D��h��"Or4�UA�� ���d��e[��:�"O ��� �R���WBQ�L��"On�8&��=�ƽ��PY�(鷏�K�<���,e��hA��ѽ=$���э@C�<��lS0�8I#��5bS5��E�<���J����2���0�Pa�t@�x�<��#�>�8��dB��xL��&E|�<�G�R++��-�A�ʃA�r�:f�d�<�&C\+����cD�\-�K�OF�<٦�H�C�̓ЎՓ��q5�E�<��%�u��d�1ʕ88� $c��G~�<)�/�(�Ija�P�j�t����x�<���XG�.-񢣋�*:h8bv&En�<� EC�I$l�Hs/�p�y�O�i�<��&��c�E)7"&xQ�}�,d�<a�+* i��j��&�@ �b�`�<!�%�6���كK���LX���g�<��!o�j�K����Kb
e��Ba�<��	Ё;��"TDJ^d,s#�\�<6FE+ ;��K4�<CY�j3�t�<y�DϜTT-��\<V��1r�&�j�<� ��!-��T��`ˍ�0�Rđg�<QLA�:�Ƚ��
 ���	"i�a�<9ዂ�9lT�DϊN*�Mj��\�<�,]A�u�Fg��ht�q J��m�!�8F�ʭb��݀IjT�6��/�!��Ma��5ib0$Z�"۳}�!�dA�a��P֎MC��[��J/�!�$��K ��T��\�(C�lݮ;�!���T'�`��H�5��Ժ��V�{�!���'1ppq7�S2f�ƜiĖ�%�!���4�+����CPh��C���ȓ"�7�C�s�Xs�l��v� �ȓF@���u��r@��7�?]�F��\y��j�N��P_v�"��@���2�x�#��[���A���j�T$�ȓ�B��˫t������!Ԅȓ'����A��3N��pcI!74̸��!�qۖ'�/R(�i'�F4�b,�ȓ:P	��֐h�<�Y#�H&y�~�ȓ8[��J�  F&��cF!x�<$��,Qz��"J�[��KUlO��х�g�f)&kN5)+p����h%��"OV;�H�%BL2�{�Zs���"OV(`�J�?gR��r�)P� *�"O�u� �8jd)���,!��=8�"O$���j�Y�l\�v
ʧf�^�)A"OX�[�f�j�s��2=Q��"O�Y�ƣK�Gh�p (۠b�й)"O���qf�k���i�	�$�Ʊ�"O�U�d�?9s�C���`&����"O��K�
g����`�?^���"O�M��-I2oM@��Щ�0[��PJ�"O<�+���_�yh��M ����d"O���	��jf�A�(,f�֜��"O���c��C<�|�v(� �j�1G"O� *����`�J� 獫z���Z��'#��ĳM�\�lZꦡ b�=^C��B� �h���?�����|���!�X8C�%?1���(��;CAX$�ʄ��F؞ ���b�P����+� �f[e��Y�c(ăC=n�pȕ	h|I�OW|�'������?1ڤG�E�䋞0Rưa%�̡�Lr����OVʓ�H�@e ѥK�X��̋��՝O���p�
O>6͐'n�t�!��lM�)����%+�V�i(p6��OD�n�՜}jߴ�?�(Oj�'E����g�#e�0i�JYۢ�Ⱦ���I��J� �}�	��&>���,כ9�L��e�����XB���W|�<��5�'5+��A���FN������c�b �>i!��ԟ��	T�q�t����z]p �9f��fY:y��O0���O>˓B� h'�Z(`��@�Ý�$��I��MC�����Ђ�|���P��4#�`5:�U�W�˟��d�<�O��'���i⾀j7,ʥd�[���w��RG���Iş8���|"��X�����N�l1dLפQ1=]�Q���3n <��ʬI$��[��]R��C󮜻z!H)4c٥^i�����Y�u��۟,��4�?I�c �g}BjR�)��Y ��@]���3��%N��D�<y�Y؅��ö/��mI��� �ⵤO&�I��m��֟�ش��I�Ov6� 6[%��e��'c�@0��D�0�ā� �<9o�ş��	�x$��S��I��P=#���{��-Wth�$'�$Mc�	�����cEU�x������ߴ��P$�R�J���S���`%�^7�|	C��io�1�����OP�O��$�OHO6%������s���L5�zR�>�>Œq0���?i�>�Xq$�	�đ���'*�'�7��O<�GoN�!�iÛ��Q�n�Z�C#�xy���'Pz���OГO��O�=+�+;񤝒9�T����:%�|-��a���a{���q#KN3wI�Z�a�!b�L$�%��g.9u'�;a�n���ɆJCb��O@�21�&c>(�!�Qv�p�o�
���柌��/�_�Ӻ�ϟ�`"����*�>��P>�3�"O�%�a�^>9@1@� X�(�T�Ę�MC�i8�I'��� ش�?q��tO��X�4L�Qd��-~8�ᧃ:�~��'rҠWx�'s��@E�MЌ)��ŉ'�\l����'�D�C$I��z��S��|�!Ef-`vF�qJ�H��$܆��'�J�h�'8(h�7�֗NT�쪀�D�~� <���d�O�=��#bF(��w!)zВ��Jj����ϦI��4��$�[���p�fq֦�g�35����O���!��$�Sa�q� @�?