MPQ    r    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h�]G���|I,N>%�
ֹ�I�<_.11AQ���F��IР��^ʵ�����;�)�31A"^�8X*�bB��N��՝�Nb�u���l4�.j�Y���<�=uTG�%�3�4�j�����X��P���=���&u���"�f'��qz��>B3*%_���:^�}�kT��;�v�W"�2XBŤ��T��R(K�j�	_�~�;	�{�Se�"��F`kb|b�[��֢�d�����s>��q֟�T3Ϧ�gͣ�6A&�t�P��3�N(Zށ�~�f�J,��*��GBj!|�l�yw�P�S��O�a�&`/Å8��x:���_(��t+����6F�pƸ
�{�6?M	��L����-��&���Ygu04@�+`�-"\ba�O��+\�iz� �8Q�ey�
łL6a���p���ҬƆՠ�H@g$�0X�e�H�ζ=$E<~|�����1�'�MKB��p���|g4`��'Nr�0�bR�ͣ{8�聡��x}V�}5�9NYH�_��!�^|�� ��[�����!�9���T�@�֛�	���%ܪv�'1�����R�f���|��!3*NK|�`���ϵy�u����%� ���26+.��K�k����똖|W�Ԩ�,h�Ȯ'zV������J�Dl��o�Ģ��s�m��K�����0<���K�c���@M�[���N��vn	��v��X�C}⟄P)n�i8�fQ�������է�tdic�b/|Dz�[��S��y���ў�^�(��p�b5r�j[%�ȝ��M�>��N����{��w�tT�w��vFJ�/�,}��a|<^W�E�*Hѭ�p�<��:��R��S���=����c�p�����pr��He�Jȏ�������빨os�&����g����J�0�Oltt�
�\�s��&6��miI��������$b*N�lͬ}_bO;�^	��@H�� �ݧ"�G��N�qsM���k�QEU�6I8X�����'�b^�7�4Л��{o �
�Aph~]��B��z�!_!�}D�>�7K'*�3fbx� 1����R�+"��<I���X�C�֭lun\]0u������s�κ�����d�l�Z\����5�'z�L$��~Y����71�<�@�ڇO:��%��`�#��W�k�9�!��02�Q��F�V�/�{��W��L�E��]<�:9�=������&˜��fd?��Jf�nR��4������Y8��6ͨ�m�����]t.�� "�,K�}h:�����uS�����0~��-��#s^���D������.�t��rV�1��~�̴�5��
��$�t�[G��u�x���5��QѺE~��,^�l6��d>����+���;�Vs{��w�����n���[����חLK�wJNS�b�����>�Fs.n��<M�Հ~X*��Z/F!�`���<��6m@�θ�␌J���_�h�.��lu�(���Fz)Yy�aS���$�s"Ng]:��D|X�SoOa�KZ�a�j�|XW{�0�?�2��!�T4�p���z��zW��2�hf5!��7�q����D{�㜈Y�V6�Q
�mHm5���U�U��ET��yGh��#�e�r 0��2��
�E!��YĤ�hF��|��~��4@HB�73WK�4�so��	itQ���9��)`�E���ԑ¯�e�1��&�,������+gJЭ1s��x�M�N���ɶ1��@��M���V̀_2Fɋ\��
䠶.n����yL"-��%}o�*4Ħ�����}5���>f�ŧ��u��"�Ô�ᶸM\ͺ���m}�	HEK�����A.�s��#��c�)��}���@�̼
 $��[��L�5Ӿ�]�������+���������e׫YE��U���ϱ�*&�6�cE���}�nPK���I;�R��"�f����"���؋~�����i�_D�\ �CZŨHr��})�b����r�$簐XwWh��j��k)$��y��)��F�p��)꾠��G�ozjf>��|����MV@j�+L����g4��K2��GJ@}���\�[	����$�h
pe@��MB>ր��p�ɧ|�©���U�X�Ax)���?��GZ��j�TFz*���.%_�a�L�}�R�8
-��"s'�d��.W���3m�R��J�@�Q���E�|�x��i�$xca��k9?���`P;~�ÌNBC��L��,��%��s9�E9AE�U�m��)��l����<'/���LBZ��p����i�e(�>�A�"�P��/�f��.(U���D�1��7�Bʥ\��-�Tz^��-��S��3���S���#�M�O��L�2����O0������}��:���(�������>� wEWs>��)ȫ�*�	�G�4��Ѷx�{�v~�qpl�X�ߒZ�;8��j�X߯aK�Ⱥ�
�k�!]X��Z���f�UIE%�� vLL~φ_d��ؠ�[K���)'�v%j�me6�l=���d�������l�Hj\ꂎ�e����Z��L����ߠ��cx�z]��-��ɖ��6,�V�^�����#�1�=N(�ٌ˘����f�3)�̷$�|ԲD�l�B���Z�:������sk��ܺ�hZx�)1P1��RQ"�|A��4h���S.��W�ɉ��<����WA0&3�d1y����>� q�p����.-$�\2L�,t�BDg��Cl`̒�v=P��u(V�o*����a&y����k{;p���`N@l�S�/Y���E�*<��	�+�wX��IB�e���{���N
��[LR�I?�O+)jҔ3(��/ ��e����$�zQ�K�`��t�np�v���8��u����y�I�`�`�l\��to!	3=Jv��XH ����):-$ +N����B�Z/ �d�طTk�l�O��)�n 8�W�j��Nf� ��zIߠ�o���P��D���������*k��Ǥ=С���e��NP����"�W�pakش/a����D*ke�{�,Ls��n_�&���C/�[� ��XɆ�{����֙ �S��Ѯ�2�,||*��z�I�'w�����5���2�F?j���;�9���$�~=�3�a܊�cq�fzI��k�f��˺3EI��	^�>!������ev�D����;�_��T·R�=j�K���mП�-�{��}�����Q`�\�b�n����V��\3�>�J�����a���gH,,6��t<-��o.8N#���t���!��,t�*;��BEd�����w��S��(���"`�	8�=d:��e�jM��И]���^���xp��㖀�?��t_��L�h����S&�BIYc�Fu�!T(ۃ��X�\� �O0=E+W�z�I8�8�!����];�a3�pf ���0��H�֯�K���n�P-$�a|)�����1Z7M�E��-ڂw���T4��f'�Y+��RR6�X�ު��]��X%a9��|Hwm ��Ǘ^� � }稓���7�����-��T���֖|{	Y�%�F��B"�2v�-6s��S�����]I*�Z�g�$�	����:cu[���1� �w֞-/6�L�QHk�z'Ǘ��W���	z,���"L#�_�a�x(��_@����O��N���,�r����*m`�����~G)���MfM�L����fviq�=�RИ�+C�'v��=2n�_����|5���Q�n]�b��d���b���z�����³�C$����nӛ���p���r#�M%y����M����N�t	��cr�2�8o~wooF%f��g�o����^RH���[\�T��<��:r�gR^̞����c������p-�2H�8�JC�����8�0[@�
�0&��Ӿ�ԓ��KO�#~��'\5�����6��hi�LR�N���Bu*)aSl29_�{4;���T H� ��"k�TնC�q���C�[�L�X��3�X~Q��0�L'g���iX47�r�`�A�}y]PZ��"����/��iD6�"7�T�T�b��� �|���q���Qh��GI4m0X�#֨Xnh�U00`��oi��u�Ε<B�zd�1��U���T5Z���g�R��4��.�l���k|��	:ZM�:�z�>�	��س��!¡z0�ⳮ�FGC1�W�{^�~Cv� �#���$<P���U�0 �l)e��_��e���?��:��Ϙ����RФ�/��b��2]O&_�W;���x].?:���S�J���~����!}��[�սK�o���ҟt	,r�X�����г��QK�z��vs����Z�(5����Y��v�K^�{I�S��ub�+�X��gVN0����쩤�n������n��:Lf�bJɲCb�e��=����T(s)*��Q��PXE��Z�� �������6h��'�G��!W�_^^o.�2@l�<��b,Fud�y�ҕџ)$ˢB"ɧ :��o|���o��KU�v��G2X�0��2t��/���I�	�@�'�K��#hh!1��5^�7H��RD�Q�#��Q��Q\%�m���7}��ψ�#�T�A�G�8#��@rtf?0���M�
b����{Y��h���w�~�@�,�Rg��t9�NMċyt�]��4�
)��8E=�FԬ������x�,W8�$L�����J+u�.ƻ���n��Cŕ��B1���@*�̾�V(s��w
r�|��	��قKL�7�� �6"H�oǬ)h���q²���s�L�=���"�Q��4��h'��9��mX�(	��9��^��x�.?�l��z�c��ǿM���������e$�Z��ِq~���C�����j`����:�"�}I�T�c���¸iĤ�E�w����E˾��P��3.?nK��^����;�~��}vf�)+��ve�~�����O\;;(Z@N�r�o��E��Y����_�1;�+h*	�j1�!F)2�&un��""F�&�ބ_/�����	o��0>jm*|K��_�tV�����إt��4з�2p]�Je�>�3�D[_�V�$hŦL@�B���ȧ���F�]M�����Fx䵒�Z{�G�	�EMT����P+. A,an�}�R�m�]
�/�"N~�d���W@v�3ha!�5�2@)�.I�~�S�+i�?�x�E*�f����7�P���ç�@W�'a$,�1:�Iú4،9���U@���ϕ��\���S?<bp�/����Z�Z�^A-��/ ����@LA؀�P�� �*�f)��(���c�����A&\JI"�O�3�]-�:���_�/}���|� ���
��G�U2���
J����ʀ2o}��*�s(X�����>p0� 2�sY9�Ϥ�k����R�{4SU0�s����",���s�3�(3���쥀��J�C�Ê�
�d����mI�(��U$J��˱} �~�!����[��K�d����v �Z��=d����x�ݭ�Tl0��j����i+
�SDɷ��ƓG�� #���.�x/_*z���-��������V�Z��	�(#+��:*N�V�e��|_Zf���'^��7FwD�EB7�qZ��ۜ	�я$O�k�V<�:�x�&�PLS�R�h������ʰ���.���t�X�����!$W�x�&�sdlfp����>�"qޗU�ɶ���\�2'Jt�:ag��]CgS���P��z(q�*P�}�<.
y�G�k@v���ہ�`	i���/��� ]�<ڬM�ơ=S�kI�Y�ec�����.�$�
���L��i?Xr�j-h)(t� ���K����Qp�`D{0�i��vJ�58SKj��������;}sP�ll�3A�^�!d;�=� �s4ʆn����$[e$���q@BL�3 nD3��+���Q�ʗ�)9�8%Dڶet�N�Zu�^��.<����^�;��h7D0�^����2�
��\�X}բ���#�0*�7yM�R��s6Q�o��r���.e���g}d3َi@�&@����:�[ã��K?�1��S_q2{�N,[�	���`�D|E8�z�쒒�*�����ţ^��y� �T�y��t3=xwٜcP���Afu���S3�`x3`�ۏ�\D^�����X�����v�Q���5���T:��RP�j����
��qr1{��V��d����`�v�b��[к������p>���U�.�ʮ��Rg�ԛ6�u�tw���
I�Nm�����_x,7di*��B �L��V_w<S����<�`�j8�X:w���E[F� ����
����,	p<v��F�?@:JyL=,�c9�&�/Y�L�u��<mVX����\���O�c+R��z^��8���S}�o��8J an� pK���V���4H�f?�fF[6!�
-$�X|�7���s1�f�Mx`H�Hx9��,��]&r4֝0'�a&�<R�b��cN�;U�n^v�359���H�y��?^2�k 8Z�#(r�O���N]�hՐT-��֑	��Q%R��]U��������ȸ�D���{*���"�]�$�Q�v	u6�"^/ ++ �(<�6����"Nk���$ϖ2���A8,��z�>L�
��3���z4׊eoG���o����?���C�cɄ�\����&֚��MA_~�jA�K�Svd�U�O�S�C��zK�n�õ����w.��w���,���d��1b%�zvM��%h���A���v�ɰ9��u�p�br��,%TΓ����tC�N�]3�Vl٨��	jw�]�F $ӄ�O�ܗ�%^M�R������p<�Xg:��R95���Z����c�N��80�p��hH���J�x,�n���kꚨ�@�&� �y)��H��fc�Ob��shW\p"δ ��6��i� ��	D#�p�9*��lC�_���;�����H:�S (�"��7ՑXq�m��S�G{��=bX9�#�K�m'���(�4F򟌱����dA&��];b�=������d�Dq�7�"wŕRb.W� ��^��Tv�������Io>.X�֣d�n�R�0�V2�8=R�i��p��$W dJ�E�P�qU=�5ĂvI�t�ڱ�z��Gr:�Ы:�.����x�Y)��M h��=!���0h��U�F�O���{-�V���+��}��	� <�cX����7�'L#���q�\�6��I��B��j� ���,D���_r֨�ߪ��;]*>���&����s�[���f	�S*?|��G�~�BI��?������V���9��@�(t$g rL���:��*6Q�kM� ����]`���������yy5m�}�0�,�]�^窘�wa�0<n+/�
�1T[V)㪔���D��n�ߜ���b��L���JD2�br���xK�t�s$ص�y�U�K@�X`�^Z%���(��b5�r��6c@)�n��� z<)�_�s�.���l뜫���YFp�y`������$�_�"D�:mj�|�c�o���KP�g� -HX�|�0p2}��
���<ܐ��H�<�m3�h�L/�P��7�>�w�D��|���QL��Q�`cm����R�~�K�p�$T,�0G��#�S
r��90W���
�>��e#�Y:��hL#��r8~t��@�Z��m�;AL��)���-~t�G~�/��)s�E����� ��[���z�`,����������J�\u阪�8�D������1�^�@�F���V����ᓋ��� 5����k�FqLXb��Y�}��:XB�Dhr�sI� B�����"Et����Ÿ�����m3��	�׼F�<���a.�z��y�c����Ȑ莧���2�_$1s�����/���P���i
��NᚨzE�u{n���Oyh��\�$�{�`W1�,��E��hድ{��o�nFO�lȓ�h;�U����fr�X��7~ ��b
���y�\V��Z��r��Ҵ�)��Qq�����ڛ���BhEv�j���!I��a���_��F��������<x1�Top�>E8�|����֔Vb��ᬪ�/l�4���2��J��-�y�b���[�r����h���@2B4�����4�? Š�J����x����u�"GPFl �T�覬�Y�.Cah�@}��M���
#��")�|dF�W�3c.l���@:!A'��Ē�.��i%�*x�Jc�aIV�E�YP�c���8^b�.�,�����2/;�9��lU���,���b�{�c�.<��/,`�ψ�Zw������#�~�[oԥ�c7A�PB�_�%��f���(�8�[��'����v@��\��.�J��4Y-m�v��9����Ҧ��;V��&��B2fk��Ń�(V����|}\��	�7(���1/>��O ��st���g���Si܍{4�F�n�i�,�x�����R������5����ӻ�zJ
]�~ȗ��5����1�U�n��rj ���~������^K�)��v۔���ۗ��͎�����Y��h�HlK�DjRd�D�Ďm�Nu�BB��[�ؠq�txJRDzSGH-�:&����l`V�v��p�ְH�$#F��'�BN�i��AQz���f��R��$�����D��B�leZ�\M�D�r��-�k���b+�xSC-PgR��]��� �5E.������'��ǝ���+W7��&�j�d�sV�8B_>
5�q9߼���O�"2* 2�?tS�g8��Cbf �q;�P=U�(�Vh*����V\y0<ވˊq�m�6c`ı@�7�+/O}���/�<��a��N/�I�!�e�������
m}L��?�����[j�[�(/x4 ����z2���VQN�(`�F$�d�6v��J85#���^o�1�QV��l�j(�h�!��q=�?�̎@������2$���B���F
B�#8 )D���"��b,g���!)tQ8�PY�`N��`颃I�ߖ
p�9fV�٬D�S���xF����j�5�sJѢ�D��Z.G�k����[P�M�R�+��*Q�*�
�:��ex��������dAP&�ǒ�fe[�F��Eǆd�Ď����I�$�d
��z�|`��z	>��XJ�I �k2ȣ����_�47ʈowK�4=S=���
��nfp��!���EX3{�5��C�^��8���Tȗv�~
�C]/��(TUL<R��Ojh/z�/�9��G{��9�3\Z�F�/`��[btK6����e���>��ְ���� ��g>��6�M�t��C̥��N���*0���X�,Rt5*1�mB�I]�5�w��[S�;Ϣr��``�8T:�AP� �-�[�՘��t�"��G�9p�����,s?���#�LP1�����&� QYFua� W���L��@�\��Of��+MZ�z��}8��n9����yMa���p��P������Hqӻ��
��_�_�<$�c|_� �,�1��M3��c
�x��8��4�.'��!�CRݢ�)��Ҹ���~8�e9�)�H�r���s�^�Kl �ho�>�1�-�Z��)���T��֌��	�c%�ʹx�n�(c���!�
���U���4�*_����4;�?*����u�]�� ��a�#�+6<A��|k��Ǎpܖ�O�Y��,9�W�P��\���ӌ�H�����<F�${�ר�K�� ��E���[��%���M����������v_�}�&l��jC�ە��xHnp�<�ZZ��߆�xX�$�<�؞�d��b���zQ�d�:�p�y�Z��+��$�7�Y�p1C�rU�%/��0J���<N�fY汔����L���welJF�}����2^�^H��;�R��L�<��T:hw|R�E�X,w�R�1c��`���cp�,cH�J9��I͸���ɨ@��&�j��x"��J���DO���NGw\��鴻�_6���iZ��ģ�%�8t?*�Thl~��_35U;���
�7H�k� CD�"ax��l��q$^�y+e�BF��GhWX���f�V']t&���4�ͤ�L�x�lA��]�;��X�t����D��j7Б���b�� Otk��W������I�/�X�-�֞��n�&0�m��S+c�丿�Kޛ_S�d��K�B�t5Ь�ĝO����ڌ&���)���mx:0k���Z�t����G���If!8�&0v��xF�{�`�8{H�"�tHm��_��D�<�(L��J��|���s��ל��o���kN��������G�@���#��]v��YiT�y�n�6�yK�!b4SE����B~i%�2~�/�ז�E�%���y5t?��rǵ��Z�<�eO�u��8��5aƨ�3���܂P��5H���k��83^��#�ҏݸ�5	+J�����V���(S8��}n����l5��+L��pJ��bMc餳x���Ss����iZ�P1X{��Z����b.����6^����U����W_T�.��ul&�ĘYFk:�y����G��$=:"��:H��|	�o ��KK 5�{2�X�-0882��N��R���"�v3b�M2��c�h����k�b7U�R�]D,t��YS�GjTQ��mya��m���rsK%TgzG9�>#�r*S�0d�?O
X밽@_�Yujh����m�Z~�Q�@y7���/J�C���T:�vt"Q��*!�)qO,E�`���>��'��U|�,Ͳ@Z,���J�cG�����Y��>N���137F@`&���V޷c__��T �{"���H�O)�L���Y��m�`!�_�2��?�h��;0\��@���s�"��I�=<����/}�m,�	�����2���.�-��T�cګ��CJB���p�m�$����
�X�F>�>����J��S����ܰ��ϳ�4�JC��f�ָ�7�{#S��>1E�.�����i��nA�kL�Nz�;͢���fM�J��20���p~`��i�͐ċ\q_�Z6��r�y��.ZA��A���m�5&����h`�j'���>�����G�F����:�0�P��LP�o�|�> #�|�2�ԕ�V
#É<����W�4^2f�JJ�pތ�6&-�[�����`h;t@MU0B����~	�z\������2P�i��xZ�&���Gˢ��yT�O#����.e6a��}LL����
�^e"�KdB�6Wv��3^3��{@�8wB��?�(�	6i`�x4o4�\L���PlQ���F����2,5"���*�O9R�U�9��Gy1��M��>cn<�v�/�Z��ZҸZ�~;�>����B����AN��P�O�� �
f�4�(�|��2	���"���g{A�\��S�E�F��-(�~���:�%0ҁ��v
) b�=�2��@�����C�_�v{�}7�zD}�(�.Ŧ��>&�� ���s�vϚf/��B��E�4�XV�i�����_#��\t�u���̥��f߀w�����
���R�_�P��Uڳ��AR� G��~���u	
����K�f6��h�v��,��F�Z��C�.�q�#Ƞlf՞j�-�A������2��=�y�#��,F�xeefzν�-���G�@�F<V��N��__��#a�:���N�Z`�|]��f�f�����
Ե��LD+��B-y�Zz�����Z,�k����<�x��P���R���8�ԡU;j�Ю�.�4��*��=�T���W��"&�\[d�P���>��q�FD�?<���0��2�c�t=�7g���C]�����,P�2P(��*F(���ykɈ�u�l�6���K`A�Rs9/� _��"$<P)2����I�`IS
Ue�w���{���:
H�L0f?T9��j�n�(��, �-�E���Q�h`z2P�_-�v 3 8�>��� }�^��D	Ǝ�l-�g�!��={��̩l��|��⺶�$�9��|)�;PB�< �c]�:D��&E���)���8[}p�[�	Nw�~�σd ��Pr�[��CiVDf�]�����
%�R��7����ź5κ��@��m^+�HO�)A=��o�E����\zeS��ݩ�D��_b&���t�t[�	�Al؆?����P���x�D�
ѿu<��P�|{t�z������Ԅ���v��Yi�W�y��7��e��̀=.�o��W�47fko��|�l��1}3�u��yK�^rì�W������v�����I)Ő�ITp�bR�CjC���j����[�{��ʎs����`�
�b}<J��P���-�N>���]y�@�;��g���6�E�t���@�NRl���˝Rq6,m��*�ݧB��݄X3wP��S|����L`��8,/X:m����֤���6�.��fc���
p�����2�?����L�E���P�&��Yt	fu[r��La1q�\NO�+H4|z��8=4j��er���Ǌa���p7H�A�H,�j����Qk*�:�\$1Q�|����Z1k%�M����~�������P=4L�`'��URcw�g��U�d�Ɲ�s9:u�HH%���y#^�� ���Y��F�$A��a�Tc�և�N	j��%�ٝ��>��9�ʾ�,Rk?�z����4*���蘻��Z���l?�u�5��� a����6����7&�k�?��5���Ԕ1,�[�����p�����Ȍ�|��[�z�q��_�"�C�W��E�������DȚ|�JM��p��d����vZiAN���c@C��!�p�UnK��R��M�I������Փ�d�w�b�z,;̼uLͯ�K�ǉ��˕���pL#0r�8�%
TJ�k��Ъ�N��{��'�c*��w���F����� ��>o^C�Б�U���+�<�j:��HR�f����G��c��s��L�p^�!Hѻ�J����$!���h̨ۍ>&���������[OX�#)F�\���V�j6�CBi��_�#P7�9���*��
l���_��I;�y�e��H�vK ^��"��G�;q_N��#~�=1̖���X���ˁ'�d��4�����9��"�A�}�]�\�s�B�O+���D�<7����w/b�w 
 ���z�����r/�I�@�XUf�֙܉ny��0a�r�n9��_��&�P�o�d����F�O
$5�n�ĸH�j��g���1�7@��O>:kQ��k*!Џр�C����!s�j0�类���FX�q{ckv���:��a�C�<!ؾ]S�A����.o�R�޲J>��Z���'y��>��""��-�4B0��4�]�����~�V9�i��?G�����S`?���Nv~D(%�m�S��	���ɀ
�}�tZ={rB�l�5v9̠�ῡ����kꐄ̨G���d��ˬ�5#OjѦV��G4�^�h��-ޒ��Oh+eMG�'(V���cҳ�zxhn�3�Ǯ�تyL��J:��b(̤�ȗ�i�s�A�/_���X��TZ�hn�S�Lm¸��6Y�"�$%��xu�r-_���.��Xla���3�Ffբy�ҕ$:b":)3:#��|D��o��KF�ޚ�W�XC��0S 2s�����Ё��ݐ�s�~s�#�hR�Mۆw�7��-\Dg5f��;gBf�Qm7�m4H���W��A�*&��T�F�G�#�#z�Qr��n0����
ӷ#��oY�A^h���h<~*#�@44E����7[�����u�ct�z�%~�)�K�En�f���(�Q���0.^,����&���J<�9_�������:씕~|1n/�@�%����GV9
t�n�ȩ#������u�,�L����3`A��d�z�ڪi���CJ�v>+�h���a"������丹H����m鉶	4�~|9A���.Po���c�����#Ȏ]��̨�o$g�����١>������K���wǚ^���빂�N ��E-����0��b֐�ݒ"��E\{��
J�Spn<_o���	Z�;*�x��L�f(���w��G�B~����K/{\�!�Z��r�.δi��� ���4�Ґ�Z�D�>h{�Jj�k��<��&�ȕ
�F��ޕ��kg�of>�- |����0�Vى��Υ�c�4!�h2�J�&��}Ȯ[����goh�
�@h�vB*���Yj����ݠ.�}��ƶ�6�x��&�GF��T2�s�!).��a�O}�8�"=
&k"�B
d}J�W�*3Y(v�F< @�p�]�����䗗i���xϳ��W�ݎ�]�P'ɸ����.�|�',pʯ�r�%a�9��Uq���b~+�X�$��<*;/buu�DZ-�hrW�Y�4�Q6B�w	^A�[Px���0+f:��(AඛM�g�>]ƣ
��
�\���@�!D0-�*��d����\G���S����8�32���;W��^���O|}W�\=()�ͦ�E>�\ c��s��f��3��Q��0=4$��dzH���,]ｔ��`����_"�V ������V
� �kc;��|!U�&�|R� ��~��N�c_،��K�K�i�v���Y�I5w���	��D����\l��jHy������'���8Dd��Ѡ��x���zIT-`�ɂ�0آ�0V���&;���K	#|��N�k팷�$�M�f�m�8�h[]DF��B��1ZU�����0��J#k�̃�n�x�ܹP��/Ro�X桐}��k8�.{��ƅzƈ�v��^�W-`6&�n�d�^�nw> %�q�����\��%T2� tx��gn[�CX�$�'��P�0!( �*�d/���y���<@
g�۞칔`:���m//E���5<��Ҕ��_D��I�ge��@��7���
#�L>�B?��l�:�j>��(��� �6�̈́����QĜ[`>��Z��v[��8�h���e�J��X��l�7���_!uw0=6�6�ĸ���|�u�$�_x^/�PB]lA ����#qG�XA��[ul)�C�8���V��NҘ3�^ �Bߌ� ��o�~4D���㮟�C�j�?���D!�w�Ӻ�~��������Cť�vCؠ�;�`���0Xe.g"pf�{�Z��&Qha�/[�෼�����"=B��?����Gw|�BEz�@w����Կ�Jǡ�v��0I�XT��i���Ɗ�=	�#�M�����ff��ח���>�3�#��r}^M���ϵ��v�8g��U#�K8�T�JR�G�j������B ={�+���>����`�b����Ǳ����ȱQ>z��f�~��W�V`�g4��6�]
t(����XN ���*O��+,��*'1�B��΄�Qw댽SwMf�(`�U?8Gjd:�^k��D���,��e���G��v{pmd�Y�?|���44L�yD�4&�>IY�Fu�4 ���Ǖ�L�=\�]lO��+C.gzo�18�������D��6�a3�pҟa�E��VBH�������5����$l��|�ͤ��+�1ƴ�M�p�ܙ���n����4�^�'U8�f�R�18"����!��$9u�UH�����_^C�� ijƓt�h�#�w�h?[��LT�4"ւ��	ř%��񴮮�0Uʙ�5��`��S��*4�Sb��ui��uǦHӢT �Ξq6��`��W�k9_�ǃiۖâ-�Ϧk,o������^��d[����Ҋ֕��L��䚟��ޛ۳�:Ft����И����7M�T�8D�b�vUQ���Є6:CV��3n&�ڬ����Uk���O�ڛ�N:�d��sb��nz���~�������T���^pg#sr<Q%��M�����E��N�ؙ�gE��q�jzw[�F���S{.�h?8^>ع���ɭ@*�<{�:^�AR�/����̇�w<c��²I�p �H�|bJ/�+���y�X��vd�&��.�W��&��&O�!�e�\!����.�6�-i޹�:��R3j.I:*�Ƚl��_in�;�^���=�Hk�� y(�"W���"Wq�^���:O�8<���Xjh�˜~�'Su��~(�4�㪌��A���A7']<� �M����he|D"��7R����b?8� ����h��+��M�I r�X�֔H�nԴx0���g���{�� �ի�d�/�A/�f �5FP��a���G4�B��XeCf���Q`:ƒO�&��Ъ�xҾ6���!�*�09���[(F�4n�v�{~ZR�j͔���亠<��������Xt6� �ͷ��%�����;���ա�U�<А;c�O���]�E��C ��1цd��4���s�S{�~K;��Z.e	4���.��"��q��tu�4r��Y�D���q�<���Y���r�qU���=�F�t5���������O�^�����L�a��+��ч�� V�����q���n����"H,��o�L�jJ�p�bឤ)���E[_s�A�c�|�gX��Z�ژI6���"��C|p6T�	�z�3P6�_�_Jtx.]ll�}v�Ί�Fa�yq�R��v�$7WR"��&:�y>|e�oVIKAd�1��X��0n(�2��^�(�5_��N}�ϰ�~$h`#ۡjd7���*�D����D=�XQ��=m�N���5�����T�2
Go�%#u��r࿩0�gk3�
N���6Y�8�h_��c�~��@�P���w����޺���DtX�� ��)'h E)�$������� �,C��^���S�J��K�O��M�⵹��Y�S1�G�@�E�����V�|ٺ���qʶu����O�L)������tk���(k���Y���ln�����)"VmC��:�ԓͺ%��m�	o#��g����.�����5(c��9z�8͢���$v�� ���*������m���,�9���&	K��6��@7��(k�U�Y��ϒ�=,E7���<d���pn74�z��Y6;E�֗	'�f��	ݖ��׬~���s�����\�KZ,$5r\���"x����l�����"h�}�j�Z�h�����0��F�>p��t��ƾz���o�Ӓ>�X�|7���_�V �� �`�-4<��2\��J���*9icge[�v	��]h��R@�Q�B�-	�4���tx��l�@y���x����Ɵ�G����<'Tm~�����.	�ay3�}�ńن
��"��d��UW���3TU5���@k��x/#5�Ϳ1i�tKxj��R��VU�P�D�1��v��T ,�����Aa $9�<U,���}���Ӿ+����<N�/������Z�3�-PG�t�k��I[�R��A�9�P{���Gf�s(�cM�h�������~8���\����;���-��z�*r��c�7 ��2V9b�3��2wv������yi�lDn}���[~(��.����>�UN ��s�i�ϐţ�q��>:�4��\�_�q�=��\�ߊՒk���9]�~߶���
�
ni���BĠ����R�U����ri }�|~�͠+���GO
K*A)���Hvl�>�����	��������hݙI}l��j�������?]��3�J�l������x���z�
�-;l�ɽ��=�<V��e�6Q�y��#�
����No�*������<f�VT��7��#M2Da�`B#�	Z0����AN����k��S�s��x�Y�P���R|������ڰ�.v�!������~��^sW�B�&z��dX[��	 �>��DqJu���A.�&�R�2���t�[�g	�~CS_Q��RbPnN6(�u:*<�ݨ�3y�e���*b1]�G�=`�Knӈ�/�g���hP<�%�28?�FI	;�eO�������
���LyB�?�����j��A(`T
 
:�'�k�Q�@`�iP�UK�v�8?������֧��<�Zlc���FB!� `=�][��$��rl��pTB$G�`��PB�@F Z��>����{��6�))%	a8�6g�Q��N-��I�����;{�ʤ���ED�z=��yf���
��Y��qu��U���m���Y��i�>[��˩�[�l�{�E��sve	�SVOz)�U�&����[/��7��H��?Z��֞:+�u�c�L^�|�0�zz�p�n�����v�<]"��'e�/�e�^���p����=䀨و���jڌfaӱ�2�&�Lks3�ݵ�o�h^(e����%u�v��O�T����T��GR
��j�t&��n���{����D�w��`$bs�!�C,��߫�c�>u�2��AĘ�%�q�_g��S6c��tc�+�v��N
܁;�2���,�d
*���B��/�Ώ�w���Sr,��ݑ`�9W8b�x:c��C�L��d�C�NH�Xz�p(q���?��#�m}Lδ���&~�Y*F�u�.��	QB��'��\ļ�O7^K+>H�z�X\8�q�-�[�.Ť��aZ��pmQ�*r����H�妻ҢXG d��1�$��|0����۱1!d�Mdܴ����B�����4��a'�r��R��:��#���Z�G���9�kH~�����w^��� $�����Cz��TnT��&�}�r	 ʙ%>1ʴ�a���F+�ts�ȍ��O���h^*p��)����k�b�Yu�7kO� �9؞i6Mt����kT���͖��T�
^z,
y �	F��&��8`��DL�Q�^�'�j��a6�y�׳�w��z�H����ښr�M���s�����vPY�݂�?)XC!Z2�f�tn��Ȃ��5E���e�5���	�}d�b��z�ꋼ��JY����x�5fr���Hp�C�r�_�%�Y������Y?N�A����v��1��u�w�W�Fl[ۄ�t��`^9��L�u��H <8q:�CfR�i�	��#�c��M����p���H^~J�����(�WgN�[ &�h����|�{[���ӲONqߣw\\������6�M�ik����m�"��	*p��l/�_;�;��Y��vH&�� �ʋ"��~���,qՎ��Jr��3gp�X��X%>&˷�'Υ�Yhu42��_j��/A��]��R�ŗ�&CP�D]=7혲���b�} �ש�(!��|�(;�I[��X�7�֏Լn/��0�qC�����U�T��@��d�c��<��V�5RF����`�2����yl޴��s�:!����#Z�����9�q�[��!��0�B���H:F�����{�i���z�gŷ��:<W6����8��T#��;�H�6� �O�У���&���$��Ǘ�Ki�j졪y%Y]��R�~��%,A�_\��A6�R,xS��R�}ա~������| oV�����6[2�,�tt���r8�R��1��ÿ׆���c�F+���?h�����_v5�`����}�3^Ӧ.���=��r+�O��f%V�2���0'찥Gn���}L�NT�L��J0p�b��a�dw��l�s,���h�7?	X�kZ%U$�Ω�������6O����#_��J���;_�	�.8K�l�]"�ir�F\k0y���x�e$R�
"0��:�i�|�P�o�p�K<�Ś�aX��
0�P�2i��vÿ�pU��G�@�ٴlh��|ۼ}�7uX�oD���*m�8�Q#�qm�u���3��7Wܗ#T?G
+�#p��r;��0C�N�`
ɰ���xY&P�h�]��^�n~�%�@����K�-�ޕ8i��t�-���r)���E�W��3]��G�����,~ړ+3����aJ�9~�#�����0�&�4��1��@1���։V����Z������VжP=�� �QL�L����&;����_j���j�%�S!���n�"�U��n����庠�m���	�|������.����+c+Nw��6X�D��P$�a���@��Wi~�o�B�5�~� ޚ���ax�τ���;a�w���l���G)���E��w���:��n2)�%�)�y�;`����!Jf�Zs�Dbh�}�~�?	��G��d�\�xZ�ir7���ߪB��m��*�F�����Jh�j�j�lg�*�M=b���Fޔ��K�����x�o\��>��|r�2�f��V�%��M���G4WG(2�ݺJb�P�e���?�[�b:��khl�n@��{B �u����+1Ǡd_���g�zC�x�^C��8�G<x��6T�E��WT�.��a���}}���
0
�"�Xd���WG�"3O�p���i@&@2�����͚��iR)x�8�M�Վ�l�P����.�_$H�n�/,�z��P1��9c�U�B��w�N�����<��D/�
����Z㠥�h���ߊ�G}`�-/EA�7�P�@�`f�(�h��>���Y��,��\Q�R�62,���-Y�n�Ex0��,��)'����W�.�I2�da�ȔZG��X�}�~�z�(_����m>7oc �Ks�E��%��L�i�yd-4ZM�Z��8��n���QҒ�<��]3���J(�Q���z�
��'ȃ�����z��GIUkBG��& �~���x��5�KE�ΧʡvG���HLk������?�t�T�l�j>pi�����z����+�.�-�ǔˠ]��x�^�z?�"-T��w���aV�&��Q��49~#�h�^NJ��-B����f��w��}D��^�D|CB�^.Z�4�0�?�+�k����0gx?��P��R��lɅ١b���.q���;�e�n���&}�W#E&U�/d�跼�T�>��Sq�<��p��I��X2n��t���g�z�CN�9��D]P)��(�j�*�u�݃5�y	��r5�]�����F`��ӣ��/;K �g�<�o�ͭ�:�Id�e
s�}��u̓
ٴGL���?%{��j�hX(3� %����F�PQ:_`K�$�P
Ev� 8���(��[L�ւ�w��l��6�Ѐ!+�o=�Rd������{��KS}$�h������
B5K �;�Y?��N�'���)`��8,�F�LԨN���LT.����߂��������ًD7rA��d����VKC�߾��mFS��m��W�=�>&��9i:Ap����~�&��e䜁�\���P�E&�0�U�[J����T�О��z$x��5he��w����|�>ez�Ö�I���5�V�� ��>��h%J� ~�ۛb��/=�,������f\�����S��D3�����!�^h��`���v�r�������T��R��ij�vլ���x��{���ʟy��2Y�`(�ab�����(���0�>p���I�q ���g*��6>�t�@����Nށ��v��{B,��v*8�Bg� �	�w!��Sm���Վ`L=�8}@�:���팀k�G�Ҙ�f��d���=p��j�8�?rϗ��vL<B٤j�;&y�1Y��FuMH�Z��^S��\�;�O��!+9�Qz%�f8n���i]�P��t�a�'Ip#S�/A�R�H]K��ɂ�*��ˋ$�X|�&����G1|3M�O�ϒ-�d�i���4�~0'�g|�Rt����>�b��@:�zdW9�;H����Kl^� 0 �뭓�p@��E�����$dT4#�x��	{�%��&��4ݲ}�Oy�O`�K8?��d*�
�����b���c�u}�=I� 2����6���h�ko���y�
�y:L�E5],�7>��~��.��4��-�̤r���D���K��Լ*w<�U� b0��Q�M��U����Rk�vK�5_ ��;�C<Ķ��n�n�S9�{�5׆��7�� ���U�d&�b��z���&�ۯ��/��cڐ��E�p���r�[%����=�{/�N����v^����XwQ�cFG�ńɍܞ�^4`���o�����<S��:T�R�!ՔD�򇾮'c�����p���H"_�J%����z���ͨ�qe&�R�����6�<��O����X\��']6�yi�fn��b2��c$�e*K�Slj�D_�'�;�>��v!H�V� ���"Mξ�ؠmq�����.�ܖ�Q�X�3��Ҹ�'I�Z�4Ȟ4mz��!k�IA�>]�~	��]���s[&D�jk7�ƭ��]b�� ;���C���|���[I�4�X&��֊� n��J0�"��#8�о3η��K�.dQg9�7����5�sA�	�T�� }���[� Hy#뷵�:|u�������=�Ҵ�B�6el!$/�0oۮ�U�FimL�4{����`��B'l�0�z<�z���R,�����Vؚ�Re��J�L�q�b��Ǵ�2��������^]q���f��F��Z�;Po��WS����ș~���?��p��3	ɑ���H�t�n�r��W��?��Q��rw#�爉ꡮ��x.�2W?�<�5���Ws���^�u��>�3��\+� ���:�Vp�B��Kl;n��"���K�	Y�L�nJ���b����a*�{�Ks���@�m��ήX��Z�����$��쬸y�/6J��5Sd��eh�#J_@��.�"l^�z�FWfy':�3�q$m�"��r:�y|�[Oo��K7x��WXt0�0��R2�X�Q~߁�kƐ��x���4eTh��Z�װ�7��S�նD9�ŵ�3�Q~iEme����Q��8Z���TSk�G���#k�r��_0���i��
D�D����Ya�^hS|�Y�-~;W@e�b��?��a4�p��&9�t����U�)� E�?��N<��q���S,�'-�'���C�JM����r�5��⫴q�S}1�@��޾�)EVJ�$O�6�i��g���+���;�L_����D���Æ��HD��W��"s')Q��VK��W�"^=�)�r�
��wQmzcU	���M�����.a;�@S�cF��/pb��~��Y�$8m����ٲǾ�*ᎄPP���ۚܜX�.�6������� ��뒓��E�W��x&�՗�n->��]��:�~;{�*��;f��K�N�QI~��)'f�|/"\�'MZ"�{r0�[��X�냊�[ҡ���u/�h�w�j@h����(�f-F�
Yަ���<`��pgoתL>��|��2�[�V�f��NE��F�4r*�2R$�J=B�����8i[�n��xTZh'�.@��:B�0��L��fʠ����Β���&xF����PG�Tfg�T�,^��"^.-�a/��}8����
�<"p'�d.�EW���3J(�W@��x�-�+��u}�iLOx�Aj�H!<���PX���I��ѯ�I�,!����@�
�9�U]U�0��M��ɯ����<��/3���NEZ>.�����/����Q��`A:VvPI&&��tfKVB(r���B����T�4��g&y\�L��1�[Ue�-3�`�Һ���1�b����)�.2-s��l�ȯk��b�6}�B�0�|(����ӣ>��X �f�s�A�φ�Ȟ'>�ܴ��4��C�Ui9��;�^��9W�aȪ8M����쩏��
|
$h��>���y�
]_UF �- ���~�cy�2�ؽ:`K`�<��*�v"���
�K���������K�lҵj�����ĵ)n�Ui�)��"����&x��?z�׷-�ׇ�3�y�s(�V����7�ð�߮#��_��SN%^��h����~f�DיI䔵��(D��B�Z槶�kP��f�k�b�)��x���P�klRr�s�L��A�<��.l�=ƖO5�)�X�A�KW�g�&0d�dΕ�?��>�|�q $��+��d����2I�t)�Ug?:�CI�ޒ8W�P��,(�*2.�^��yW̿�`�X����`k�+Ӿ��/�N��B.=<<�l�hC;5\I��eņR�8h���
��<L��P?�{@�GjO�(�1x @Ƹ�9K�!��Qu�n`� 1�K��vll�8��=�Ce��0��]T���Jl�[��z!��_=ggQ�]c�h�X�&r�$�b0I��OABnIP �"��tց��P6��r�)��z8�o��GN����h0���4��n��/�D҉���o(�Tsq��+v��Vź������u�٨�4��֖��T���H���
#e�gYɂ}���K&�&bIX�`!�[eV�-F���DĵUPf��0Ի�+c���n|�l1zp��$�9�p��r�!��uQ��;e��_���������=��!��.X�CfW�/���`��$�3��e��^��ݜCf#�[��v�?��
;�|�PTܷMR _�j����VZ����{����������`C�GbiǷ}���<�4����>k_��w��,!~�Og�g�6e�tٳ�̬�N J����>d,٤�*���BB�A�Dl�w��Shث�9�`a8�۹:Y�n�gN#��>���������p����S�O?�8\? Lwֱ��&&t��Y�gu�>���8��ݳ\:�OmKP+4�Pz�kQ8)���SQ0F�ZC�a�� p� �T���CQHe�5=U��~$f�|f���y1�"�Mڠ����V����#48?3'&/p7mR� �S��Y
��P��U4�9&�H�/���<^Tf �ܷ��x����OJ���Tϭ�s�	֊>%���'Ͳ����*��>0>��@����*&���,��@��X�uX���� � ��
ƾ6���#��k�ZR��Δ�T�Ԁ,,@Ԯ�����Ҷ��Q���w�G��ݾ��KFׯ8��Q2��a����;�h�GMcj������\vF�i�K�еn CWN�\<Dn�а�>�T�T!���Ź�M��dA��b�z���a���N���A���Ϙ JIp��r��%v���W��%oN�s��x>ƨO�,��w̔HF"7@����9$^/��c��q�P<n�R:�4R[J�A��Yz�c���Z�pJ}�H=��J�3�������� �G�"&�\�?Qg��$���ODp���(\�_´³H6���i!�ȅkb���,�xM*&�6l�V�_:4;�ު�ѻ�H��� �n�"��ճu�qKO���A�)��X�I��텞'�ff�H4����SD:>AH��]m$����v}���#D��7#����bP9� �h�^G���ަ���WI��GX��%օL`n�6�0M���ڱ�K?Β"� Td��2��w#e5w� �$m��V�����	������:���W�#�����/��<F!_�0
����F�9]~{������0�kx�<�����|��#3����qVK�>�?��1t�Ft����Ɗ7f���$U��4�o�0]Lm��9[���UXc������S̿��s�}~�s�Y�v6�����p��+W��3t�i�r.Ni��m�̌����c�����Q&�3=z�M=�����5��ђg�bL^�db��W鸒��+��!�/SVK��O���R�n~[�3�+��}�L#?2J&�b����k3��us+�r��~XX��Zr�c��8θRs6E@gΐ���d�7޵ _��.�4�lM~ğ� FR��y��S��g�$�n�"&��:��b|0�1o'v7K2^�B-�X/��0� �2_�a�,Yo��Q�}�jɂQ��5�h>����$7k���[�DSz*�`�.��Q�d�m #���f�-:���CT��8G@�$#f�r���0�ܾ���
�)轇j�Y��h���T�H~���@ g��T�#�-�K&�a��t)a��24)8}�EZGv�i;$�=T5�5,���a<���@J�hCK):�P���&�h��/Z1ZP�@gdf�蜼V���
�V�4>��'A�-K�vy:L�������P�lZ����Uѷ¯U�b��������`i"g�z���T�%5/����mUAU	 ���{k���d.��3��caZֿ�ɘ���̔�$Әq��^�F���*��k�i�uI%����׶�Ϻ��1�-�Z���<� ��OE�6��2X�p�Cn(s@�1���);�@!�zv@f�N4���G���{~�m��&��7�\�i�Z�T�r�A�U+H��"���m����0�gh礖j���C�W���C�U�FԠ��Ơ�`ӈ#oRƋ>g��|�q�Ԝ�V��	�����4�-2͊�J>Ì۬�4Q[�����h⥒@Ի!B����-��	���F�����0�lx����eG2QB��T4��� .��a���}���*s�
��"K^fdiӫW}I�3E�[��-�@�����o�!��P_^i�l!x;4�Cy>�g�GP��d�����$�,\�{��p+-9�MU]�������D���:^<�6�/�[�<�Z��b^�G�ş��=D/����Au�~P�+6�T�f�.j(-�)���4�	x�����o�\��u�,��h_-ϡC�{䜺����ja�o'l��$P2��7�'~��ʜ����}~&~k:(�Ob���5>�. O�gs^:�D}��
���4���PN��N!�InQ�0@d���u��n�B�߇ư����
������kZ���!U!�(�h�= N	�~���<6�x`qK{xr���v���E?�����|ak�������6l�}�j4��f'���ʷ����$���}�Š�0
x줊z5�X-̽K�n�����V�����l����#��	EuN ���z��(tf��r��j��T�ID�5kB��[Z������aUk��캄slx���P	�PR��3��|�*�מh.g%��+��U$�\�W��&��d	ca���>�Eq[+ˍ�'���2$T�td��g��CDx?���P�g(.�*�F�9��y��O���*S�	�Xoy`&!���/1r����<w�ݔ��0łIt�e���Ss^�k��
��L*�}?[��J�j��e(�P� [��u�:��jnQ��2`��u�F�v�J�8pO��^FNQ5�8�횀l4R��{D!��/="�"�0)[���I���$�|��$����B�}U ��؏���D�Ѝ�\�)�&8b<ζBtN>VH��̃�
;�x���[��j�Dm�q�Ϛ#���k����"�c��|ͮ��(�tK�/ݜ��،�X������[e�R���K� �F�&�) �[��5��䆆�J��)�ޘ�+`.цn��}b�|�%z��f���yԫi3��u���!�r@��a؈���[v=u��9���;f"fR���C]N�}��3�ޏ�P�^�u�~����Apv�,�e��7לT��R{Q?j��c���X���H{�KZ�UȈ��~+`^��b�X�z�w��40�>f���҈��N@�4g ��6��tG	�G�lN��v�L�����,�t*��B��
�wWc"Sc�e��&	`¤�8���:�3�B<k���ɘ5�����iD�pY}�n1'?h�7�yL��>��:J&o:Y;�Gu��0�\1������\u�.O��+/V�z�$8�k*B��/t�52�a��p>&%S�(H�ԟ�#xo��U恟�$X;L| ��G122M��O�(�Z���Zh�4sj'���R*[dly�tG���ო0$�9a�pHO�o��w�^��R U�%�࠸��þ��$��KTjk�n�	1Q%o�k�;Ų
J����y1���i��޼�*�a��?=���>d���eu3���` h�G���6^�w��^�k�C�o�j�/R�ԻC�,�®�[~�7��P��7a)��3ߢ� �hz�J�����#�φ�yw�V�s��veM>\��$���qvA1:���p��Cr����)�n�mX�y��T�#����F%��:�d\!�b���zsb���\������?�F>���_p�c�r��%QҼ��?Nб:�N�<���&��
��GWWwGc9F��J�? /�ԁM^*hw�]v9�,e_<�1:J0�R6�������e�c�GW��D%p�WHX��J�T�k���UH���7&ц����,���=�#��O� p �\ږ�]u�6�̴i|o#�&����}s�*0*l���_�`�;��=�,{�HW�/ �p["C9CՎjq��c����$��iYXV��s8'?�=����4㐨���z�A���](�������X��АD�$7�����b�yt �Z��y
s�rN����IwRX\a�ր8�n@��0�ˣ�_�Ɓv�m�+��-d��#�-Kҹ�52��?���y�ڮ Do{�`�뭙�:2ؙ��^�&jҪ�(��2!��0�/����XF&��{�V�VWu��J�U8<(d}�锣�;�D�I���f��mƲ�~���秕���mv�.)�|�ب�[)��~�]'es�/-��ۡ�Pg*���AS��8��N~�����!�_�����G�)�]pYt�lr�̆�|�����k�������)�WM��ky�hC�2\�5j����{8�N�,^�sV��E_�M��+��̇�C\V&�ɔ�.��Y+ny5�����`L>^J�.�bo\K��0��as���#x�hNXu
Z����] �s7��.O6@����ϐ�*�g__6�C.�ٙl��^�:�pFM�y�Nԕ�MU$��"�+�:j�|k�go�(7K-d���dX��0ڈe2�O��To�!�P�U�S��%�h����w�7�{�t�D��͜���)2�Q4��m۩t�����[Vm*\T�#[Gۥ�#a� rL0t�b��
:�׽bf�Y�U�h���O��~��@���*�+����&���Rt�*��/O)�
EoDԄZ�ҸV,�w��,/"��p�����J0��%�k��/��,g1��C@���/�V �0��O3��]��������L����Jf��W5��齪д���e�$"f���!"��7��R��@ `���m0?�	[H��\���.���c|¿%C����H��p�$n�0����h����s��1˂����%W����UQ;�,������A�P������3E�5��(~��$n#�E6&9Ȱ��;�����Ѝfo�,���U�NJF~�?���E���$F\��Z�rrȖ��������;�W���:\h�j	�U���βȜ��F�V��\�7�������o��>BD||#x��7֗V�H�^oj�L~�4�P�2H�J�Ԍ��ω�[��u�.�h�ܚ@��0B�����.��%�5�U�ܜ���rx�CE�2��G�m,ETY[t�( :.���a���}�8�EW)
���"&��d�WÛ3@I�zY@Wg䫙!�H�+a8i©;x���>�܎�r�P�v��Ya�����G�,��0�!��p;9tz~U�D��w�� @�`�~<:��/i���JZ��Qs��/Y�������A���PQ>�-�f'(�Л����V6��/���5\"N+�'���-�0$��J��IңÅ���g����2��B��*����XV/}Y*����(0�#��'$>H{� 
��s1�3�|���{C�*�<4+b�KS����� �Kg��W�������}���"j����
��ȴm>��}F� �U��a�3� �b~�yB���3��K�up�|Kvv��$���F<�^�wǪ�P��݅��lf�j���A���+v���Dߓ����%����qxx�z�$-�ßɩ[�ة�_V~����c��e��#Cc���N۟ ��F��T|�f��J��v�T/D���BddZ�?+������}k�f-��D�xp�1P$t�Rh��Z:O���-�r��.b�J�L(Ո����w�DW��&槕dDPԼu��>�(q�R���t�i�wH�2��mt�|�gu"C?k\����PZ4(I
�*(�I��^yͲ3�C�Ni����`�.z���/��.��s�<����P+N�IuCe;Ν�n�<��Z
jn�Le�>?���۞j�\(L�v v҂��V��sQ��`X��A�v"I�8+��yG�Y���M(ʊl�h�v.e!<�=����K��^j����$3�*�V�~�"B$�Z F�>تdQڿ����f�)^�8�(v�=��N�՝}4҃���󐞮6�U�j�D������
��̘�0f�����W-�����*� Ka�G6��X���!�eu]Y?/|��A�T&*(���[�<_�#�=�a`��+�Iw��&���3�8��|)Bzf���^j���/Ǩ���C.�y�۰Q�ވ,G�w؋=P���tQ���YfM����8^38.�[O^�,��j����v�9˩�s���T�sR�c|je<C��t$�I�{�#�ʰ���cA�`y�b_b�3���������*>a��-�[���F�9�g���6ϴetO���❟N���͂����,e-*��cB�]���w��'S^*��~�`}�8�q:OW�JC��������}�c���pl���&?����L�^�;��&j	�Y�?�u~U��.|"�[�\�y�O���+*�cz6��8�p0+�xGO�A�aF�Lp�W�����c,�H�dP�>�13
i�\Yo$�0�|�����۱1�a�MP�� ����X\�5�!4��'\N�	R����菤��F�ڝ49�؉H�����=r^
Q� ������+徯�o�@�TI��i�	���%*`T�5nŲ�����J��R���U��*�<K���<��\�N�lu���?� H2� �6�����0k�L����
��z�,v3��M��g��@�RUC�=�7��lg������y����;,��4_��q�a�^9Mn��_T0�#�v<��p:��+49C��4�R7�nm*0��#���݆���׮���dwփb�P�zN�̼׿߯�ì��]<ڡ��v;�p�\rv-V%,���ͭ�LpN�%��./���Ub��w�Q6Fؒ�z�!�o"�^%푸�e��<��7:�i�R�9��)�q-c��Ҳ�p���Hs"�J��F���C�C�}u�&��ݾ�CҀgn��>D�O:��Kߙ\Ht_��V�6��i�#~���9�W���*ܙ-l�Z_p�;�~l��Z�HW�  ��"����iPq��W���.�S���X�j�#��'����ŧ�4L���)~u�A��2]�����"�lT	�;nDI]�7Yp�ib�q l�6���I��K����IGH�X�Y��{Dtn�-70Ì��.=�A��H����d"2m�("�-p5���Z�#�LV%ډy
V�J/�;p:��\�͖}�1�j�%�=��I�!ե
0@iD��<[Fz2�}-{���ɋ�����R�<�����T�cr���(��**�4+��l�X����B��üpq���7`�����e�8]}�j@��Vr�K�Fa�[�>OLS@��ic
~f�;�ϱ@lE����3ɢ||�4t��Nr$k��W)�� w�C	,��T��������iE55E���
��E^����OT����+Կ�	x�V�Ŕ�m���'nt/���&��:'LY�J��bJ�ΤP�!�L�2s���Q�}�#>�X8\�Z����w����L�J+�6;@��F�4��uB:f_��$.���l����PyFHy8	��dS-$�ȼ"��:Ei|�=�o]�K(����{X���0�0�2U����n߁\nĐ�B7�D��E6h���(
w7arOO�"D�\��O�$��Q���m�P��*l��#�H�$T�1Gv�<#\�r�0/ ��i
�"�=�LY��h$�6�JH�~L�6@����E��e���׿�t_*�L�)�ՄEжԟ���3y��R��,j�q�ŀ����J^���5���%��[��I�1Р$@�Ý����V[��Oc�jH���xⶼ����sL07*����U�.��֪K�=�e/�3���������"7u�Zƥ�[똺�0m]	�!�]��z�F.r�V�q�c��տ�܉�y��
U�$	P(�����â �[���t�k򜚀�u�Mu���'ƫ'I���v����H�88���E~T��c���}n=��:��k8�;�N��pKgfJ�5�0�w����~�A�:�FͭO\.N�Z���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸���p�&�1�#l����_�)��ToڬrN�'|V�xcĔ�MS�'
�x��� J�恰 *�y��%ّ�'=�F-zӬ���	3��t(�ن��Dq]4X�$��T	3A��"<i7�lӠ�7;Dl�ᣄb� J4��@V�|`'Ñ? �� � ?a���#��7M�r}�ҿr��hd�
�!�t��1�X�r�Jt��i�_yR�O�pԫ3�L<I�
.BV�%�q�at��1)Ct�<9T�Y|����`.��|'���h�l�<!҉�<>�J��<X-����d�<YB�K�ܕ'B_�]� ��&e�^�<ᶏ�j]̩�s��A���s�"]W�<�W��?%��ᦃȯ��hs��I�<iFI�(q��@A����P[�<a4J@�Z¢��a��	V�bHd��^�<�C��L���8����x�Z-C&`�\�<�1�B�n�TC+ֿ -��k�Y�<�C'.�(
#�W�Df�is���~�<����D԰��d�ǭ8�̹SA�֟�Z�Ox�r�}��c>Y��c��;u�޴QDU�^�D�;��]"���'��Qe"�U�'� �O��5�2�� ���Y�x[|1�@Z�l"��ɨM�h:�ʂ�9x�R�+އmu�xz�0D�T!�@   �����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   �  *  ?  N  e&   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�%J�L�TM�P������PČP_`��7ju�r�d�O���<�'�?!�Ov�up��O[��S5E\�]KXl��_�&W,X��wJ�:�͇�/|�a��lP*��<@� 	�'��Ї���X(p�1/jE	��<=Ӧ�*e��O����O��d�<�����'�Z�Q֨	�δ%�"���}!2���'�.�!�ϑ�*����M��rǠᩋ{��{Ӣ�d�<�F���?����P
�m�rbj}k3�P�\.h"� 
��|$���?��`�V ��'�(�#S��'m5�E�qb<r��
�n��x��*��M/ `Fr��㔛p�ay2D^��?Y�����}���z�ŋ_V�
P��4���O��$5�)�S��p��U��EG�`	O:}�:C�	� �ؤ�s,O�c��u�K'2��Yk�ʟ\�'��T�t�mӬ-�ah�O|��H֝�_d��5!V��`r��ռco�����?y0��?1N>q(�剚m� ���'sx��`s	U"@)FOv�"��ֱw��,y��׻�h�H�S�\�I*�a�Mk��I�x�N�?���I�Ov�O��)GY�����M���D1,O�\���N��]�6o\�`���y�a�5��'��ɸ�M��i7�' �����x����*�0z#�d�5O��ħ<!�b�?U��ϟ��	}}뒊/�� P��Z�|\�%����'�j1K��l�y��6]˘�{e�N3frY�>�!
�YX�L`Q
4vO�Q2Q�(Y�~��Ǆ��'�v��S�g�I?PB����$��%���C��NB�.W��	[W�#yѤQ#fϛf|n�'\"=ͧ�ē^�P<�uչVڎ�J��(��u�k�R7��O���O.ʓ�?)���t�"O���!b^�~�@Y����>C��G�#(D�Q��	-@�yrk�
l��Y�#�)���E		��rd� �BYB��Эl��yr@�S�ڐ�u�ϯ-��0�!g� �J,9��?I����'?��p�C���4Eʲ(����0�]+4"Or=���T��vX� ϲE�H���Fz}�U�d�5i���M�g-���M{�Ȁ�2�uC�ǧ
3`<1��Ѹ7�"R����ş�ΧB����2�F+o�Ig���4���Ӏ��Q�4�w
L�8M�]K��'��3iQ�X���*��G�U�fy�b�H6�XL"��*,O���t�'^����mvWH��ЫT%��3��'�	Οȇ剢b�l�)У��0���8VB�/�\,Xff�H�ܭx���,������O�ʓuUp�hg�i�hd���'������0�c%�9{�� 
�'..�� �'6nĸi���� $^(n�#���O��K��L ����[�5�h	�4�^��{fms�o�	h��q�O���(�@	�k
.(�v�8
l��aQ4�xj��?���h��6�C�ui��G9N&�+JJ�*HL ��� ��$S�{ӊ� ��K8�������0�����Ń%=V`�',�r���4j�@����?�E�c��m��?!��蟴֧� ��Y�nQ�&�.��g�(T�`�����A�w��8�AZ�'�\XI�p�ƙx��eJ�q�5� 扁U&(Ѣ��L<���V6�,�2�C�;NP:t�C3�b�'���D�CY��,O�6M�7>`�}���[ � i�I¹T��)�ēV: ��K�I� xcc+���v̦O��Gz��O��\�P���LFʬ�E�R�(��5(9}��U�{��'"ɧ�'����'̄�Whtes��ʋs@��������83�%I�
ZlȆȓ(�X|K@���t`�W*��xPl-��B��e���:�CÊ�aZ���"i����ңv�,����˼ZI���=�����v�ć.Q/�����V�F�r�@I�i�|h�Iy�	П"|�'�L=�B.C2v�Q:�A.���'O��#vO3+�E�cM�=?.eB�'/�$��)�F٤X*�H=1zH�
�'�� *����-�2��-�
 �	�'��i�o��C�6�Jc��aҒ���*[B�'��Ë�i�6@�N�!��F7[U-��E	�"��h����4��I\:�Y�  ��R���!�ΰB䉓x��pzg�$L����/W��B�I,]��@�6��3OM�C�PC��,K5jD��M	�xxs��&l�.��$I�'��]��l�"�x97�F58*C�'0�ʈ�4�����O
�>q����Jw<5�$�
�rąȓ:P̙u�˒7��W�J���ȓ��� f�8mV<"I֥r��ȓl�r��m���9�呸g~���4���s���3�|���e�)��ťODGz��4,��~N���w&ыV�(=B���hR�T�Iݟ�&���(,ID���3�N ae��iH~T�"OHh�3�$jWc��^;J-""O��[�☏���(a\�1iC��y�,@�@cX�	W�R������@�y��W.,d�ƃT����7m��'��#?�1�쟐#�� |�<�%ID���+9�?�J>�S����;_͊Q�O���8�s��	!�d
�]zL{�@.?�FQIьs!�%U�}�A	1�$@�C�ÚD(!��%�\R��>e����Œ���T-}T�T�Էx���gS�"&�ํ��:4Z�>r�4��=���۬�b0��+ա�?A����>��#Ș>Y�9��͚(@M���l�n�<��H�>%��	���/j��89��U�<1�A�$��k0�]2tN�b2!�T�<���	!Y����`�`G��*���S8�� ��Lu9"3�F��z��r���R��G�J=����T��I}r,��>V\!!B�w{�m��G͂�y2-x4���J�>�Ji����'�y��L3Jh<(c0���5!��!���,�y���>O�B��r���~�4 i5ȅ/�y�	
�P).Ȼ�
�-*5�T.��ɫ�HO�ִP���c��Mjwok�ĕ[כ>a#��?)����S��3��� ��WJ�4�7X�NC�3hq�[���#�,\K��ި-��B�	�6��}1��4Y.�-A�(����B�	��JI��a���'(_ \y�B�$sE����gѴ?ҡ��2Q���x����WmbO[$`���iNr@����M���t�D?�d�O>˓,��,)p�	.v�@�2E#<=��D�$}�\WےoX�|���E� <F&��3 Ә\Bh �ȓ k��aP�	V��ɶ�>p�E��J&ꬢD��Kǌq�WI��:&2�5�r<G��l5E����5jG�+"�p��L�4�$�OV��� �ً��@?2�z��&e�-��7"O<H�a�a|q�0iEyH�ʢ"O��yGiX����
-8[�"O¥ ���/��lB���{*r$��'@�<�$,�<o��7i�@pn�����x?��@���$�'�P���ƌ�u6*�ps���Ͱ--D�Pj7E��iR2=!ŝ�q�l����,D��y%�$3h�@0���g`8�`�#8D�D�s�ܽ!�,�x��*Bo��c@7D�h�"�]�,�r�Seϖ*��6�/}R�5�S��=�rU�"
	*$<�A\�/��O��­�O��D<���$-�?E�(A�s��8(�̌�C���y"@��r��\�raV�7�$aK��T��y�
ԻQ��0�DB6:�b���f���yd�,X���F��,W�a�"���y�)Hw���3���!��c'�T���'�."?�"Ǐ؟԰u�ɝ8���*1�E��	2UeN�?	K>9�S����+�P�bŠ�Xv�#�+�
�!���K�.��!�^��[E��$�!�d�;}��Ҥh�/%o�a�d��:.�!��(�~��b�?9���Fh�����+m�x�)�!@�e�^]��������8��d"M��>� �07�
E�5c�?[^�`*��?q��Ӱ>�]'S�%xd��5[��P�X�<ae�Ϊ|Jl���/v`�P��Q�<��F�:i[m����D/hL�WoV�<�������AWu��$-�]8�q��d�q���Sn��4�ƨ�U���p{��	!�����(��a}�l�/�ҀI�)Y�Ȁ����y�DU��"�:ĉ
���1��A��y�,�9_90`�B����e(��y2c����:�KO�8̩U�Y-�y2��t~��+C��,.@�ZP&����
�HO���R%e�Wvt�I�5J���>7�M=�?	����S�%9B#���S���4(� JpB�I�!�V��U�ֶ�n��7JjC�	��FTbNо�Q ��ǂU�PB��`M|�Q����s����C�I1Iz |`�)�d�y1Vo7K�v��P��$�b:�n�CQ&����|�-��͘*��d0���O>˓<����Ik�.��A&�~�V��u�di� �
*X�`x�E�?<����'2^���n	<�
�7.Z�n��ȓT>D���j��O��3kV?X�2i�`�R��	ױa�XY��*-��a�c7�cn��D�t�R��)��Q�bBF��W��W*���O>���ڡ!)J��X*@�`�r/Ǡ`8!��9ª�be�*�nP�$�ǅ'�!�dӣ;!��pF�	!´k�D�44�!�0�����:�:��e�z�x2)<�S
�́��@��F%B���
E�H��c���Gx�O���'U���g��#�슐9�e���;?xB�-�z�臌B�]�����ʒ�f�"B��F�,"���4'���
>A1�C䉂z�,�˵��*��`�d�9��B�I�ws�i:��˱ulv����;j
`�'&#=��@���tA�<�6JƱY¸��FK�D��K3L����O��O�O�B�Jq �xz��Q��8r��a�'�}�Qc�+�d��Imr��*�'n�@y �g� ���%0�b �'�a�5�T�_"谙�c�= �ֱ��'��!�5�D!H��1(��7��Z�{o$�A(����;Dx��K� q���Bj�Y�����?E�,O��1�c���8�nL�i�x�Jc"O� ~���j��u@�Y3$��!9�"O�lr�đ�gnМ8��-p7�E�e"O݈rӴ_v��؃���]3�m s
O���`�2 ��<y§�bgl�)��v�'an�c��I��9���Ce�8�j�;P5��IȟЅ�	B�h���A��D�F�B@�Ԋ-SzC��'ZyfLk�a 4N5h�h�\�C�Ƀ�*�ñd��$*�D��� 7D��2��+*���'5Uc�B!O�UGy�k�/o�*`@��9'{�	���8�~�n߼�O���O
���>�f H�!w��P)Ԩ-��A�x�<�jr��9���"*��8W��G�!���\q&�jRƌ�jN�z�!͆�!�$�?F�&)�ӫ�=mF��$��<Q'!�JN��Ab�Ɗ�D0�4�+|#�jƑ��?�Sf�aC�A���B�6��|xB�.}J^:Il��'pɧ�'hT��	�ҍ5ULl�1*F� ,Rq��!hj!P�ħ7R��"��M�
�����$��l����
� P�A7+ �ȓ��][�`�<�A�*8H6��ȓ{[�l�r��Ljx�4e> ��L�=aE��I��d�o$�zC.��9���S�U0���Id�	�"|�'%�4Ȁ�� "�"�`1,�8v���B�t���>u�|P���3L�`Ȇȓ
���C�M�o bP1�C1':�ȓ:��q�-i�ȅ�Ƙb|�P���IĦߨu�<-0�,)PΡ�b�2�;�pE��-G0Fx捳�� p���!O��p�d�O@��D��T�\]1�N�`�hC��L�)#!�� oJn���&� Mb�<���ߩp�!��$;8)��
(2�x��*B(�!�$N�N5���"		$��H��I���x"�7�<e��Q@f�%V��E�!��=&@z���M�LEx�O�"�'P�I�K��)�VK��uh�m����/Q+�B䉧u����pgB�e(����KHFB�6 �X����(}$��0�cP'I�B䉕?�xe��ˈL����&E��e�B�	J�у�W��ժ%$�/g~J�'Q"=�Rwn�&�y�� �x�!B!��Y��ޯ3���D�O�O�Oy��{�OF��5�2f�5�>�
�'�2y	'��"P1��")Q�Y�'C�#�a7|��"��?j36D�	�'e�����V~�A2҆�c����'
`u���Z#+��	:QdG�S(�a�{B�>�5�����-�t����	��88qƇ d.�}������?E�,O��Jd�+;
��E��^(:쀳"O�4ڄ+J4=���b$L�qo���"O�`���
I&�aq�N�.WhCw"O ʵMI�BR��Yä�0R� ��
O��ƭ�	�`h:N�^��+S���O4}c�-/L��m��^�ȩ�M��s������?i�=���!�Ɇ1a�����t�9��@����a
�ڐ�!��F;��t�ȓN*8��dO�*��)�eE�5͇�� ���d��5C��K�8��-�㉧�(O �*AfΊ��U���7"�)���O�Is��i>Q�	şh�'k����e�K;�x	�ʍnx�
�'�q@n��G"и��M�h���A
�'�(���Mʅ4pX9q�H#m��D��'H��;v뜬*���A���.�@�z�'�*�;�ɝ|+D r"ǚ��D�L�t�������a��Q��*Lf�
ܒ�b�%e�M3���?�H>%?	�o��6.�m(�I�8Z:vy(v-)D�|(ӣ�1dP�My��ئ@�8{dF+D�� ��$C��7�^�a�-���r"O�}Ӡ�K��l�ŉT�S1��ڒ"O.�
R�Ks�� �")�
6>�����d�'�:C�dD�x$!�[�^�o�=$�@F�'�'%��Y�����ޚI�Y�$M���񃡥!D��0�m�+'>Qd��,<�h�c$!D������Y�x8pM� �F����?D���D�C�X�>j4 ɶ@��\Ї.3����-� l���"
5�lC4�M<�Q�,�W�?�'v�p20�ĺ4J��J�a_)z��`��'���''X�B�.�"r�f@���>:����'�����GJgL���#Y�-ؘ���'��u���Z+X!D�ी�V,R)
�'7�		@� �-G��"�B�S.�b	Ǔ|�Q�\���?
(�R�R�N��4�W�'&ԧ�����Ol�2�9B�H�GR@�����;��U+�+0�]8���OL�m�n�g≉"��"H\�eơ�'�P~rNP���*�;"�'����!9�3�P����@+ � YV`��|�=��|~���4�?�'�HO�p��I �LyR"�ߊ�,x0V"O���f'�ē�!ZN��y��>q��i>q��Q}B���c���;֍�
]N4P�]�Q�*�9���	�$��O$P\�`�o���pҁ�8e��)Ә%c�ى%O��|Pt� �'3����5�L��I�V�j�+�F�"	�6�"��Г)�B&�'�0M��K�3|>�#j:h�`�Y� �$�?���hO�b����W�Pnb��5�������.D����Q7h�&HkeQ"C�I�2I-��.�M������'t��O�V���Sl�I6�A6BzdL(ϙ1�T�Ĵ<���?Q�O<L2cK��&u���A�C���w��I�pE�Pn�wk�r��]q8�,�V
��^5 Vl�@�|��܊V��`�C�d�q��:k �xR`��`�	R}�i��3�`��Fg/0�(�� ��#�'a{��I_��X$f�w_H�
�Px2K�/M�����)��gv��#H˗�\����'�剞vb ,{ٴ !��K����'�u����lHі�2�P�)��Ε!H����ONAX�.��0�� ��Z5��Uϙ���tW?�k��'o��d�FÄP����'�L�� ���^�
��e	����|B���J�X�'�	�>\9��S��1<^���O8�}BشY����Į�!��=��D�q��[�d`�mԁyi�zV�F���p8�����䋸X.��@d�'�|Ƞ�I�CF����4~�v�p��?I�m�?9��ƟH�If}�!Q="�̑��G�vhݫ��80>�M"3mP�#���	)K�0b�1�3���*��Pz��RM���(X�\������F<&����X�f���xrkD��>��F)ńE���Ɓ�t�"��%?�!�Cӟ���>	� �A]���R�W�G����t,PA�<�W���D�h`�`��@��e�����'~�I�E��T�m)hi��g+��(���'/,�Z�'1��|J~��)_�!�$�pd��,�����*�X�<�%>Sx���hɰ�6T�<�aɒ;-2��׈0[�時��g�<a��ҘkyVu���]�j���Zi�<A!۶���)%��5���P"��^ܓ"���tB��O�9�(PǮ!��	�6�v�(d@�ɟ�&���)�gy2m�z\��;�f�T�t�҄��y"���P�pi� ?HL�${5<�y�N(J>�RW  <'Α��� �yR��T��Igd<b���� ��Px��*�:, l�6MGl�����r_|`E}�A��h�����A N��,r���5;���B�럀��fX�Pk�㔻��}C[BX�$�<f$!�D�o0q˃틛o`1hFkJ	!�/��8 |�@�@@U'�!�$� kr�L���Ӽ~8DБ��"Z��x��,ʓ#cD`XdT!H@ya �� �Lm�ȓ
�*� @�?D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  5  �  $  )  4  !?  J  �U  _`  �k  �u  �|  7�  �  W�  ��  �  O�  ��  �  s�  ��  g�  ��  /�  ��  ��  !�  b�  ��  ]�   W � � � d$ J- �3 U6  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9�ӄ1Z���1.*��5�����)z� B�4��E��c��q�B�s�'$Nݫ�%�a���%䀄�r=�
�'�P�1A��BC�a�M�z�l��'��yS�H_���R
\�wz`A�'R����,'3��:��^f���'V�s �^r:�r#�ԓf*%0	�'�6}�Wʈ���¢G(M�Z �I<Q
�6����hGy�؀AK&�z)�ȓj�B��m٩���2a�(
��ȅȓ�]:�L�6�ZA���f#~8�ȓ������#'*XAc��Eb*��ȓ>� q �IH�p9�U1g�Z�Y�)�ȓt$]��_��a{p�ӆ-��E��|�~�w �b���:��k��'��}�ˇA�~���W�@Ġ 遱�yB�L�	��R4�U*P�(7�[/�y�F��M$��W�NK�����y⍄c��#��ChʡE��yb( <�*((��݇py�xI�
�yr�'[�ЙS�/��Wy�U�s��
�y§_&M�y�%, �LϜ��BB��ybk	.^☽0#�/���8����y"A�2Xɛ�,�w�W2�y��Y�+.���d��<,:y�F�O��y2�˪P�$��e"ٙ3Z���U��y�'�4�����$�J�R��S�yr��dq���V�#_�m�fA-�y�L��LY��LI�1ch܋a����y�GV��ac'턖:�x�׃��yR�߫XX�di)\2��tc7����y���[2���E-a�nq�Y��y�%�y��8Dc�WӸ]6뇑�y�凖B&��)tFZ.7n�a���ލ�y�J�.n���I�߼W�Vй�b��y"��Z�,�"3�	K��� ��y��E�*�����P'H�Yw�H �y�	"u]�@�ӚQ�왒6Fݺ�y
� ���6Q�,N�L�c�1LiVฒ"O�1Ue�Ji�m�r�ZU��"OJ�#Eh3�4��I�E���Y�it�"=E�ܴ�਱�c������N�XY����?����*lYS��ɒx�l
1ITv?q�xL�Z��߃�9#q� 3�����If���|%�9:���_�r�$�wl!����r��� ���QR�"�&d!�׃���jf-Y�w�����*.�!�d��O��3Ԅ��z~@��	L��'��|2kS�p�\��g�.;��=�I�:�y@֑,\�����i����FAE��y"Ǌ�a�L�J�i׌^'A�$�ȕ�0=���Mw�xcgmz(����yB�Ļ4Z��%a��`�f:Ը'5ў����[��&4d��� ��6��!��"Or`&'_8)��� m>��ѷ�IkX�� ֋�Fئ�	���l7��5�;D�P�k7���������@�O0B�I@����JQ ^��a�ʙ&yJC�I�C��|giE� ;�m��	%r~�Y��R���1M,C��C$�Y��̅�TD���Aǘ&@��Cb�<Ԩ�ȓ(��D�G��8����Z&H%�F{��T�����HܖsT��r᎛�yR�ܺtWd��AڱZ��������yRf�8^n<YvH�4L�p�6��4�y�DJ�g��EԏC�Lx���H��yZI��Ec��E�U��@w���,C�Ɏ|U��g�/j�@��^S�C�	.@[�S%\�\�� i�B�	;>F��T�S����w 9W��B��	�<�g�$&�����(��B�,�m� 'R3p�re8�ۿWO�B�I�H�
Q��u�xI�4Z�	WbC��6� �ƥي�T]1#�"�B�J�(����1Y(]�G@��i$tB�!$�4���7c�ֹh�FO	{jZB��5
kҹa7�:&��鐒��;vC��<R�44;lK>B�<x7E�<u��B�	?�\�P-I��|h��Q+�hB䉐{�
�[�dZ�ڙ�r>�VB䉣6j����h�܅�"`B�ɴaɈ}��e@v��Er��W	f�TC�	.ac��v��9W�l�)5N��Rk|C�I�V$U��f�t&��ZV�Q�1�FC��<3^��5 9Jc
���*i >C�ɦVr~�y�&�?rr�QZ�ƒ2w�!� �v9���ٰA`@���ѢX�!�d��m��	�O�m/Ľ�0��t|!���	/{�Gj�4��AMU�F_!�d�2nl���m��!�n��5����!��݅�F�X�̂� ̌�1�D�	A!�"y��Cff@	s�~�8���*[�!�D6L�y�<q��4*�ğ�)�!�ԄXT�y�����~�ꡃe�j�!���U�M�#�K�#�V� ���d�!���PFe�Q��Vv���7tZ!�W�Z<TZ`-_�:U�u8ፌ�	O!��1��pCV�@?cS��;Э�}>!�
��)��Eގ����H��!򄜅QQ������e��x�g�R�d�!�ز\v,Y�M�9L��8�'S�\�!�8����#�7��1A�9J�!�� ��X@O��L�f<���әDL���"O�(#"��
$���k�{X�P�C"O�E�P�A0Txp��W
�Fq�m��"Oz��a��`���HG��R`x$"O���W�[�h��d���T�y0�3��'M��'��'��'�b�'s�'C����F��[P�	�}w����'a��'n"�'9��'�2�'B�'o�$yB�jd�	sPWn��s�'�"�'.��'0��'R2�'d��'��I���a�.������^v�)3��'"��'2�'�r�'�b�'|2�',���1��M2U��_%� �'g��'.��'�2�'�2�'��'X�����	Fh�S$��J�1�7�'��'i�'db�'PB�'��'٩����@H��h��]�U%�����'�R�'aB�'z2�'~��'Y�'�p�2�*ʘ9��N܅,I�}R��'��'��'r2�'��' ��'����ǯ��EQ�Aw�q����2�'���'���'r�'QR�'��@H�	�<p��	ߊ`���«�3�B�'���'���'���'vb�'����C������]�w|�lBR�J7B�'�r�'�'���'J��'=��[M�l5R��#Q�&�����u<��'���'~��'���'��'6B�МS󴸋���3P�ȭ���@��'�r�'}r�'��'�7�O�ĉ|�xtQ���}|�2w͐<&�l�'�Z�b>�5țF(ދ�,��D�7G5�q�-�7�yRY�lzߴ��'%���?�
��PA��S!J��9r�cζ�?���MߌU��4���g>i�����S�=���@�
�8m�����-��d��c����ty��=�!ӖAO
ED��� �ɐ?d��OPʓ�?���/o���Z0M��k�̢du� ¡�P�&x,�D�O��`}����)8���<O����܈xW(�y3�;�=�08O��I�?i�?��|B��g	4����4v�E��&		4�͓��$:���g��?�բD-e1�N#7�Ȑ���ҟ��'���?1���y�T�<MC$E+���hOz�b���%?��O�*8��f�'O�(��&�?��ɏVf�C�䄙����Fm�!��$�<��S��yrC�\p��8c��a�D��Ab��@'BD�>q/O1oZP�Ӽ3�YH����'&�,T,VMC���<����?��L@۴��$v>=���gj���\-IL
� �N��6�$�<�'�?I��?a��?!f� T��(�VD@l�}a�&����\]}��'.2�'��O/R#�=vr anƫ�	�r'R�]�.��?y����S�'V�R%�s��\����2X��&���M�Of`1�cڼ�~B�|r]���w��0v�҅�Ӓ"vh|��3�O���'���]3/���%�[�p�8��G� p�҉~�p㟌��Od��O6�d�,�
5+�!"�%�¾Uy�8(��q�
����92˦?�'?I��.i[\ѳ��:üI� �N�V�
�I}����f!��w� �	�Y�u>��� � ɟ���ٟ|ٮO�S��M�J>�ƄW(c8�H��1m�� KFO�����?I��|�4�Ώ�M��O��\(G:l�h�`�M�`����fuҁ�#�O�Y�N>�,O��ĸ�c�N""�'A�	JS"H�w�'Q���՟���ʟ`�OJГ�U 	<�u��nY!I�-R�O1�'���'�ɧ�) C��!˂n�<0iAG��  1f+��a��7-ty�O'�����mwz���f����Fi�^�I��?y��?1�Ş��d�Ѧ�R!��q�d�P�ǊH�zL8��o���'�.7-#�	�����O���(��X��4�&%	�}��Cs�<Qs���M��OP�;4�ϳ��wH�<� �@
``;T\Xo&@H��<�(Ob�����e�MI��7b�U�0@S�N�8�'���'������睉s�BH�
_�_���ز��Dbh����L&�b>5%ĦΓ~ު����E��1�Q���Kz( �>��Q�d���x'�|�'��I>b��T#/.� 8��3d����h}��'�R�'��h ��N���S�,¼��9����S}��'���|�'<EҒ����h�)�P	أ��čR�v�p�b�$?yp�O���><��Rde�: �2� �88����O ���O��d8ڧ�?���!U,�DJmM$thna�ˏ��?��Q����؟ 2۴���y[�D�:�Ϟ97��0٥�ф�y��'���'���*�i=�	?0bvUxџ�%�eh�4�,��G\��5�a�;�$�<ͧ�?!���?����?!���|���F1"��t�����T}�'7"�'��O6r+�:+a�!�s.	�-�|���.	듳?q���S�',0n����S�_�  ic
N)M^q!���M��O6y��M�~�|�V� #��B0_%�1`��)=�^����l��˟���͟�eyRL�>)�oM��˓2�VĩW���#������ �����o}R�''�w�"`�6F��X�ۂ.�%lOF���]�ep���8�f�%���2�	��� f�*�(1<����a�#t�y��3O����O���O(�D�O��?9�f`Y�LH1��n��؂����ӟpa�Oʓ}����|��b�TDXH��,�ơ�ҡ7��'N�]�����Q妵�'��E!(D�4>�1 ƞ �倲�T0�F��	+�'��ʟ��Iϟ��	�
�8�X��9 o0x"�8r4��Ɵܗ'f���?����?�*�l���� tUb����� L`��2��<b�O���9�)"��Չ���P��1\CX�8��L�2;6�h7Eِ%�́/O�i\��?93'7�$N�3�\���8Gn�K�!H�0����O��$�O���ɨ<��i��a1癅RT�<���ލ}Җ���'tb�'��7:�ɉ��$�O��$#�6o��c�D����Ҧ�O�$���7�(?Q����%ן@�W4���#D
\>��퓬J��M���D�O��d�O����O6��|�w�4bB`E����(a2��gg��ey��'��O��e���Dk�&8�W�t����8C'��d�O`�O1�0%�im�&�I?T ���fFMX��fd�f_�	�:Dfhش�O��O<��|R��]$��a��$3l��zQ����V5���?q��?�(O:��'=2�'��R�FY���!|�8��W��O*��'���'��'z �����УG�I8T�����O ��E�׷:�D7̈́L��*oq�d�O����P1�$\��dW�e���vG�O.���OP���O��}r��g�R�1�ɋ�-v��/�^X��a�O����O�|n�]�Ӽۂ�ϵh� �X���%�l=����<�����׹UZ6m,?QГ~+d�I�5(i�R��ǋ]�8���"�Ҩ�H>�-O0�d�O`���O��$�O���G#s������F�.]�@��<a�X�L�'7��	W�s��ܐ��d/r�S�k]� ��'����逌>�nT�t�׉&��䨕��!&ʴ�3�EJ#��/��(��n�O"��M>�.O��1��?�DT��)��F��eVM�O����O
���O�<�a^�t�ɉ�2A�%�ԅS��&��8|\�����M���m�>q���?q�9�n����ք,Wv,�6!�'���EX��M;�Ox���O����t�w]���c�+9çĝB�^(�'0�'r�'e��'�Р5�,5Tx{���}�� &�O`�d�O��'�I,�M+L>��英n"n����]7;��]�d�;���?���|R�Ã��MK�O�)z`��)j��|Å	�`�ip��$ ����YH��O��|���?I��[�6�+#��}��{1�������?�(O|�'@�	ɟܔO��5��C�HS�ĉ&(�ޅ��O�-�'{��?a�E"߃t�(�2h���0A�Y^�}k�O,~�������*��|#�+d��dᦤ)l�p��F��O'r�']2�'E��d_��ݴ(��#���6�͓�"�Y��	Γ�?a�p)�����K}�'b�8��J�V����åűQ�ű#�'�B��78(�v���b�է`����<�b�Ei�N)*�;]�-�3C��<�.O����O����O@��&��U>�h��x)�
���B�4�-�����O����OH���d�ަ�D�q��W�b���Ձ*b�j��Ih�S�'[ Ա�ݴ�yң�p�<3)̈vw�b���yR`I�1�Ƙ�� &�'�������I�s�,�*�/�<��)3*F�3~2E�I����	ʟL�'����?���?y�O��FVđ�CK�^�Hf���'��꓆?����1�	�2���0�i$%������'"	�3��El��+���$����+2�'n.��d눸*�1���C�q%�h;v�'���'���'s�>���h�8�6��.i��'�X�ZA8L��-��ħ<	g�i��O�V,u��hච� Z�x ��W�~�'���'ܚ�0P�i�I4��bP�O�\y��ªt�v@��c�\q��g��ly�O���'���'�2j� �����@(y 0
1d^6��I���$�<����O�|�B��t���-
��)��>y��?�H>�|2W�Ͳ|J�<����6<vr�����D��L٦$�n~"�	"{�x��ɔ]P�'��	��}�a�]!�`�vJ��g���	ܟ(��ԟ��i>E�'b�듛?�ЈT;�:�⭙�ISH�˶�ʋ�?���iP�OV��'��'B�K]F(*�b���0X�'O��Ha�i��	�<KVl�����)!��ܵMs��k�1"؄E��.n�X�I��p�	ݟH�������W&+Z��U����R6"-a&���?���?�dP���쟐B�4��Vx��9
D?
�����k�LqM>���?�'NS0��ڴ����Ix����hG�w^��qC[�r���PBa��~b�|\��������I���#�30Z%��
	�Ȉ��i�4��hy2m�>q��?���	��6��bs�[�{��$��,I��I�����O@�(��?���K�a����d�� !5�����>��d֦]����P?�J>��
{��0(L��[�(�A�?Y��?���?�|2)O�ul�!X>��qR�T�l�^��4�l���Iޟ�	�Ms�bʳ>1�l����j��s�>C$
3Έ����?F�3�M��O���'���RI?� ���H�yD��3,C1+�5(12O���?I���?���?����)�$>�(�hp�Y��	�`�ֳ���'�B�'�2��T�'+�cޝAE�-)Dr�A�� *�)X�O�����IM�)�9���l��<C��'J�p)ٷL=�{u(	�<y��F����1�䓇�4�����L�{�CB�g#��s��:G���Ox���O����ȟ���0�HP���R� �?Q��d!K`��s%�	�	�lg��7C\�J�x����A�x� �O���ppgZ�B�ѰI~�P��O����c�J��gͰ:F���2�H|��$H���?����?�-O>�I�ZàL1�lN*Ic܌{�� �2R�I�����O\���즉�?�;}H�My�D�#S(��z5a
�T\ϓ�?1���?�E��!�M;�OLM��E���d�	+z�9R
�Hަ( ��=^��'��i>M�I��������	SL�A������b��$K�!���'G����O��D�	j{`�����(|1��Y�L�(Su8��'M��'2ɧ�OɊ|9��.kn�1��S�І����/���O���K^'�?�%�-��<q��� N3
��B�U�������?����?I���?�'���H}��'�^��N����D�R�D���Q�'Tx6� ��:����O�ʓ-T>���@�P�.T�e�ٸ ��]HSCB��M+�O <Rw!��/=�����8�vBI�3�aB�ǝ�Y+�d�:O��D�O����O��$�O��?�@A��g�����P4�F!���ʟ�	ϟ���O�I�OUmN�	�U�X��NTK�.i� ��v�vy$���	��S>;���l�H~�a�5��]Ȕ�ɻf�bQ�d��iel]����D?�N>�,O��d�O����O^�#6�E�8~\��s�� .����O���<	"_��I��	]�D�M����V86�r�)D���dKn}��'���|ʟT�h@�O9���{��NL���.4���N_�r]�i>���'�d&�(��R�S*͋�"���a����I蟌�IƟb>q�'�J7�͋M�� q!
� ��A�H\�R��<�b�i��O�A�'�C������kԮn��1���I(��	�>��o�K~�)2`�B��S2M�ɞP�l���ʃy�!��m���{y��'���'���'Sҝ?-
p`��|wR{ ��%z�v��n}��'O��'���y�u���#A��Y����:rZ��@�E +�<���O$�O1�rlY�``����25�L!�Q͚rp`�B���*�牢u��!W�'� ,'�������'J� {%f��yi�	=q�����'"�'�X��H�O����O��$&�v�(%�	f�e��b�<`´����O6��OԓO\�@U`BE�&8�qO��h����Ɠ�DpF�^�l@h��1��*lE��˟����S7j.01�fA*gL����	ʟ�	���	��E��w;(�2s˗�@��I#ǡ>K3�t��'���?���B�f�4Ke�C�C���rЭ�M�L�Y4O8�ĸ<QcW�M��O�ia���beh�x�<`�Ů��K�d�K�I��?4ĒOn˓�?���?����?A�
�����)�
y��� Y�sd$�)O�M�'�2�'����'Ķ�PĂ.i������T�3���>I���?�N>�|���D
<T���&�#^d�A��I�(=��<RB�	a~��Ql]�IB��'n�I,1�9� �
p;u�P���<�	��X�	��i>Ք'�.든?1�A�k��!���:���A"�[�?s�i0�O��'��^��� �_�؂���>�ƴ�KQ�5mZm~��!,ol�S� ��O`woC))]�	V�ԓ>�4�J"����y��'��'���'��	�[*½S�J�o
<�[ǁJ	k����O��$Ew}T��Cٴ��<�8,�4-�H܍R�/N?cC�a�K>Q��?ͧ&3|�iٴ��D &K0�*��ߎ~Q��� kL�.CȌB��/�?�e+���<ͧ�?���?�0뚴<���2)�4f� 4�0�?����$�l}B�'Zr�'��S�T����%QVuc��?Y������ߟ���[�)��2D�9��̘ot	Bc�[�*l-���M��O�)S��~�|RaA�[���0 .DdR�,�c+ ~02�'���'���W���ٴf߰��G�!� C$�ʗ9r��?��t�����\}��'�ܤ��*�X:L�Ab�;Aa��?Y�*�6�k�4����������`y+O���ƎW���"�iCYQ��P?Od��?���?����?�����O�wؖ,�U��"~�*(���$�>����?1���O�$7=�$������QRd�!"�4sN�O\��>��	ՃK8�6�j����� ��*��O+�B(�6�x��"o�%��d �d�<��?1��.?�})Ҧ~��D������?y��?i�����L}��'�'k��e��;tH�<{AH@K�rE����o}b�'��|��K����2[�`��	���1��$�f���(�(P�f�1��� ��c� �䇲\���H��R�Y�̠^���D�Op���OL�D#ڧ�?'cT�W��J0#�%Q���qf���?�qV���IΟp��4���y7"H.A	v��Ѝ�.K
ͫ^�]��'i��'�fL�f��l(ԭZ a���  ��c�U<'�����9}�n�%( �ļ<�'�?9��?!��?)��K;B¨0;��Y������$`}�'��'��O��`�=<6�3���&�D�5�		�*��?�����Ş�U� 䅅A�2hB��Q�N  @�A��M�OD�K��A�~"�|�P���4�Z�)�X=��h�.ɒ�D������	͟��By�>Y��G�	ϕ.G7��`f�PC@T@�J��v�D|}��' �'�.a�wE��GX�q6�N,o��1�R�ql�����I3Ō2K�Q>��/Lu�I+ͩc8T�5'Z�P�������	�������}�'9J�i�$��i����b$��}P�����?��7v�i>�I�M[K>�c@m�L��Խ)r^]�D@	>�䓙?���|�E�ƫ�M�O��d�l�1Z7`�*k��	�Fթ*�$��'J2�H�BY����?�����o]M�ay�h�5鲜�� [�H�	Dybŵ>���?����ɂ$:?�T�#B	_�"ͪ���{���O"�'�b�'tɧ���';��8�h��wѾ�Yp��0i��9)v�H��ܕ*��������1�̓O�x��ޜ��0�ЭJ&�.eP��Oz�$�O����O1�ʓY��H�;iN�0�whԩdm��"g��y��'��x��⟄1�O��$�?g��<���
�!�	ȓ�S�L�r���O�H�~Ӻ�;O��˒����OU�h��,�1#�p�`&��)�&��'���ٟ��	Ɵ@������Iy��!U�.����v/�	�pp;"AO�.2��?���?�H~��V|��w��"W�p���r���'r:̉Cg�'`��|��t@mM��5O�M)q*/	�c�&F$`�ܑ�=O��B�[1�~r�|�]�������PBfZ�S��<�T̝&e0�!I�-��������I^y�>)���?y�l䊥{�b	�נ�A+^��N���rH�>y���?�I>����%?�9�ef�%���� HJ~���Kb 4��e��ΘOk"$�I�NRr���hGΩ C��!Jr
p�'㕏:{��'���'.��s޵Y�'�]�np� ���9���O؟X�O���O��lZC�Ӽ�� �vi2C��aP�R��<��?Q�s�(��4��d/�����'E��y
�C�>�l�G�	sl�h� 9�$�<ͧ�?���?1��?����%�0���k��TɓF�Ĉ���b}r�'��'P����1!�i�F��I���� 
}}��'�|����f�����6���ANҒ��0��i6�˓r��x]�~��|�Z�0��I:7`\1�Aꅃ*gJ�Y�����Iğ��Iݟ��wy���>I�]�8E�"��g�]h��^�#	J���-����J}��''��'��Y1�\ z��aq��(,����"3p��������Ai��+����,x�S��|df%:����nE�g:O���Ov���OF���O�?!JFHY�AXGf�� D��⟤�	ǟ0�O�	�O\�oZR�	67&�z���c$��êӀr�A'����П�j���oZx~��߀Ip6���l��dQ����7��F�>�F�D��䓿�4�n���O`��ɋ"Y�B�
=:~����S%5���d�O�˓W����X�	͟\�OLI1S�
)k�N�a�K�|[����O���'�2��?!rD��TwLi���R1<�ة�U E"G�q��"՗x�F4���I�˟4A�'�軶�'�����NϤ�ܘ��"v[G�'�b�'`2���O-�	=�MۥIP�t� ł"�n̤`�$K��<Q��?�мi��'Q��>���=M� `���G�=H�Đ-6ȵR��?������M�'���&E�f1�#���D'4jv=[�n����%kD*R�w>�D�<y���?���?9���?i,�r�we҈I��Ɋ5�:C���K6�P}�_��Io�'9���w�"4Aq
֛p� <�e�J)3&� �`�'�R�|��dI[�&:O6��WF��B�̛�*�2����?O09�`N<�?q��!�D�<y��?	Z��"@cT�ú�̐���O(���O����<)ES����������$��u��2J6���b_O,Z��?��Y����ڟ�'�����ضP�r� �&L ��$O.?q�F�lV	"f	�1��'nX�D���?Y��`�"T��ʆ�O���Q֡��?��?���?A����O�ՙ�mڗz1�$�ec��X��g�O���'a�I��M��w�`���&�UN�A1c��S<.�(�'���'7"d,ϛ����%�
,�$�C�"�Yh���X�t릊� =�!'�x����'Z��'���'�~��jɘGg��£�ܫ��7\�X��O����OT��,���O6p!�i2{+:���Ō�!l6d�s��V}��'&2�|��$*f(�0p(/�� �U�!$Lh j&�i��	�#���1�O�O�ʓu����Q�	��EAч�3�x1����?y���?q��|
+O�4�'�r��0 �c�$�(�J�vaV>�y2�bӐ��Ox���O
���y2��zAh��2(`u�Y�<���t�`�f������J�L~���j0��K��0<���A �!�L��?)���?���?�����O�M�`��\�SmB�+��C�P�p�	����?�R�4��s1��c�.�u��%C�R=��<�����D�H 6-=?�0�s�? VX��C7�4��e� �4��5�?i1i*�$�<���?���?qQAw�����_tȘKw���?I�����U}��'n"�'��S~��Q�81J�[� �\�P�nv������	`�)��/	��Qv�܏+Sf1r�;Z��p3m��C��-���G����[d�|��1������V86��I��%Ȳt���'�"�'d���\� kݴmLiu��( ��y`A�W�����?��]������y}��'eva��
:9"Hx"d+��@V�'0b�=�6��Ĩb��q�$0GP��0�{&.��qH�"0<O��?��?i��?�����iH7{Bщ�	(���"���'T��'�b����'�6=�� �+:XLjWJSNF� U��O���$����Q�6-t�03d��<&m ��3�\Q",v��c��!u�˅P�Iiy�O��`�R��4��Ԧ4p$��H�R?��'`�'F�ɦ��D�O��d�Ot���$(Y�L"���?
^0�$�7�I$��$�O �d=�����yST�IgƉ��*V����΀c�O5T �c>�kG�'*�5�	�� k��H|�dU�'���l����������h��O�O��H0]Npa��,K�ֽ�&N�(H��g�>�.OBm�_�Ӽ���]�Z<%['�"����<����?a�$!�U0ٴ��ą�lŬa��'s�J��K^8e��\��F��y_�d�ŀ$�$�<ͧ�?)��?���?qė�	��X�e��� -�f�ؿ��Z}��'���'z񟮽�6+��
aV�h�bWx�
8��(MZ}��'�Ґ|����V�i���v�4t64�`q����S�id���s�Z8p�O�Oʓ�����5R�J��fwX1����?q��?!��|�(OBA�'�+�)SN���+Ɵ�X��3�['D��/q�v�y�OF�d�Or�$I \T��Ja ����S��ܴc�R�w�d�s�%���?a%?)���)��l���η�T�`�薑	������Iş���ޟȗ��OCع@$m��O:����^�Z�^,��'��'����|��BG��|�,Bk�(�8B1j�Q��K��'*������۪yt�星0�0��=��r3Ȓ-h&Ȫ ؿM��x�C�On�O���|b��?)�	FH2���k�J� �C]+(�f[��?�/O¤�'Z�	�D�O�d< �◘�rH1��ȕb���Ol��'@��'.ɧ�I�2V��i3��T�y���Sud��7�p)��W�'��%�Ǘ���+<J2��\�	�
^<3�RA��ˢ�ٰh.nT�	ʟ���㟐�)�Sjyүd�����z$iBcS�1W�Q�3O`���OR�l�Z��K!�Iğ !EG�/ ��ٲ�B�g���ʟ��I�w��mZ~~��:l�|�����t3m��B9=���ɓ�4���Wy�'���'w��')�_>��GE�:n�ӁJܖ[���cM����O���On����Dܦ睺r�q!JbI���ÃO�,q���	���%�b>�2�Φ���b�:��'ƀla�*ߞa��=��X �r���(&�l�'���'��d05��	
�rJR	�I���'FR�'�BY��)�O ���OL��ؐ�EN'����3>��ģ�O��D'�ɷ+�%�u`�&tz�����%5�M� 
�F�9'K`�L~R���Oj���xxx�g��8Op�j�OY3'ٚj���?���?���h���$���|e�e�F�q��`��2lT���PZ}"�'r�w���]�\�u���'�z��ѮX""}z�I矀��۟��jB����uw�X'#z�䡛�O�L$:�Y�@T(=S!H1rl,&�,�'���'���'���'��i���S!rV��b��J�P��j�[��i�O��D�O
�D*�S�h��(҆��+�D�S T<kQh̻�Od�$�O�O1�܌t�II��kr �gTH��TN�]�.6��hyR*\�r�j�������Q�{���i׫��H�� �pn������Oh���OD�4�vʓ0�I�����<���+&ƥS��
ŧ��8�۴��'0�꓋?�)O:��w@#l,���"��3"��5&"6N�6�4?JјK������'ϿC���	z��ӇiL	��(�J�<����?���?����?��tkT?��uP��B��P`�$�]����lèO�I�OHl�t�#[H��j�[ne���iOm��&���I՟擙w�ʵm�t~�Ȗ�m��|��B��5Le`Bh0ў���
W?iJ>�-O��O����OL�Z���+"f`��#\
���.�O:���<��T�|�	ɟ4�	`�#��>�^�qC$4ݠ�I���D�F}��'�"�|ʟ�0�`+�?h�P�[�j��c9@	����%��	�f��`�i>���'�:(&��k�*�F#h��;ixbb�������I�b>�'�:7M�<o��$�^�*�������<�i�O<��'B�(
>f�T��
ݶJ��. #Nn�ɶI�>l]~�˨.�����`��	�a���HκKk�(��#L��~y��'r�'���'��W>yZ��&J%Tiu,ͩ0���%$˫����OH�$�O2��J�d���|���!��(���0` ��K�������&�b>m�Ц	�S�? �h(���5(��@�C���L�?O�1��b��?!�/(�$�<ͧ�?���[)> ��_�Ti�3E���?����?����YF}R�'_B�'?v9�eZ,
�r$m1K8�H���P^}��';�O@�A�P�x�
���۝�a�P��`�,�uV8� !�Q�pR!�ß��uĉK�$��%��"UxT�
RhDȟ��I͟L�I���E���'�u*�HIw�:f�Ӕ�t��'����?��Q����4��1�
3\��(K5I���077O����O�iD"�@�i�i�4#_����j�5=Z��KA�W8���ݳ|��X'�����'v��'���'}6�)F-
�vK�,ta˂$���U��)�O����O���)���O `�eF�S���GY8pBHE�"�E@}B�'�|����ύP�8A����o���`ĊʮgNa�&�����G'ژ��'ܰ�O�ʓ��(�b%��R����B�<x0���?����?��|B*O�u�'%�*��|ּ�[�\,򲥉�M��2X��D�W}��'[��'x �R��[+�P����RĨLJ�F� C��&���2,���t�I���Yנ� = .�1-�q�e4O����O*�D�O���OH�?%��OD�= ���a�&*X�Gß�I۟�B�O�l7���|��v�2�e��b� `Ь��''\�z�(�����'NN�a��������D�B�6��k��q%���\H��|RU�$������	ݟ�Z��(�έQ�i�fA�B�����	OyN�>���?y�����A��t+L[�T� 
�lt�ɷ���Oz��S��L��L�4\����B��q�͗z�9���:�P�x�S�_E@P�I"@��l�C�tv^Q�Oݦuʮp�	ПD�� �)��Dy�v�yd� ���B��&D��T6O����O�pl�Z��s����k�털(5V�ّ�u�|d�Ռ�ߟ����y��m�b~ZwoV����O�|D�'C� #wنX���#���H�'���؟���ٟ��	ϟ���p�T��Jl������O~�Y����j^듞?i��?!I~�aJ��w=THa�h�z�ء� �@D�� ���'.��|��$�i՛�0O�r��Q�]�Hؠ!Px�|�=O��%��?Q��(��<ͧ�?����VQʠC�>���A��˪�?���?A���N}��'���'����c+ t�&BbT  R��D�E}�'��|����(C5�ފesL�;uL��$Ƚ8�P`W蕄�H��zh)������M�H^88��Ԫ��}Yb&;1�����O���O���)�'�?��/Y�̠�B@��EE�<u]*��� ����O��ě��?�;:��]��˦�ڙۄ#
�����?)���?�`ҡ�M�O�n
	���I޵],�:��!|
�QL�!6>�I�O>I-O����O�D�O���O��"�㏣e��\3¬:Q��SpL�<Ir^���Iݟ���_�ݟX�r�O��>��+�%̭{Q�����O��d<��i��3����L*X:v1�R���uԽ6 r�4�ʊ8�n���%���'3D�£�>�$MF��}������'f��'^���DR���On�KY�������� Z�n��m�I��M��2�>)����$�)�>��" I:_�|��L�gr��!�n�l�}H�mQ*៪H~Z��?�T�؆|Ռ��fʁ06zB���?Q���?����?�����OJ:$�ebֿgE��{Qc�_�؀i��'%��'F�S���z��O4uI�#Z2PZ���1;�P�����OP�	����4��dS�??�:�@C�x�\Q �� \�ȑq�A�*�?��.#�į<���?����?�SJB�\�֔�T*3���J�?�����$g}R�'T��'��S�ew�h�F�2j��ȇ���Ơ�;
���	F�)�N,~��`\�Jk��:%���p��"Bk��M�]�擔Z��2����&ls$�$?�4yq*�<Jx�d�O.���O���ɺ<�c�i~����2ul���L�:��,
�'���'4�6�6��"����OZ������+`F�	��Hڕ�楹<��O�
�M;�O��&��1��<GoL�#T~����G�,@�Ti���<!*O��d�O��D�O0���O��'n|� ���hT�S@˝�ͮy�U�H�	��	O�SLZ����gG֓qq�x�t�FjбB"����?���S�'h��T;�4�y�,H*���H���!9�>�S�e���y�
^�T���s��\ 9*:})�k�<�)ƯH;��ur�#ђ�> API.��� ����Ā��T?y�� �H�	:3�i�b�~��т�C�@���@�	6�>O8��E�S�����C�!�}��Z��R �K�Oy��TiϨ7nQa4�$䐄T&K�K��<�a�EdL��M׌f�9��1!����GW'�\}���M�	.��"�e�q��AJؒC�4x �
+8In�{B\�E�b�1�-ʠt�r�h���)3jٯp���H��!_��pqfFZ�"���g�Ó[:�hӎ���O�u��-G6Js����	��I�������	H��������.)�I2��K/ӛ6P(2�[�)�L7��O���<����i�O�d�O$���	/\H��ٳ�߆}b�93bm[e���D�	v�v�IR�~be# 1)�ԉ��bR�k$� [����'�ny�~���O��d�OR ק5���0�bT�̟$��i�V���M��?1�R)��'q�� 6�����>�"G� :&>]3��i���h���O��D�ON��';�ɴ8[�j����l�@�9t�g
�+شP�������O�5{����*�ReqKN���iJ� �Ȧ�I���I՟ 	�OP��?Y�'����"�(y�8pH�NL�2�qX�}���Y�',2�'+B��/]P�C��/u�X!�-�o��7��Ob�$�K}r_����J�i�M�G���6tH�(���(�>9���8�?I-O��$�O��5�4��8M�<��Ʋ6�DJt��/�M� W�8�'>2�|�'?��ֱ�.q�glʜN�P����]'$�a�|��'B�'��O�"��n�$��+�.@�����FN6DZ7�<)����?!��f��'�<e�'���)�/s;�Y��g�	����O0���ONX&>Y)��F��RF\�RF�x�Z� f$^�&n��D$�H����!�lɟ��O��P�Ѭ"��#�"��D�>)E�i9�'����3�����O$�Ӽi�ڑɢK�x:�2(��l@O���OH��r�9��[:w�R�.=(tx�`�pB�8"�a¦Y�'��qӖ�D�O*�d�ON8֧5&A	�vC��#��	�y�6��h�M+���?ѧ��'q�\}
��N�QL�-e���X��M��6���'h��'Bʡ>i+O =q�E�-���7�Nm�Z�12k�Ʀ����U}����OS2��6w�b誢�T�t�Н��Ŋ(N�<7-�O��D�O��$Kg}�\�d��^?�1��L�����+R��H�6�Z�	L*�HM>����?��C��ӍA!�;F�C���)H�it"�'/NO�K�ɝnX����fĒ����ɘ\��̀K<Q�����O����O��O�\咗���O�T��C,� S�!۴(�'��'R�'�i��P� �H1���`y���h�R�ĸ<���?����'ID���(��9gŞ\� l�H��lZ�I�����g�	xy�O��G�?ڶ�ר�T�� ��Nq�O��D�<�.O4�'�?I�MZ��A0aS�Pf`�V?ߛV���O��/���&�p�P�/$ hK�DY,N�[�x�F�D�<�(O(ʧ�?���?�1l��'��u`<� EA�>�&����By��z�O뎂>�UW��P��-_�'��'�����ɟ(�	����u7cYCs����� ��Y"��*�M����$�63j���	)�Hd�[� c����W�t����p�	ϟ��	gyʟ��+�	�H�a9�&�0��0A,PX}����O>�a��\g}���Sn�|U*:�N��M{��?��?�.O�Sa���PfRݻ厔2)S2�HWO�@�lEx��'�S������h�'�{&���Ƅ��N5��lZ���	ryl�~���M�/xZ�HU��p�,��z4O�����������	N��Śx&�8���:�ARA'ހf���$���O�d�O�ʓ�?i�Op��Ң�
Ѩ�ÕǍ�2�&؉۴�?1(O&���O�����?QG��+ [J!�T�2v��*n2���'@�$�O�˓�rUl�	�ε���
����E-HN�듖?���?y���T�1��9�Z|h@gƧ-�H���Ѕmt.�nZ۟�$�X�����'��hu��1a�I2�:I��1m�`��syR�'l��:���Ok,\2a&�#dN �T�v��V��_�'��I��k�s�֝�w�Z�3�F�[D������&G^7��<��	��6�'�"�'���>��\�<D�p��\h��!��C(dO
�n�ǟ��I�N��ICy�'[q�����E��zU��b!��he�p���i���j�2�$�O���O��	�O^���O}I#GR5	�@�@;�A�͛Ϧ���@ٟ ��ay�Oe�O�r*�7/T�y��X��x��2JL6��O"�d�O��DVɦ��������ϟ��i�]�G�5 ~x��b�,${�U�Bp���?%�C�<�O�'�R��#x��rI��k�@PL"1�6��O��d|}�Z�X�	`y���5ƫ >/g8I�dH�w�$ٚr����d�9S�D�<	��?�����/B�R����
��=~'�%��iT듄��O��?���?y4�͝E�q7�����ua�\3#�1͓�?����?q���?Q/O���|�Q�ҧ>���6LY�=N�P�Ǎ��q�'�2U�t������I�yjx�':�޸Z�ˮjD�`3Ǒ� dl�۟���ڟT��Ly�O�X�'�?�1%�(�ChK�6�~53uK�)n��oZş �'���'2O��仟3v�PcBKO�{Bdѡ��N�gz�7�OR�d�<����ҟ���ȟ\��'�G���ǯa��t������O|��Oj���=O��O~��fi�Ebc�����qP���7�<�eg���'`r�'�"��>��3��ɕ抸QT|��AH"��Ho�ӟX�Ih4�	[�Io�'N����� �������i��4o�ҟ���4�?���?Y�~�IEy�DF��6C�*C��4�B7k�!y�7-�(%��\���h�;b��4x�p���EK�k&!D�i\��';r�'|������O���=`r���	#`q���1J�&k�7-�O���O<���2O�ҟ���֟��� P�CF��{ �#WXvLb�i�r�'xx�����O�ʓ�?�1):N�˴�!���G�'���nZ�pB
h�h��՟x�������F�\ce"�*$M,"5�P
�y� �ߴ/���';r�'��İ~".OL��ݵc�|]�R E;�Ȑ.�>O!
��>OZ�d�Op���O���Oʧvś��Z�b���ĨS95R�M �-�y[N7m�O
�d�O��D�Ox��?��B]�|�.���P���0���`d��8@��F�'�B�'��1�Z�5��⟸����)�����i�#'�ݡFN��M+���?q����O��<��'�!�W�q# ����a�hр޴�?�������O\��OJ��'nb�Ԛ�4$`&lN2`s����(R�I���?���?Y!E�P~W�(�'q�q�c��<~�9)��K�z��mby2�'�7��O ���O&�Ka}Zw�Z`��V+6�4y��"�'9Nt��۴�?a�;���Yz�s�t�}:�B�$���A�O�/ajr��1�@ۦ��	*�M���?!��?�rV��'+�ɈPjQ/���c@�W�!��F�l��6�U����<1���'�:��T�}�"�C�������M��M��?���?�#T� �'qb�Of�IQ*p>x�UW�|��3�i.�'����i�Od���OP����)Ov��e��gn��ԀӦ���ş�x�O�ʓ�?!)O���� 9E�Ьp���P	?��aRV��@c+?q���?����?�)O�N���D� ([LYx$Sz����>�*O����<���?1���ܹ�q�ÕO�:+G  ~F��\~B�'���'�Y�擅��d�C?��}�ԦV�,o��*c��M+O��$�<��?���Yא�ϓ3~�� �`F)x����ïAZ2@[��i���'���'��i>]I����d]D�8)�؇Pl�`��bz�\�d�<����?y�7�4��>Q��Y�kf�� ʊ(�0�� ��Ǧ��I�@�'r¹~����?9��o� A(�)��7���SQ��+>q���TS����ʟ����KvT���ĳ?=���opЕ�_n��PC�f�\ʓ�?Y0�i�R�'q2�'���Ӻ۵bZ+5!0h��J83�8�j�KĦI�IƟ�H);?�.O��>i��H�Y��-hC���M���dtӮ�d���a�Iş����,�O:�kE��fbI�B<���ʍ8]�|��G�i"|dӞ's�'������N)" � ��9����L�D�mП��I՟�������<a���~"%��Q:<�$x�x �4i	�Sw")mZ󟌗'��J�����O���O���kR�B�l9�@�E��*0��m�䟼�ɮ��$�<q����Ok�>d[�E��ٴW�(`&��	-�ɗݤ�I�D�I��h�����u׬az���3���9��$��M\���'+2Y����韨�	!z�auI[�d&D���J$ܾ��c�p���	�����؟ �	Ny�O���++������w(9�T�V�3q�6-�<�����O��D�O���6O�	x���"�:5(
{}�����%�	ҟ���蟸����k/񩁴PQ|�cA�=,SFP� m��m���L'������X(�G�ȟ�O-�g�v1�2ȕ+r��,; �i��'V�����K|*��?��<"������U�Ȃ�	�#d�'%�'0�`��Ĩ?��ŋ�#e)��f��u��j�z˓�?ّ�iL��'�?���a��	�r53G�ֵ/��7"\4$�0|oZğ�I�����G��cܧi�\��˕�[����U!��F��]o���i�4�?����?!�F�'�R�
%9\Ir�/��Ra�b8||\7mGQ��*��+�Sޟ qt�ĶY��PX3�J�3� ��M����?Q���?aD�x��'���Oh��\�0:���"d�p��i��'��T���'��ݟ���ҟ�6��S�AE�
X�y�C`19+6M�O��p��?�M>��G�jPr6��v�����0\���'�x�S��'�	̟p��؟h��29��:�4}"��qL�Qې�iNdO��D�O��O��d�O�`҂IRn8����Τ/@� ���ӕP�&��<Y���?�����':T��"< ۢ�3V` HDc F�	ן4��d�Iן0��$�"����R$!֠��#S���b�\.s��2�O(���OH��y�S��ħ&�����&�+U�iI�CT g0��i|��|�'}2*�y>���� #i�E��` "�<a�C�æi�I��'�� ���O8��� ���X`��
=�	c!�`�'���Iʟ8�e����%���'c���B�FN�Q�f�����s��ho�YyR�'�6�v��'�r�!?�B�_�h�Y��Ia���gHG������������$�b?��0��I��5�����jcr�J�ĚզM�����I񟸨�}B���?\(D(։{_���7n��L�۴D���2������O���=L� �c���&'G��B%����7��O4�d�OD�d�~�џ��J?�ŕ4J�P �J�8@��W|�#0j��M>��?���W�`Aa�e	�j���pBD�#�	Z%�iMR�'�HO�:�o��e�˔��Œu�Z�Rl�%����}~�-Ԩ-Vs�?}�V)0a�Y�u��0�w�L�%q�)�DiȯQ4X��	�cs�$:Ӆ�B���
�Ā%���Z��G�	) I��oŵ:9��0��_��%��!���G"�"<8�ݣB+Z@���� L�t0Z}"CB�: ��q��P/?h�P�E��A9�O�g�� ����ԥ`�:�C�R�{����-��w9d��(δ ¥js� �*I�T�ۻ\�����_�8d0�r(��[a"5��V%^Ȃ��M�#�s��Q4.^D1�̷}�0�"�eů:O4����ۿ2�p���/6W���#�ު"�%�AJ�V)��X���R�_�<	��?1�m�$%e�
�+�	'��>�O��˝&:��K�iT$N�,`y���ȍ-�ά#�� [bP�}�EL�T��)�*%sr�b�
C�'��0���?��t��0h��@&U
MC�D�6���y��'۴�HG�	)��0jӎ]�&���/d�'N��[@�ʆ}�  �4L>�R�И'�z�$�>������?���?1i\�ar��:P4���j� ;��#�.@�|�*VV+�*��c>���e�v� ��^���Yє�ZP!�OJG(6�ZaK�{0r��)�� �� 4qQ��qb� 1�ʕ�WC��SH��I՟��䧃�k:�����68e�ķ\vД��Z�:)rЩ_�=�-�d�߶$� HDxb+#�S�4N���<���w�N���N�9�R�'�0��f�t���d�O����<A���?�cX_����@�\3V�¸��ng?1�c[���SdD�A��x���'�UJ��0x��������~�M_�KZA��	P�<P��P�#T,1'��.���aߣ���I9a���'�ў$�'kV�'6g 	5�%|m���
�'�L�a�k��LHl3O�r*�!�$;�S�U�`�˝,�M�E�9p�����ݢJT��a!����(�I��'���'����X^��MУT�v�	�Ɣ
XH�hU<X@�\p�JC؞��D,ŏ<Μ�h�b�-kQ�
'l�v�-��j�tntd���^��	�%
u��0sA�k��K�L	b�'�џT��@Tj���C1�B���$D�̢�H�0j�&麔��)��1K%jp��X�O~˓	��h�Z���Iy��E�Q��������³�yb�'@2�'P��
c�Ȍh�р��T}*�t=��,��U�R�11�(���g剋$Ҧ�����E��@8��4�^�K�p�(2*��A�����(O��D�'y"����S�D����֮+:�	X�6O���$E) 긡!e[�S!4��g�J�a|R�:��	F�l�nѡX2ի�B��l�D��l�����h�埸�������N(l�a��+��V�����k�=T�(4�eLQ��ē��)+�9OFuq�E�7+�J'��M*0 ec�N4ȑ����;D^TA��n�"~�I�?#B	�bd�?	B&�����?�:��#"�����i��&�';?�䊕��-A�T��T�E�6��O�˓��<�G���nB��(?lQRL#�ÆJ�'ě�`Ӿ�}B��J}��k�!Q�0��2S�B=�?���ȶ�1�ij��'��S��ɟ�z���=80�c�(����i�f~�����,L��t#�K3LO����1/g`�q �1���;&oR�*����&V3f��"i��P�����4b��r���]1ഁr�«D_]rv���4�N˟\�ɰ�M�gy"�'�剓�lIZ�*F7"�&ಥ��1R2�C�	�t���#+�>�ta�N�vX"�Q�4�?)H>�,��ʓ
��̻�������pj8l�%��t��)���?�����4���v>��@�=zY�LZa U|�V�pt$9PS�;��|�E�:]�L��4[
e6!pal�;krD���ݠVnJ��	v�����O��Q �(U�b`I� ڀ���i� �O���<)�������L��	�/�&�ޭ`�IU:	�!�d	Q��H�ޢ�.���G_�k��D������Ey2����7��OR���|:�.��WJP�2��cwH,Z�.I�<!��?9��M�L���Ҙ��g�0�"��t	�$M4J�Q�\�G4��.s$���h�"��)V�1�a�:��e�Ig�OxX��Z%�|�ah�i#~ �	�'tq¤�G<u��P��
4�z���bX�'0�i�@㑼>G�@����(y0�'�jL�b�o�@���O���B���O����a��u#FU n!X���7#>�au��O`b��g�'j�HQ�?&*8�1)8R*�2�A��"Q�"~��68 �Il^Id 
�C���
h�cZ؟��<E���%�����=f�� �@a܂���'�:���կ@�{��/Fm�h;��DR`���)�)2x����
��uhz����0v�v�D�ON @Q��Ц]�I�D��Myb��y�'=����� �
|����{4�U⒉؈6e|4PK-�h���O���<١/[��� �tNU<y.�P�OH�9�p���|��E�Č�k�\��'aQ�(�vb�����	���R0t��"��x@��O��&���.'�&���O��*��Os?��S�? ц�OhZ�� d6n>8��Sg���	�<i.��<��`��8-
�㚢+���3DC��?���?9*Of�$�O��S+0�D�OJ�I� !_������9cY�5�'�'�T�p-O����?��q�� �+H,��J��'�"�����?��W�	����� 	����-�:�?������O���'_W�$����=9`�������ȓ\��{f��i��sE�Ip�=�����'��I�"s����	柬�O}����cށd͊�:��t��[�'7r�'Bf֤Cb�T>-[�(Ps5�}[
\�Q�\x�C�(��T�F�Ƈ����ִ�б��"	R��Ē!%d��.5%��V����"��8,҄B�ɻ W��cG�m�V��S��kZ\���Kc�	 ��(��ڊH�0p��C�
06�I�PxЩ�ܴ�?����'�?	���TQ4X���w�\�9�R�JЧ��R������������7�@�K��ȈI��U�׃��6}˓��e����e^8~�����~��԰��B1DQ���'�1O?��F
}8�9��/2�����E|!�ď~/�@*Uf�&x�V1@����k��Hj���?!��t"���DX���5�6D�(�i�09`��P��5z�-�4D�@�VȌ7=(X��	�/4�.]��-1D�jA�*\��Qcu���_���.D�XwN�x
D������i�c9D�<'k��I���TDJ�Y!��/9D��Y"�x�� 9у]����[u�*D�I����Dy���ș*���S#D�4�S���*e�rgX�6������ D�d���a<��h�K\"�,��s�3D���)�;})��8ǆ�'\$��-2D��!7���d<���+)+(Tc��2D��:28v�2�K_2��h-D���v��tO�4qW`�6>BX5�M*D����l�'��(a�ܷ9�\��0�=D����lǫI���� h�X���:D��)& -\B�!�kU�r\�p�:D�43����cU"��qhX{�J�1�G:D�tӅo�.B�p�`��k�.�Q�@5D�y�У|� ���݈D�@��1D�@�0䎌qA&��SN[�zd�O"D�`��K@��r�0�L[)9$����i:D��ת@$lL�i4/Y�u�H5�:D�ph0�#���!���5K(���b:D��J����XՒ�C�8s��!�j6D� �� ��&-�%@`��W7���$1D�D���"u��9��_�$8�|{w�-D���Pi��2�5yQ�ݑB>uia*D�ԓ�E��6|ꃨ>Ts
��qD)D��sT��%$�F�����@���M%D���YexBd�$�@������#D�x9���f�,prc��e�
�x4�4D�|�._
�t����� �oc�<�C%)~`𐑡�TI�v��'��V�<�2�	9�m=�0&Km�ʀj��V�<ad慍Y�0�Р������U�<i�̒0(�J�	�369�����RK�<QR,�XODx��E�O���P�GND�<���,|��X2�4�!#1b�y�<����r��� EQQq��*��^�<9�JT�3��)��K�(9l��LZ�<��T�w�"��M�'�h|���Fn�<郮L�%��b��<fE�Qp$�k�<��3��b7h�!�$P`���g�<y�'C$t�`�C�EH�"DjT���d�<!��Nl��@T#*H`z&�`�<� �pc�ڴ8E8���ET�`2�\��"OZ���d&��ݨEK�F0���R"O�q�E�֥�@o�p*�ܹt�'�#�	)������X�fT��	v��$wAC�IT��Q����N�����j�3?C�'�nQcsI�|�S��5s����	C�ִ��mV�Cl����~t4�D�ܹ[�4�P� M=ZP,�=�) ��@�TH���E�.�D �DM� ��$N( O�9R��,	P]+`m�!On� bpĞ!�x"	_;&<�kǬ�/y�xP�M��<�W�X[�1Ox-�� ُ5<Ҙ.˸Q���"O&� ��;W�^؊��
���"O4�%�J�J��(نl��:�D"O�H����ZӺ��pl �]I�qZ%"OЅ1a�C�*Ĳd����^f���"O�i P;p�r�1#�M�Je���"O��f�3?案g`X?TR@� "OJ��a��-f bjáěTL��1"Oa10a�*8j� y� �A�(ʥ"Oj�xF��
�H�5.������"O���ҫ#<�h��O?���ۥ"O4u��.�z����K_{ܠ�"O���ICm�"$�M�\���C�"O*tB!�,Y:� �ΟͲ�@"O��!�?J�<�V�O>Vbe��
OJ��M�#h��$��;W2 ��`H�\B�IH0�qbñ�H�P��{������S��t�{�[ #�t����[�IN�q���=�yBb�#��!g��H9�Q�(>��D�
r塈{���H�~�ę�+�8tb5���9,�!��X�u��a0���M�4�a��5Z
1O4�c���p<y��S���	q�[�{Z�#�J�|8�hjцL
s޹��념q��aJ��ē7i��
+9w^	���.a~��|[�-�N��$�5.F�O�����#y��Y0b�.$�H*!�?`s���QT��	��.4���t(D����s�~�*7�� ��1��O��{)z�s3�F�2SP8
�,G��w�"�X�A���h����-��'; ��nL��p���b9L]�K����Mk� ,P�R ��ۃ6	��x�'/z��qAP���)�;~�,���`�|DH�k4���
Bn@iJ2��H����P��2��#���d3���'-$5·�R�zO�c'��!E~,�O>a#��%a�~-�SJC8{.4���^~�OÞ�e$дFۜ���.ۇ7��	�'�l�2ȟ!D�(�0Ś$F42�QB��6n�8  �+#ѬH䧘Ohe�<�|D���.O�R�ӲjX,^e8�8�O|h*6n8B�!�c�C0]n��0d��<I��1OAt�sˀj����p�'�.��gO�����!��v�F��ӓ���Wm�3#|A�s�N#DN1(��ǥ
��Hƃ4U#:�2F���|]�h8�O>1�Ӧ�Ńv��آT��Md6(��D�
�M�&�/b��ԟ6p��D� 5񄸣uB_�!�XԐ'"O\9��-.�F, �C�"��1X4υ����d�"p�$)�P��>ia�`n��*�`�	HP��I��ƉW��� D��y(��	�yKq��?�XԄ�<��%���X$hA3~�� ȤkPb�'w\$�U��'r������8�t{ד\b>}2f(��A]��s�LF]��]��,@��iwkI�I~���Q'�p�� `�'����l�a`�j�4#,���{2M�1VI�آ��Ɨ ����H3��ԟN�@nD�^��-ڷ	��y4��0T"O�X�� s����UR�8��䫕șha�0s�H�u ԉ�g^��y��)a��6�:C h�u�];��ӑ2D�lkpm�*�(�0"�O�@��y����FW��.c��5{L�WX
�i�
?JQ�t"MB%q��YB�^�_��D�Ǐ.�O���C,�>�:��"�_ VRhL�֧��n�T�b�M<yf�`!��.�
��
�;�bL�e�>1��=6�SV�F��>�P�şQi���5M��uz��X�$�P?��jF��BM�7��P �i�p�����zǢ\R#+I鶹z�A��d�s$�%�����f��7�%+��QƟ�|�{�? ̋��ڥy�XL��i
!><t�"OBI����t瞅W���|hh�$�Lߛ��̓0`*��k�/MM���HO~�2�	��2��t1�&X<�R���'A�᳑��z�0L��Jr��9��ߊ0���
2Ĝ�wCd9� O�cJ�����R�F
�7*_�͛ �'����@��B��9�5�/Ծ�3It����p�������&"@V#ĂCp	pC�	72 9�!.��v_h�!
�j�$q#���\bB�h󍖰_" }�2F"�矴QJP+,V��	��?�}x��0D��`�/H$���'6*j��� .�v�j����'8:m��.]-!��9��C�BV2�8�'�:l˥�/�R(�t�4Q ��	�8Z\� �,��L�}�'ޣL5dm�G���V��3���0<�%c�e��"�Y����@ ���*(Wl܈��H�F���<�*xx�@ڹP�4A�II�=�'!,�k��-t�=9OE%O�I9�t�'K�Tl`G�@�l�2G'[��Q�ȓ�h86�̦b<hj抳  Л��'C�m(�ȓƦ]s� ��Om�O2��&�!Guj4x�@!=5�O2�Y��-�e/ǅC�9�!�ܛU���D.�"~b}zP&�#_�μ[ab(,O^`� O۟J�j��D%e!�S��'Z�UHP�_�`�((	����u��@��؊ N�1q���7ذm!e�0 �B�	�1��2яЈ<�&@3���/B:�9�S}�ʧdO�O���o�:��60�����*͌w��qض�K	X-�B≉1�� c@���_ � ��c�!n�e+�}b�K':Y�x���GC~���L���Z�(�����jO0��0�_8q3�qE~B!(ݜTy���	}�e��M�gm�fX�1`�+?FTqiŎI�~�F���c�%^���gL�lay�.�� t� ��=F(ƽ	e���yB��@0
�a�j̻f��s�&����O��H��"{��pŨ�D�&��ahH<	��>$��@�%ʻ,S��'G� ���AV�d�'ߢ��6-��8Bp��;
b���Ǉ�?�NM��.�"1��	7QrcՂ�<l���J�Aj�;�$3-���P�����}��i�/>�J�
V�o��0Ѷ����07sF��r�(+�Ҵe.9�a�q1c�
wB�`5 ]f���	r�  8����\1�G�"jj�cc�7�̠�U�j��(l�pd<@Bt�	N?v�;�ܕ.���z��
O�\�ɑ/`�uPd�;��y0��_;΢=IN9v(@�AukB�� �ᐇ�McG
3�~��$��'���dC�b��]�!a�.p39y�	���6�DzZwE��4K�"`f�ݒk�2�P!N��!Y����a��B�I�L�Th۔��,(�  Sŀ$<�T���$��d~0�Ҳ!�
�PIC��?�AuӐ�svL�'8t���D�Ut4�2��'����@�E-E�4�0�;OD��ȟv�A�'ű<0��P�i����^Ht��:�fx��T8g"b��Ma8�@3��#lO�h�&8(��y*�#d�Y�vF��fl��m��8!�ORh<y�L�P�<�b�d�`�d��C\�A����pB��4�=���A�82զą`���$�X��B䉢F]>�Y3{�e��F�=r(h���E1 @2�oIf?ٔ�>q�g�?,ڀ*v�8J��}h�DO�<�dJ6�=��Lx� :dh�o^d�<����(��!��	�xH*I����W�9!��I�~k8C��$!��)�E!
�_u�U7��B�ɏ�\8"�ر��@Ǔ?0�C�N�	��޼rL��A�$��B�I$2Yb8A�KJ�1c���F�{P�B䉔}f����ء_��#��
h��B�ɧ~��w��hD��4�=HĞB䉼!�� @,S xg���!&`��C�'a�N��)]#y蘌:%�@��C�I�1�H�R��0v�vH4	�<dlB�	gw\�ר��P�*0����`vB��B��1i�nO/
���/ҝ3EdB��D��ҵ���Y���
�x�C�	A$!h�"
@Q X�B�W.�8B�??x͚g�^�5��|�J�5d�B�	�r"mQ�UZ�0�eK�&F�B�	+U�Tٰ���	���H!FѢ.��C�,�V����ՃG�35Jl�B�)� ����M��	��ʕB���v"O��a�J �����LQ}�*)0"O��bON�K
��A
�m�r��&"O�<)�<y�2i��B

+��Y�W"O����ÂW� X�� y=�0�"OHQ�Ae�'��}� �/s�૒"OVPi]��:i��Y9�8��"O�1��NQ��� Rg�=�|�	�"O�*��ΐ�����H�Ӷ���"O$��e`��^�&�i%�@��AA"O�G" �!(`d�U��a�j@j�"O�l���$���9WIZ,S��z"OBu
���SL��p���C�"OBM�Ц��e��sGM=!����@"O��R��(*�t8�(� 6ӦP�D"O�-��F)n\<�m�s�z���"O����O�x�����.��͋�"Oj�ˡ
ÖO�j0�נ(�\!
G"Ol�ڗ�Կo#\� p��2ܘ��"O�(�b
�i˨Ec�_� �"O�|j���s�Ρ����$_ r�c�"Oڱ��X�d�VQ2��F��"O����B/O(�c���@��C"Oؼ�ᄗ�3�H=9�&IG�
���"O*��I-5� Kʏ?Ѵ�@"O�@jr,�!Y1�QCv���ҘM`U"O��U��z��W���B��:c"O��R��H<,�$�ڴn�x ��"O z5O�|���c.�z堅
E"O�ّL��)k�	�k2�z&"O��YS$N�S�293�̕�mJ��
D"O����.� \�dٛ���V�]�5"OP��F�ET����P� �x��"O��T�t_d�x`��9�nU�"O��PcHOJI�L��-
p��A�a"O�����]�~ь��/U�1�����"O�̩���N����-K��Q%"O�`W#��y�pHc���=��"O0�*���GI���«��e��Y�V"O��g,2>��A��G�g�t-�u"O���s��4-0�d�I�IL|�"Or}���V���(���"���h�"O0k0���P���B�ԭ���"O�,�qGV�a(.dK��͕2e^�q"O�l����K�"�	R���ITFPsU"O��Thݢ:��!rɅG�Hz�"Ol� ��
V��ѻWI��c�
k�"O�	�@%P�cF�=�r�J5uV`�0"OT�i � <�+��ɻ^ZLJR"O�ea�"�ZeT�G�.�naA2"O@̢T��6� ��3%��Q��"O@���?x��(�d,�e�*uk�"O�,X&�����i��9���a"O�8����IH8L��h�1���D"O��r֭t�@A[��޴[��Z%"Oĥ�)�k��9��9
��¥"O�@h��$ߘX@�d :V� ��"Of�[uᆅ2���2�^�ntp+`"O�`J����l�^�s�F#s�$�k�"OV)�B �,g0�����*ġb"O,x�Q@<PV� �����J5"O�5
 �D�p�
�i�!0����"O�h+c��c�p��!���� 9"O��+�/��Q��%s�D�������"O� ���a'S�h��X�3b�@|Y�"O��1!��D��({S�Lo���0�"O<��CƏvl�\����S�R�"OL��f�7�.Ay4,؀	��M�4"On���
�'�f-�J�0�x��"OJ����D���J�)����E"OT���ʜ�Ǆ��)�_�N9����\�O�aS)��CK��;�ڲLӪEj�'��Ce�Db�b;;�"HӍ{��)���_� ���#�aRJ$���W�Z�!�d�U�� D�
�=G�)s�
~�!�2�Е����w6a��f�&+�!�$�&W��p��l#`)� #ʃE�!�%tpB�k�`	(s�Q:#�@+F!��^�~�s��|Ҥ"e/T�w�!��+vi��.P�	m�PR. �!�d�8J0@�@N��N9���E<h�!�D2Eĵ9��#$�)[�%x�!��1y��@�T��.e�A�A7^�!�4
K5B�$���� i�e[�'�(5-}^���b���l`(HPN[P�<�0�1�:C$>P��hY���L�<ْ�ACᶥV$�!��)�D��G�<�w�Me�5J���N�F��H�'M�x�-)F0�啂0̃���0�y���;^(���@Ȗ,wJ�T�c�Z��y�$��5���o����(�y"�='�uIw�N�m�����d���yB�\)%Қp���X�`�]�GiT��y�o��l!)��Y'ef8�j�C_��y�b
O�2���.Ͻ*�|�z��T+�yř
M��)�$&J2 ��!)����'�a{R@I�?RH�ӠAU(�������y�K�O�z�!��[hg
4�BI��yb��+7�BU�d�g��������y�-��:�3C��5\��m&�yRiZ�o���I�ԓM��#���y���J�pKc�ԛ����FC��yR=Pu��(�&L�,��JU�P\�<I"+E�+�����O�>l����&�c�<	�ۘU���:92��vʅt�<�E�O�7^�1U� ;Oɪ$H�Et�<���$�јG+�-k:z�S�MT�<a6oQ���S�-�.H�3��j�<�3��`��*d�˶1�(%{vO�d�<�`/9mq�͈���18-����J�G�<1�*��a��q�����؉bd�T[~��)�'L� ��2��q$�	��%�;t��[Q�1閯US��ܕh�`��ȓ<�P�	�˙P��j E���݅ȓL@8�U�X/R7�`���nx�ȓs����"��7c�j4�FS�8�~���_����e�A2P]I���)
W�y��W���ٵgo� q��yv=�ȓD����F&��)�lH����Y!��ȓC����/Ń:� ( �> �04Gz��'I�dC7G�6�8�'�J�d�
5��'G���b���� Jf�%%E<M`�'�f�Z��:��4� D
0N~��`�����,B;B��E�.t�}�ȓx��]���&c,��q�'>�Z��ȓ�<�������'�� 8�bɇȓ_lH 1��؍;�jT�QAV�*�VX��@<9
t�Ҿ�!��J�ΰ��S�? Δ	r�Q�7���.E�x�QAP"O�	�S�@t��$m�,O%���"O I �iR�_�jt���ˋ(	|���"O���Q*�0BZ8�C"`[�D��"O��3 ٤A �!!&��]��I�"O~hz`�Z!�4ˀ�^���[U"Ot�"wτ�y���Aʐ�` ���0"OR����=/!�MkèB�/�|�"OD��%lEG �#�Ɠ�A���`t"O8�	�F�#q�"�^�k}�bs"O���e�� �.H�6�ـ5�d�y"OTL�"E��"W�)Ĉ�&x(�"Ob�P���9Rܡ������"O����J�7�J` ��Ϳ`���+"O60` ��i��Yz@׻f�d�"O�D�Q�Sn2�a��x��y��"O�A��k��y�ڌI$��N�T%c"O����G/<g�]��ؼ~�uaR"O�c�l�q�F�Θ�/u��+E"O��
׏'z�V�Q��Tn
P"O���G��r8r5p��;bd`�"O�xڠK^��a�p�ņIf�\y�"O����K��N�9���BO�"O8Y͒���s6g);�m�"O���#ݜ	���W�[�K2���"O�2r�V w�	�#��E!&�""O��ɄC� l������h��`���;\O0f��?[e�����2�~���'d�L5�!�,h���0դH�2�P�ȓc[����;�2 ��5&z(��IT�'P�x��8sE�A�d�L-޶���'�@�i̄YO��˴�	.O����$9�S�4d� Y��MU/B&:�0�݊�yR�H�
ҘU�d(S�"����Gғ�HO��=�OÊl��9% �j�D;N�0�
��	)F�4��FQ96'�X8�GQ!|P!�$�,w��(�1�G�-p���*:!�$S)MQ���O ��Apń�#!�䘮Kbl���M���	۶U	!�d�3F�X�
0���{!���C�Z�}�!��_���@+E(�����2�Z	�'>�|�H��)���>A'D�7O
/�y��#̆�)-.\Fإ	���6�O�+4À�)������ON�r�"O>H�CR�6�p�i���#;�|�"O�Hyde^%.|�r��� $��)ң"O�л��֖VXɣ���Pd-��"O�j�e��Yj���ğ�T�P "O"u13�Z<]D��17��0?�=:�"O����l	TQ��՚|�L	�"O����D�Rug����=S�"O��!��+����v�'�4���"O�����Y�> Z�T�- 8����"O�U���ո#�AB��h,�0�5"O~��Y1X�I�I�1R�B��4^�<!��@'lr�D�7R6Da �XU�V\�<1p�spĸ��{�4�'��s�<Y�ᆒ-���H�̙;��}JI�D�<����	>9��>`�����ZA�<I�H�,l�a���@"<p�N{�<U�oOƘX��Q:C}�AQ���R�<!2a�e�0e[���7M�^����\P�<a%$__3�=[㢃-?``����u�<�c&��X�
T���13�8�(�}�<� "��@J�d�<��F�2�d�I"OH�)v��;��)��@Y��"Or��Q��&�90��t�G"O�����M)G� Q�詪�"O2LZ#l��=r2��K�	z�����"O�Yo�>�"��䗌ax�H�6"OPԉso��/B�q�1䛀l0 �"O+�!FR��e#�'o[>�ps"O��hj��.o�tpa��Sd]B3"O �
�������v�o�|�"O�LAAM|�`�0���:=�4D�"O��	�B�"J-
ŃakY�h{*H��"On-�1)�3�f���)ӆ(����5"O�<K1��LC�͋f5=����"O�к$��o��D!��J�mt�Ӈ"O:�́�,���tJм7e0 ��"OD��ƟSed�ʳ��?��a7"OL���CƦm(�b��X)@��9"O�A3�KRi���tF�1O��\��"O� �f�
"m3~@ F��>q����"Ob�$��f
|}hXI¬b+�i�<	5' �&��=�e̞�XO0@+��k�<�7�8yxб�b����q� j�<�e��R��Y�.:7j�:g��b�<�&L�_'���4�H(�lt��Mx�<!q��4)�� tE�&y)��kW	Tp�<!�*��[�*�@'�O�z]l[�i�<�S-N��Z�Z�cUI��lS3�l�<� X�NTd�Āx��Ȅ�R�<�4(EM ��h⌍�%�֤����u�<�恟�_4�p�я`��]B�+Z�<II~�(F�.�bu:D�~�<(�!�"�(̏+�h��@GR�<�i\$��\Qdɮ1��NN�<�#_��ԕჁٻ��Ѧ�t�<�s*N�*��mH����iZa��Ur�<p-֢9�@%
�׎y�Ԝc���p�<A�eԄ?�� �gϦ3���hk�<���"ޠ�0��./&�1�Mh�<Eɓmf0�h#�P������b�<q��M��"��Q�Y$�Q1�^�<aR�<�ػs�� �Ɲ�@A�p�<	B�_nHYgCŃx��(� bCU�<!��/Z9���ـJ��1��*�Q�<����
�v4}�dhG�UT�<IC�X�Z�L��*˱Hc��!#H�<q6�E>��H8 ��)��X"CQ�<	��f1�s�N��@���� R�<�Q�� VH�6RW^�����d�<����(�z|#r�üYh��U-�w�<�g����ؕ/ 3l��y���
H�<90���Z�ls�n�'!&>l`R��Z�<yVʖ�*eĉ)�~��4`�'L^�<q���/�����H�?-le�#B�b�<��K�6l=���N�7z�a+T��U�<Yb$Z2k� ��!(]�72���W�<	� M̾��p��2���!��M�<��ϕ�=f��ǌ/?�( r�I�<�e�
1U�-��N
�I-4��%E�<9�@��1`c/�&L#(㓁 z�<�!�O�5���)P��J�.���h�r�<	Wnܺ;_, G��q%���#-�r�<I5nC=A�%�����):������k�<i�e� ��`��щ40a'�@�<� ����
��C3��g�G�Z��=B�"O���uB�85���S��׼y�2��w"O!96K� on8�"�ۦ3{�b"O �8B��t2ꅤykf5 %"O��珇;WD��،4W�y�g"O ��l�q����-����b�"O�إ�S��L�Q�X1�4k�"O ��&�>V��a��
�vOH
d"O�P�j��h}�E�<4Tz@"O4P��@�C����N�K,�0d"O�Ŭ4PHJ`�#���d�ِ7"O����������ʎ�Z��V"O$<B�b0X)�	�8=���2"O�쐱(Q#S+�͠ B�O<vt��"O81�*@��VYH&���I&dq�"O��Rk��G��� ��@��e"Ob��N,�&]i�xBb��"O��s "$dK`Lڳ �R�Ip�"O�pr6*�>oR(9� ��ҍx�"OB��f�ǂenФH0����M��"Oy!�,&���L�%��<�"O�I'd�8�fhኻd*x�"O��8��	�T��I�6�.-�"O�3�T*l�LT񠬄�N�4%�"O@|��N�*j|u@J�}d�	�'��Ę��ո_�P�Ë�a��
�'�Ph2d��3[V���BT<+ߴ�9	�'pl�y���"�\�Х��.*Z���'�(��/ҪjVZ���i ��R���'b�	�g��8E����lD��'�z!a��@-[�l���'�rA3�'�!��D�F�|<IUW�����'�氻%��0��D� ��z���'�h� M�\�@�D�^oR���'
h���A����ƭ�"S8��'Y�Xa���-&
Ԉa'��NI8d��'jd<Ѐ��"�ER+��G% ��'��Ń"�W%?�"I'/� U�@�z�'��س'RS��V�I$�M��'��8&��KHZ0O�$AY�E��'a@Ѓ\���)ZGJ�"8��Ț�'ς ��/H
f�6��irQJ�'/>����9O�����ظYv���'�>��p-R,Y�.�Ӑ�E!]�b(p	�'���N� 0V��6�
�Y�V�r	�'�.���&H�g�nI���0R�B���'���	%�6_�,1���VE�u��'�"�б��/�~�+� 	3f�$
�'%4h4��B
13WI�%P%��'���G !^1�C�!In*�Q�'�"�b�,s:�Bv�B�A�x@��'��'��uk���`�ڜ5���!�'3���c�"kd�LhW��-�|Mk�'5����Ŕk%�q�Nʊy�z<��'���J���Rh]ڰ���r�PP�',�y2ש� ���r�'@�p� �'^�����(� ]Y�*�M�����'@���$��3� �e�;Bo8t�'��jׅ��C���U� ���%�'\���1�����z��ع-E���']�1Bs&K0�	є��/t�e��'e�hz���6^d�ӌE3&�ٛ�'L�]A'��LݸV�
Ј�'�԰��(�1*E M���5~DH���� "="���f�~�E\*	����4"OH�I�%F�R�!�>G��:�"Ȏ��X�B�*�I��Ӗl<a"O�@�D�s��!�ED C�`eI�"O(��%o/\Y��k��U/ �r��"O�5{�ˮ,���	"#�7�h)�"O��0��%�܁*0HZ����"O~U�Pf�<p$���g۸&��M�q"O��#4� 0R������&�`3@"O� #��ߠ]�rl�Ҋ�<Q2�$"OZ)�ˎ-P��a� �~� ��"O��*���(�vU�7�ƧEb�h�"O&E��(�:��;U�E�i��"OD����4��¥�ǆ<"<��"O�L+G	���+ж\�D�Q�"Op(j�.�,�Y��;Pր`Hq"O���&�W*)c剧I݀a���q"O�u�4yl}h�j��W�D��"Op���H�j~fu��A=sD+"O�0���Vnf��	<CFx��W"O���`ë0/^h�b��+<	<	��"O�����7��*g��
��0#"OR9C1��7me|���oO>A�"O���3D�bХ�s���	E�E"O���F�R�>��=ÑmA�j��Q�"O8QpA�W��iR��="j�� �"O���`�6j�d���5Nn	��"O���W p��%N@1H-� R��E{���~ԉ3H3+תՋ0�#Ly!�d02���Fŕ��V ��ai!�ɘc^�M�Ů�(Oά-ڂOZ�}u!�$�^���pA??Ѣ����`!�$��^�Z@�+KϠ���^�Y/!�FMἼ���	Ġ�JZ�N!��a�r�%��0�d�I�8~�!��Z�"PA���Y��A
��֛�!��r��Ȳa/;ll�Bg'��)��	X��D��m�?���	8~t��#`�:D�\�N��q����l'(��4�R,;D�����F&fd$ ��n ;�ڭ�e�&�O"��1��H0� L�"��I�@	��I{B��t�p�P֪�P�`�h��� 4B�ɼu�$�d�W��`AB"
�-�B䉾��]3.�<,~vS�*��{w�C��>/6"�⡊���I	��-'�C�IK��Q�kW!*i���QM�|�B�ɜU&]��Ȇ?�(M���2�XB�ɢ)���q�_� ����!^`�C�	����Vd�7%
��ݱL,&����ɥS�上�lZ)]m�	�&g�{���d7�}��L�e�_"s�J@[��Z�t}��5n�X���X�_�F��C��"P��ȓ�~��/�F�.��Q�"H�R��ȓd����-vG�`r�ŝg����G^�(TN�j�^m���"~��� ?�	��c�Np����A��̣t��T�<�H���,��!H�Sb��j�<���	�a�d����r�~%:�)�A�<�B��2W��,"��H��f�t�<B� gX<�D*Ӏ@�4�E��I�<�Fn��/"�IVL� f��%����<��	&K�J�ڄ!� ��l��Kbx���'��Y5�^�h����<�TT���Ib�D���-qe.�`"!۫����A�:D�� ����ݖ<��2S펃-�\X	G��2LO|zg/�}fx�Z��ն�r���"O�A)௉G-zqSs�g��l�"O��Uᇟj��3$K���8�S�"OZйń�4i/r�x� H��8��|"��,�'�� �u!	�P6�b��I����M��6� ����a� ��ȓ^^=���͎W�
,	�ʞ�APB��'Ra~�a��R����� [4I����y��BPz�aBT��|�|��/���yRe��>py�Q�)�~$
ů�8�y��B1���"$�	�$��1�q闟�y���5�r��	#PZ�I�h:�y��
8�$X�F*�@%Hs.���=a�yRL����,!���)����D�4�?a���SJ#pظ#�T�h�dIX��,V����O�mI�Y8J�B����/Z��y��%�<�g�]�kG8�قEE�d�����JT�1O�{�jQq�aK�]�̄�&N�����O�|�"���Q1���A<5�;u�}B��[�&i�ܑ�&�|�<�A��1*�������<0#b,z�<�R�
@��ըW7���*�l�[�<�s/��F�$K=h4f8���~�<9����)��MZ�0X�=h��O�<�Љ2yp�����5s�M�T�IM�<Aw UaZQ�3KN�NN����M�<b��
�L|�Dυg�����DOH�<1�=X�zm�5k\�	����(�F�	E���O�(�� �	�"�r�7LV��'[��!1Ç+q/Ti���Dz����'~ԩ��
���mS�?,f-	�'t�\tBS�4c�}���ʆl�p{I>9���	����]1d^�z,�Hz!mI�E!�$�&4�M�El�WC|��Ն7I*�'qa|�HO$�� pꜱ?\�������'#��'0?�x�$(>q�y!�B�XҒ�9u)3D��S�Z�5Ś��t��%�pL2D������=p5l��b��>����D1D�Ȩ���[�Ɲ�)[;dV�H���"D�,p0
o���A�>:l�̠�M>���d.�'/�P[f�¶U<�;�H,�F���.�4���'�g��J΄Z"��ȓ��"�`Q/��jg�4����h����8L�
 �O�r�ƥ��H��u:��u,�%A`O�YbP|�� �����O  I����
���FR�S�RR�bK�+�R�S���>T�B㉶eO��!�e�S!�sc�'���F��S4w�x�� .V�a�ᘳ	�f��C�	�t4#�핌>G��6ɗ0j6C�I_�j�:A��4X�"Q+��ֹ!�C�I�24���؆�D�c�eU"*�B�	 wAlT#M�s��q�œ0��?!��iŒ[��0��H?}�%K;e!�$G�r�)�� A�A�u�ӏS�"2!�D�$sF��@ˏ[�"����q�!��ޓ��Yq �nt����!�d�Z�r@�㔂!�	sVS�Pt!�	\��x�Of���feW!�䁌7erh�c��t�~m ����!�B�fsJ��F�
�t� ؖ�Qm!�ě�p
Ɖs�.��4hu�̏B��O����|z�@�<HNJ "J7�d���c�<� ��2��H�"pf����H-���J"O�0���m}&�x���b���#A"O60�"��,�� �@I�X��'|,�@��l�|`a���{�p�
�'�
Պ�mJ-,G�!"�� �eL<=2���'��p�.ĲP���bc�ҕ����)��H׹*[\0"�\B��4-J����O��Ex$H="��a��B�	��*R
ţ�y�@J
%A<$�����5�����y�"��<���OV�qF��@ l��y�`��gF�h>��2�+ �yRFQ�[��$甏k7�<.4 ��'�@	�b֠M�dY9��:ig����'�ܑA(�����s�"D\i�`!�'�9�/N��H�C5M��h;p}��'2�,A��m�L��,>a��}j�'��u�DA�iv��i��^�Z�Z�'�:��5ǖ&��- �Z$������O�"|��	�I���Z��`IFr�<��E̝ �\a�D�	M�mst  q�<Y�Ɓ�r����TF�7�(H3�In�<�Ag�8���`���2&d�bDHDk�<�o�(m������s˔�q���R�<�2��B"Ȋ��ń]�~!�p͝Q��d̓��Lq�
A u����ϓ]��=�� ���I�,Y.v����uӥچd�ȓi�@	ꁣS�kN�<�&�١cw]��If~�Z�0�-�pE�;$���!M��y����dÖn�Zt��LR�G>�I�'Hp��!��.�3h�=�j�	�'J�dy�MN?/`T	@�_���#�'w@�J���=�b�9��P�E�.����x���+� �C��.�z�+�F���ybk�"-b�V)�$�T`��c��hO
��DP>9��C����&�.���Q�T���h���0uڵ@Iȁ�άq����=D�L���u6�A�!�]���R!�<D���%"�1z��-�N�;k�
ǌ:D�dJ�$ٿqnji%f�$vHL��E�O��=E��l.vH��K��6�=��+�y�!�$�tH0�7b�=��ՀE뗎�!�$Q9I'�,�1�'7Y������'3!�$U	kW�=�&��=&W�L��%�f!�G�;t� ���O]0��!���
8��e��
=�T���g��\�!�$>0����xͬ�b��YA�y��'�1O�,�䔨sm2䑰��LD�(`"Op5�� ݾ2�9�� ;�Hrt�'�ɧ+�3�$�"���Vb�=��1��OMy�@SN@�����]4��"O����G�\�u�<IV�� "Oz}�օΜw ٪G��>������w>��#��0^l��#B��M�ȹ1�1��?��	O:C$� ���vo:�(�,��Y�!��X��ႁ�̴��*0I0a~!�$�';$�Xs@�΋Q�>�Z�'Ң(��O� ���-�HI���0Qg��Y"O�X���׺P��)� ���[
a3"O���I��RR�D!Oa���"O���F#�5$�]0w%�@^6���"O�M�Ǧҏ[���
�EI6v�Q*�"Oz��`��vؾ�k�j���t��"O\i�3�?N��l��ő�@8��"O,��3@M5pgTp1Q�0/S��y
� 0!��1p�P8S���"�~e��"O�R�ovR@�`�D}Nr��"O��DJ[�}�b ��>�tT�e�'x���BG	m�Q��)�H%���*D������1Ai�l0��W�\dj��(D��bi͢@Yʝj �ٔK>�C#%D���vhJ1L��R�����^;�8D�H��a�~��`j���!	9Vp��k5D��f�J8M��1��	39N��.D�X��嘞3FDpz��L�4�4tʓ�>���?y����Q�\�
]HX��b"�>P!�ā�y�E�F-\
?*��h0Gُq2!�;hВ�Qn�]��Q6��$!������Ń	w	���D��!�d��}��=�F��Q �P�bC={�!��]�z�Dc)��͆�R,��'�6��B �zjrIB�NGZ�Ty�'�����L�?.~�ԹR��R��!��'�Z92�!JB��!LA/W� ���'H����_&�b�K��P���
�'bD��h�-���� �U��u�
�'�fthb߉J�];�D�Mf�i
�'��i�7�F�a�^L����5�l��	�'E�d��% jʒ�י6�&`	���'�� &��2}/�L�'b	e�<i�/tG,�{�͘�p@ÖK�<qpȏ�O���Y>5����w�QH�<E`LN��)�"�8t���EaO�<9�l��;
��{�lC�5�ś!m�N�<iQJ�";榙��[���ۢˆ՟�G{��IQ�$�\Z�B[�E4Z�b���b5��,�S�OC�E�禔�e��1J�H{٤�i�"O|�s�61O����W.9�$:��'b��'T�a@�B+x��)�4K:#Z��D1�S�O��a��D�&e Y�բӬ&����"O��Q�@�<QJ�ؐoE/!<�89�"O(���n)�\�*H	�D,!�#"O�y��7*�^q ��B]
LY��'�!��yZUJV�ڪ7Ȏ�JY48��'�ܴ�E՟i�4�j�a��1�' čóۺ/Db��),ˎHy�'�\�:#EXR��R�a��v<XA�'Q����S�9��AWI�s�����'hJ�e�7 �u(��� �v��
�'�jlk�b	>&P҇hH�t߆�P
�'�F,(�����b�Y�ky�D��'i �0ڃT1���F&�Rq
9����hO?�@,	�&r��X5���}:�Lc�<�NU'��˒j]v_�*�,Uv�<�f���o�Ƒ+5��d�Q�O�v�<)):��@�������1V��Z�<�T�8�����+zNTu��YW�<���D+<����B�o��}+��L�<�m�w�x��	P�J�U���P�'a����P"d��F�֡V�ڭ�5�A;��D=�S�OL���̽/�ڬ!�㊐WC*�(	�'Nl��!W	@ r-9�+s�9��'�fu2��M�8.d��v��%ll���'{�<#u�@;	��=CQJ����Z�'5��y���r�ꭈ�֢�Pk�'�<لa�u%���� '\����'��)q�ڗ\�2A��� |+����'�`̣VF%zPJ]9s'�}�"��'���2�n��	�h�iK�Y8
��� t�J��=]w$��e��X梨�W�'31O��cweB��VQ�2O8h�*TR"O 1J�� �`@��[��m�<"OpY�U�R,��1�g��%�©·"Oe��%�#;�P`*J�n�1R!"OB�y@�Y�֭a2��u%�"O~=�F'H5A ����Q�"O� kTˏ�1����4���r"O�s�*׆N�P�q0!�������"O�t���L�@�>u�$Ixe"O��ap͐<��[�Fϴj�9�"O����Y	I���jF�ұfOxy�P�\��Iov� YfKF@����Q,�C�	
z�A��L��$HIi�zl�C�	�q�$���O�7P��� �G+
���D~��iv��8g��@	
A�B�2�3D��S���3�Tt���-��sd2D�k�%�x�|���E���u�n�O,�=E���:M.(@��<��Y��m�i!��2	b�K�e�F�����E!���"p���� ��I{� s��A��!�ʶ��8	�Y:BʜC�,�P?!�$��r�T53!"O=S��1'-�8,!��X���Aǝ�$)VK@�m!�d�1V́�LہD�v!GI�7j�Iw��(������}����F"�M��DR�|��)��::2� t&̍W��)��6��B�<G�r�1�G�5s��p����/]fB�	BVx�񔅙�(�9�`��M����:�	1`>�*�,Xdy !�j�1Q!,C�I�ߒA�5LԊMe��2cΟ7$��B�ɒR����1ŗ:=�}J�A�8�B�(`a� �B���z:��	���?wVB�	-6��3Qj�'r�p 
U�vB�	�h� a	� ,:���3�b�wHB䉋Z� u �)�LL���4}6�=��� �\�"�ُtt(�Ӧ
�fP,B��$�6�{#�SzJHW�HH�B�I2$�Ŧ��7#:8��@F�A`�?)���ǔ[h�h��A����ۭJ�!�70�Y�cR3 &bC�H�!�©H|��7�+K�A9�/گvl!��,B���i��{�����ޮ4��2=O��b�._2��%��V�Q�"O���/Gv@�7�
�D�v�r"O"�EOƩ(�����:l� y�"O:��ǉn�Μx��ҧ%��2���|�rA�I�%������ضK��9z4�'D� �fJ
�_��C�-˲f ���2D�H
��'NkF���N�{��iB1D��"2G�x���Qစ$Bf1�$�-D��Lߍ@�x�i!l_	P�|�F�6D�� ���1�bqA� ~J勓�6D�L��߮{��YY�.�E- ���O?D� �����x�bvl�1E��� ��"D��@����x�HQ*�+R*8d\��?D��Z���DJx��E:�`��u�!4� S�&��I�!��b��k�#�G�<y��Ь,q6�S�iv�m�Q'�@�<A�-�aj`1x7�ݿ�����|�<����h��+��:�Ľp(B|�<Yu'Ew�����J�*�釫Q|�<ɳ�ɂq ʸ"R��1*%xbO�@�<� �ً94�"�%�#>*�C�O\z�<� �������yQ.�1a�l�#@"O��rD*	�C�}2m+鎅"O�|���!OF�|�3��v���B�"OJ�`�JW� ސ��C�&ӊd� "O������H��[0�˙?2�)� "OJ�Yr�C�CJys�'Y,l	��"O��sv@�>[8��g܃}(�TJ��'z�IX~2�K!D��@Dǚ�6(ܥІ���y	A/Q�$u�F��+�BUi����yrI�.��!�OJ%O�M������<9��d	�21BDQ�&8�M���B�|�!��FH2�I�Oѹ3�(�Q��Y.!��s��y+�N�+���K���/!�0U�P P�y�*��C08�!���M[�C��Ϩ`g�к ��'�ў�>�w�'�n)b�l���-�4�>D���Em�9Z��I��"� !S\��H D��[���'6��X6CK;���g<D������}���[�a�/w��5��F9D�ĺw(E�_��3׊P7l�|<VC䉖J��|rѣ�/���o)z> B�	Ӣ�r�X�Q��tCWM�2$��C��I�k�ۧ_�����Nҵ��C�(Y��!ZR,�/���IT��D�C䉲qf	�P�m�:�KՊ<Rk�C䉏N-���*Q�|g2M�����Y�C�I%�\�C%��!���aaiO�v�fC�	�V�f��҂���ʉ-p�b��d0�I :A�HY�h�8/�4s�K��,C�I-l�a��B�J��<��gO&`C�9s5f� '-C��s�BΚ]�NC�I�?�tHs�o�rJձ��+��B�	�%����AC$5Z�V�%pB�,3�.��5	٘h<�h	q� %لB䉅W'Zp��H�r�zĈ�k8S��x��H���4+,*>e�f�65���JB����0>q0�-h\��BHI]R�!�VQ�<�G���\���R�_�@�`aC\u�<	 �!('�@a^�vd�V�o�<�a�R<љ#�XlډG��j�<��*kD����X8؅Q��M�<)G�Y�<��xh�%��J)pQ����I�<�%J݇�b�U��>�r|���G�<IU擫�<�)��"{D�Rc��z�<�֧�!��Y���Č+�6e�T)Pu�<������`#@�Ҟ{���Eo�m�<9ө�5a�8�cU�rA�tC]A�<b�اݔ��v��5@�����R�<!�)�R��B�je2�����d�<���V�_���W ��q�,��e*]�<I'MJ�ivh�w#K2hL����Y�<�#�R䤁�gOdk�"*��B�ɨcn��1���8Nu�4��3PC�0���Vˁ O"|�R�Ɨ�5�$C��3l
>�i�.c�r8h�&�7-6�B�	��Pt���\�  ��%߬b�"B� Ymzْ�B=Q`'�.^�HB�I�t-@u���" �Q����E�DB�ɘ4Q>�z�-��?� ��S�G�cXB�Id� �˷�uŅJ�̜==fiQ�'�4��q�0#��h���~�J���'T�c�I�d���Q��9�b�a�'DQ��j����n	����'� l��C�@�D�zG����i���� <�҇�֊@4Y���M�fܚ""Or�r⢞1�h���w��AX "O���A�`+N��莆"����|B�'�Q�!��m��a(vg�	0.�p��'o�T��̂��@�T+P����'��X���h�8�b�̖�N��83�'�|[�b���ʀ�PfUJ�i��'�f�+ub�
N��ۄ	�Hs�%�	�'~�,Ɩ=Sv��N٦.��+	�'�I�6A !��4��?�xZ�'�8$�oǨ�5�t�X��L���'B�|��Y.)��y�UCY�L��c�'_�m����.���6��3��d�'O�؊w$)v�<8��Η*�0�[
�'�6����ˉZ�x)���L�|��'c>1!f&��D7������栓�'L��P������4	��(R>1p�'��51"�8]f�#��	vq����'��5�' �q�h�`3�J�d���R�'q>� kJ<���SIA�^L�P��'J�t���֌����g�X$�'G�a��I0�5�d)��I���j�'p�*��E�ZTD����Vz��(�';(��)�'�����ʘU)|�����+O�M��
^�z~���cT��r�)�"Ob�K���70�$�S�!{�)e"O�
4�ە4.��`M� ���b�"OR5 �kW!u�a��L�iwI��"O���TlI�z�ڸj��FLwL@T"O��1�kV�iCH|8#�
�#�"O�����K�~��р���:v
�2"O~\ځm@�'��)+D�}��<��"O��Be۟}jh�"dD=Ab�Qa"O�m��͇92C��-���b"O��c�u
n	��ŭs���I"O�)Sp,�x��<��gD���"Or��`�r�Fix[��eH�.���y�[�L2����&I+��A�@��hO����&k������V\ݪ����c!򄃳�)�&�G���4%Þq!�$�H�����K�.k��c�X�!�D��?`P��f &U�M���ŋ}�!�
�[��I�t)��>D(tR%CH�*�����(c4��Q�ـm���{VB	��y2Щ�n�;�.ЈR4�h����'�az�)�>M��@p M�9���@��X��yB�Q&V]b�9��ڗ4���B#[��y2�	49�x��B�(�:`�Ò	�y��[�x�ʸSu�P�*8�02�$�1�y�[�H�\0$�!nB���(��'Wazb�
�K�D쉗͔����q��y"��Rꨕa�I��/R,��]��y��+2��<3�@�6ቐ����y�ƅ�dhXg��7s*�@����y����N��Gǅ�-:�������y2��1Nb��J��%F�uZ�A]�<��'�Te(Vf�2�b�[��e$�@�/O|������`BA�	t��"��H-(�!��;2��A���G��Dx` /�5~�!�$QE�����Z�+u�1sm�;:!���X���$ .�⥢Q�
�!�!�d��A]� �ʈQƸ���D�i�!��(��ҭ@D�~���L�!�$��DC�X�F@���u2F�/�!�� d)����
i�@�a��!7n�� 4"OբDKE%F�n���E;Vh8�H�"OF�	e�7; �[�L:�=;T"O��KQ̓�jHS.ϕU-k5"O�cS
�/0�!����@�(3�"O
E�gKV�L�r6-Սh�<t "O��I�#I�+� �X�B̵\��r"OjАce/'�i5B�4CM��e"O���,�6/â�S��X3�Li�S�������CI4P��2 ݑh��B�ɦ.̈́��bJ�?��9���9�B�IxX̪b*ƻqs�ա�L�J7�B�ɎC��gK	
C��Ě�Ĉ�`��B�I�T/���Qi�g�h@�.��tB�	�*&���G��<t���k���<B�	:�6T�Ћ�"I]�Y�6R�R�B䉟O �d�'(]�n�#�71B�I'G��P�-��D�V�
�j�o��C��:/���Ȁ�8��m���9��˓�hOQ>!��E�۰dpL]>�^��Ai;��S�� �C�ύm� y��[$���@e-8D��{4'Օ�F����7J����F:D���7��-�������0a���o3D��6+��)�8�����(R^x��R'2D�4�@-ֻ$��"�.ū��ӈ2D�,�����3�y�*�9Vp@�'3D�R���@ca�Z
Q	@}�S'D�|���ޡ1J�->v�:�� @9D�lZ�l�)���3aI�"*�I�7-<D�t�Q�R�cbTm)�U
K���A�;D��{fGL�A���	6*S�hD��rC�$D��I�-�(�؈e�O�],<�XFO#D�+p�9��9�(��
H|���!D�$��G.$�5Б執!�h��$3D� c'��P������E8�aT�+D�)�O�1+����}�*D�A�(D�X[��ǘ�LLʅ�U��H+:D�iel�._=z�!gO��]��h���4D���4)�Fq��{��1HƼ
�# T�\����,T{"T*O˓K8�u��'�ў"~BtC�+�R���A� ws�C�l$�y���X���F߸~��AZP���y���H��J�fH�A+�mB`��#�y�/��#!^(9��
.k��aMX��yB�]�h2��XW�Λ\��crK�/�y��#.Bz�0 �>Iz�Ѡ�Q��y��q�̰GD�+�h������y�FܷAjb��p��W�,�l��yB��GB�ٰ��W�},X{�	
��y	��$ �k�o�x��L!ţ �y"�Z3�H��U�p��!	��Ǚ�y��F�yf\����<a�.Q�s���y��A��X�!̆.�r���M%�y��"����֡ۡS)N�!쉃�y�!�o�d�� 9���bbc�/�yҏ��;� (rO���ɳQ*��yrJ��k�H������9���E��y2�W�B���w���d!� �yr!��C�fHaD	�;�
G �y"��8E��Q��҃�������=�y�]�v>j�����_< ��r �y"6S1!�dA�[m��q�EE+�yR��)�\��sfN�j���� LS)�y��ë#��<@���_�LiW�<�y
� ��Yb����4��)��)��|�e"Oi��ֆL>�0���8���"O�L��èyDH�'�!�(Ar"O��a�'ؙ#ڮqh�Ǚ�[_$R�F{��i�4w� ɐ �ָU��ArŌ3!��H=6\s7��_98i�A�s�!�d7J{��4��{���H��!�dՙT� B��ަ'~��h��nf!򄐃!������6�%XG'X�mS!�M�Fx@ds�ĕ8٪Ո4&Z5x7!򄒿Y5��$)ǘ|�.dd؀#5!�DL H�P�	�*��#$��Y�!�Z��ZD	{��9DC�!�$�D:�a��F�B�"��ǳ>�!�D˿+��Qk�)M3,A�T�И}�!��o9�$�cLɜUNdu���k�!򄕜�T�Ѧ��&����*U_!�d18$�\@5*W��4Xjb�6-O!�$A8!{��
e��[�V��ֈդ^�!��[�M� �W�. ���6'M�!��M_Ba�7'�\i��U(�!��.>� ��Ɇ\W\�2��x�!�Q��B42�NA�!"~�!�d�&Y׎����78xZ��ڇvf!�D�]��D��U�"	Q���$/!�76���F�Pw&T�7�U
!��;�$�HW�G;}\��r����!�D�7;���c	�,S4u;`(T*!��m/$��w�!H~e�$�ަ~!��8K�� yA�M1F�,dFL^�!�3F�A�!W�
r��spJ-5�!�䁥[}L��!�L���HE��(+�!�Hsi� H��W�ش�ul�>=W!�$+f	RmSP�W&������_�m�!��:�H�zc��B��8���GO9!�䒇(������ P��3�!�d��Y:�	���'y��8���'2�!��K�Iۘ���K�,p���� �B�@�!����հ�=�%6�P��!����� 
�%���(�K�>�!�D]�O��&G �J�V`�1�!�d�\"F�붏GG��y�2`�4*�!��1��y��I�+�"!p�NY!��-$��8��GnrlhD�<�!�:Rp��`1�ΓFm��Bׄ��4�!�ɀ;r�0X�OU�c�ĩ�VA�.bj!�dǣi�D]	Ao�7�t���L�5^!�߱\R8h 1�B�c��V!���K��y��剅0�*ٙ�A�OL!�����݃�j��+�6CG���!�R�P�LŀW�,��&E�!�d�>�17-
�<r ɘ%��t�!���C�	fE��VO�E �d��ig!�$,F4\R��
(J��ӗ�O�>^!��6P��mq���n5F�97>�!��G!m2�c��� �d`�1rA!�d_n|~�A��j�d�C����4!����*��N�Nm&eY�ɺ\�!�WE���
SΞ�%M�k�`I-L!���'��Qy�R����	{ !�D	$3W&� �K֣A��$��G���!�䄟LHS�ŇC�te�sL��v�!������t�prr�r%M���!��ڲu�f�d �KlFA;�L [�!�� ������%aޱSD�
�����"O����MH�gP��G�Ѥl���"R"OBUZ�!\F������S�?��ț5"O.�1e��X@�8x�׷mb��"O��YUÎ�#�N��FK��_W,��"O�,�	�"1gh�r�	�+e�@A�"O���)�_-�L���N?����"O���Cf�'��i9eH
9.�S2"O��&�H��~��F�c��P�"O����F@�R��9¦B2���B"O���1E<ntąӥ��ղ%"O>d�v�ݧ/�@<�v�E�'.�A�"O����W�=�(�1�熴 Xd��"O�8i�a�V}*WMJ�B��x3""O��3j_l� ��Eӈ.ؐ�SA"O&0�M؋Jv����Y�l�rb"O��1'�	QS~܂ň�;�N��"O����7_�b@��@G��P�"O�L�c���}���k�`-.���0"Oʹ�.�3k(ڠ��G�2�J�"O@<�Ah
�g�����>����w"O�"w/��QY\��-�+�̽�A"O�<#I��'f����Ӟ M��S"Ot�8%� 29쬉��ЙS��U��"O�T�Ӌ�V�� ��H�p=��"OPKc��,}���i�&�UZ
)�"O��#�څ4�9�3E(lG\u��"O�t�#��b�2%e�{�����"OJ�H��G�5�0�a�����"O,����0Ƀd"ͬH/t��S"O�}���ՐXn�:���\��u*O�H��kD�*r̻ ���`�'p�kqd\�����+6�4��	�'�
h��(
�fW a�!�[���	�'���Wd��f���W�=J�:	�'�F��'[�_N�LX��M�]�Y	�'f��0B��;��0j��۵Tݪ�i�'5�E�Z�y`\���F�5���
�'İ��ࡇ j�\�c(�5ΐ�8�'��{WZ x:��3��#�'e�;���Z� ��RQ���' �$C��:�EPGBԞC�d�@�'���q[����	!B`�%oYc�<�pNت�n5LO�Y?��!���`�<i�e['l���˱R|u���cO�]�<����F?h��N�Fx)��Z�<�c'�3�*�����+��]W�<��"��p�`v�ˋv�
���O�T�<1�&Ǐ0X��Fop�0��K�<aԨ�~h��󉍔F/$���jMK�<�U�T�&WZ�!Q@��B���[�<i�8��K�a� ̡����c�<Y�c��1:�g��p����"Ni�<y5EA�4�~% qk_S9Œ"H�I�<���K4�j�{!�/K�!���q�<1$Q-
M�'�V�#�ʬpLj�<�7��{�QL�-���X���l�<Y@��>�oˋQCD�3 ��B�!򤕓DrP�E,<%N�CQ.�$x!�䆹CrZ8�L��d��jk!�ă��%)EǒiT��sl�%pN!򄆎3���B��G�SL��A!�$4}����SmٿC<Z���.�!�dA(!rH�R^,��anW!�� f�y3�dVfi`􌖐w�>�P�"O�nQxd̒�ī	ΰ���"O�|y���	Z�!4�ɖ���"O<X�%K�%ISN�{g��.�2�s"O�hɒo˳c"pD��]'n��"OX�+B��k�ΠC�+��8�t�"OT�1Q���E���3��88�8�"O&��5hĹLul�r��貢"O�qI�鎜/�2Tj��@�j�ҩq�"On��(bt��oěw�T���"O�!q"��	n��#�G?t�$Š�"O���C,�XSV\{�ŭ3��=�D"O��ph��iB�-�U,��k�$h)"O�4�wș!Ke2���k:;����"O°Ƀ�U�2X,�r�@0qc2!3�"O�����ޑ&(�PM�9Z��c&"O68�C
�$�a�p,&�!�"O��3���
���P̆�N#� 6"O��Z��S�W� ؠ���#x%�q"O�{4�O�F#L,��, D�"O\@�̏�+S�1Y��64;��Y�"O	�!i �����ʕ&Uꅂ�"OJ�,[�c<6�S�ӉbBn��T"O�H@6mΡ]"41Jv.7�I�"OL��ޯ#��Xi�ꀌ](@y2"O�	�iհ<��Y�/�un�"O�0Z6`z���Xw���3"ObD8cO^-��J6C'�V��v"O�e���>�M��ـ?^<�E"O����)�c��1@�O�br=��"OT��ڼ2��ٰG��#k��}�"OaЗ㒕U��Q6L b� �8"ONEapf��!�����z���KF"Od��A��<'J,��Ζfz�j�*O|�0AB܋ ���pL�3)rxb
�'x<Dz3
*,Dm��a�D
)h�'r�򒏏Dt��;�����a��'����Kq���	�,O�O���)�'�|��d�:g�(�q��G���
�'юE�4�j��F�<VD�
�'o�1�.��H����ԇB��:	�'����쓄
�J�I�$8:c`���'c\8sO�Q�X!���4�ZMA�'��/۬G:�Q�-����'�Xz$�7/t��U��o5�	z�''�a���/ruJ���"Q
�')<J�L%QE�pa�d������'2vxcr�ىo�$�ݞ6�Y�
�'��ݡR�Ɛ @�Qs�gHZ~	{
�'�@p��x4=���
�En��
�'Rr���1DaZ���; *��
�'�Xy�dh�%!�L4`F 5}H@@R
�'KjI	D.0Zy��)�}�Vu�
�'������R���Q���q/�l	�'p����`D�:fe�D��S�T���'��Q�R`�$t-�4�@#R�4�x��'�Z)q�'%V�z���&ߟd���3�'�,���H�p��{W`�e��'p����!tM�]����c�4A1�'.l=� ���[v�
�ݞ[0���'��X@�ִ*\��B�S���C�'�|�6aM�$C�	u�<^�H`�'2ĩ�ҍ�nJƩ�d)OXҀ��'G0PSN�d�H�(�%>"�~�A	��� �-he�4��d�@OT��5"O@�����J.	�g �kCv�d"O �@���.~&�`���!LMȤ"O�	�E�B�<�q1��y9�"O�D�_<3Xv eQ��\�S"O@��T_�uV}b��5Ϛ�J"O��p4O� w6,���K�$XleR�"O���T_���BiJ�%`�؀v"O(d�/��q�ͲB�L@h�!%"OhYub�<$=@���D�X��"O���%oG2���!�-��"O�P�f�M �<�,�w1�=�"Od����:Rz�Mhg�U$X V��D�x��'z ��'c� �� =��X��d>����X��p�A�Q�����*?D�$��B2[�PR��Ά��i��x��F{��)#�,ͩ�KQ�B� 9�ՠ�?f!�7Knm8�h�>K�:���)M�-<�'��|2��F��B#�^7�f;�	���y3f�d��nʁr���D,�p<I��$W�k�DE+!��*)X�#Ɓ�8P�!��ڧ+�F\�p�E�5"=�MR�Q���hO񟢁YG�C��Ȧ�H�Ȕq3"O�HyvhΑ-�<���Ĺ���s"Oy�A�1>��j��y5��&O��1�,ōf#�Mr�jPac`0D�<��_8#{P7 Ň;��H�$WҦ�'t�܁����@u#x5�ɔ	��E��-,a{��$r�@H�@޺i�K4��B�Oڸ�牓PV���5��*��cp�O2�8C�I�r���&��o�di����kcb�'3a~©��7�p`��'�$�H�!�G��y��ݖ;��q�sKQ?$�(R�[��yҍ�f^l��		)#�F����p>qqɐv�VE��c_�V`(�Q �zX��Dy��>�PIb0�Բ�<�"o���';az�d4] |b�E�l��6�L��ē�hOq�"��$*	i���'� j_����(D�\p����hv^\s	�qW��c�d2D�x��ˬ4n��@4F��M9&`�=,O�,�'߉'j�1��g��PЋ�
}�$�K�'|��QG$�U� �A�A�`�pp��'H�D�C^��Qʣ��-d�50�'qb,2����p�f��cI�:Z.`��'6 Y��*+�u)bo��Ph.�b	�'�F�J%�B(�b�`�Ț{�D���'�B@��iʤ*7�@��C.���'����
���Ȁ ۠�\xu"O<� v��Kx���oD8.K!A�'�<+�_-pq�	9��ܜ�� �=D��y��X�� �R"�g,:E�7=?���ᓪ9gJ�y4��>�>���l��_�C�	�j�cʂ��8�6�2Th�=�ÓX�"\@��_cN�#1�ʸ1�݅ȓs4���sm� ����	7�dE����0 �M>zN���֮{���j���d�-R� A�F�$�.8��O2��ӏ*oAH-�7!�k�D�Y%��#�	R��ON�i.Xo�P��՟���D
Or6-�	93$m�1
Ƶd~xMC�׮"W�'-XqFy��?�$`F�8,�����Մ&��W��84�^��d�k�'7��"Sϟ�&Yh3#A�E������'r�u;��T.`���8b��#�
E��'�8����:�x*7T1C�l\j��n�L��|���� ��JQ��,a��mÓ)�|^����'���C�ĳvQ�(��L�1O�T��c�ODC���H1h�+�E�,�����I˙4�c��Gz�I��+��A;�mV��(`�m��h!�d�%�T��a�݅u�jq�7��I��'�j��	,'� �@��m%���4�S(3Q"�����M[���7U��Y�m�xr箌i�<ңB1\�(�e�<�B�qg�h�';?�;F����	S2KGm� ����3D��z�%�6r�\M��kуr����#�3��hO�S3\���p����r3���u�ݹTw^��%�L��4r aE�`>��gh�5
8��ȓ����U�)a��1!�#<@e�ąȓ^�xɳ5
�r,��`w�˾`��0�	s<q���(<R� .�<k�+n�,��y��	�-X�E v�P��l�R���P[�C�	�ECVH;Ta\�2���X�K^�B���O�=�}���O�y�`�nAy�&�����_�<�》(�AҍS�Iܮ9�׏�W�<A����T���@DFN3grH +Ć�VX�l�O��HP
?Q��ۥ��p�\x"O�Ȱ�9�%��K)gP:,��"O�9��ހi�|���	�B���"O"�;󋇶#C���&$�ٰ=O��=E�4�Wh��@��M>��A!�yb�Ix"���M�D-���L��y� �+@j)I�*��>�\��a#@+�y�"D�%�L���`�;I��y2DWO�8�1�#NX"2������y��N�G���2�ߴK�Q#�N��yb��5{ȝ�"!ٝrqه����hOq��l��j�
�xͪ"N�P�L�)�"O`H�������P��G���d"Oj��Ã�r����FH�U��0�c"O��(6a��&�Նm�<���"Ođ���g|�a ^���"OH��n�*}��EcNԕy��AҗP����	>�����,,�Arj��,b��G{Zw��9�N@*�χ?"���,?6K����i� � t �7�j�1��8��B�	Q�QR�g!]���c��%�B�I8"�Ja�Нv�2U���[�^BB䉰0X+�E�dd�K2��}�LC�I,W���pa�� �N)���p�B��?��e�́yN���猹֖��d-�L�q���
�m��~�Bg��]�!򤐚e:�����j�n`R&B!���E{ʟp�WAL�;������,0��M�"O���'c�kl(���U�9��u�"OqcA*��nA{�M[�{e�p��"O�Xz�i0h&�8sp�l!��Y7n!���=P<=#��*e�#׃J%>PQ�P�'�'U�Qu��nǴH���*$f<²���Oz�O^�/1f�H�&� p�L�xǚ�pF{��)�54Լ�Y2M0?�@bƉ��_���G{ʟ�u���	;���0��m޾
��9��4|O*�ӄ�A>S� 	s�Cb��Hz�
OVE#�Ś�U_p�A �&szN��b��y�#�ObƉ��$��j���0��y�-[ �´��L��(�g���y�KW�2����76h.��6�ن�y��̩o�!��ۗ ����.�?�yQԡ�`�(
���A��~��'��Yq׎]�K�3[4��#�OK��HODO� �Q��ڗp� �R�O�}Ծ��"O�9�j�0Xj�	�kݔ̖���"O$A����}I4�J �l�A�$"O���T$܃)�8��w
� fo�(r"Opu�C"U!
�^�C�f·�hC�"O��bFȷL��$HW�E .t��x�"O�uHE�3&�D��ĳ	M�1�W"O���4�ѫY�b���dI?(��eb"OV�z���;aVD�-�"�b��F"OhuK���egHWD3�NY:�#�k�<�ԭ�A��ت��S�\(�p�/s�!�d����c=.��k��F��!�șz((h���P�N�����T$!�ZUҪ�˱O���݃���:�!�DG�$� 5�񦕓b���cW�h!��>Ίɚ7�וMFPIa��[E!�DƌB�d�&�1*�,{5
�#r.!�dF�pt8�7�^�����.[%=*!���.W�]�A���r xfgPZ�!��B"FޢM2!�8{�*����+#2!���4i�f-Pyܔ��$��'�!��N�nPp�yb�]�w��x!"�<j!�:F	�<��%�;�4pAaJ;)A!�	�+!-N����	W�!���"i�vK_?VɜD�wĘ �!�䜯s�`��&�zi��O�<�!�]13��AFc�J���!Jt�!�$�%P�����oY���ꖀS�l�!�DD5>���P�5{�Y��,@��!�ܬb\$��O�ƨ�E:#}!��^����G_e��d�9P!�dҲ�{��7� �RbDne!���,%¦��<@�� L|!�]�B��EӃ��
#�x��D�~�!���M�pR�-��;�m�g-y�!򄒃gBE�5�ea��=_!�$�aδ�P۲;9���~E!��ڋ)̆��H��I�)JЊT/X!������@"�HPq��?�!��[.�>8��*ל7�T����6|!��w �uyэC�����&^�!���;��10�✼P��Q"�c�!�d��B!�Q�ָ="ԫř?s�!��9C�*�Ã݉O$!@��Z�!�$�5<+ԅ��(��q����8!�$]�Ɇ���yuX�Y�فhR!�d�|�ȡ��֟_m�U[���HN��gl�	?a~�A2F���P�G�-�h(�UT�y��U/:h��i�4.��у�U��yr��X�T�	�i�@�ˍ�y"È5Y��������1@�U��y��߉��i1��,[�@j�����yR���p�0yǏZ�	��r��A�ȓF�)�΄�>E�eH�mh}pl��{f.��I��A �!Pq��^[2!�ȓq���&�3f� MAgn�����ȓ`�ʩ���׎�(s��I��H�ȓi	~9��O�.�F�b�#5�V8�ȓ-��,�dD�:|N��"7Y��u�ȓZr����V�X�H@��^� �Jчȓ,u�=Y�� 8�(��U�c�z��ȓ�e[G�$�����٘�\���

��7�I�d$�;gjښ5�B,��5u�����/n�IA��]�^���S�? �@�BEVeh�P��\?��"OxBr�Ќ+4h���>$@�"O���D�ي$ќ��aB-D'DdKc"O�EICm��X	|�C�Jf�p"OD���1^&�����2i2s"O8��u��7BT����ƪh�@Ő�"O�3T�ҷb��A�������"O�qiKѺ*#:�c�
�h8�"O� !�G�O�@��կ\���Tpu"ORy����n_��R��Q�ᘆ"O�}Z&"
�L],���/�!ߊ0��"O� j�L�c>݂�)�p���if"O�UY�}T��Җ�ͯ7�ma�"O��3�bS�H�u�#o�--��<��"O�i��P�tpg��4<��ܲ�"O�����J�
��d��j,x`0"Ov��oN5W0��V!��%��:�"O�I��-O>X�*�1wa!e�Ra`4"O���q%��[��=	��#"OZ�B��N�~��*�M�3��x��"O�yؗ��`2�p�X�H��4"O��i�ٽjٞT2���&J�y��"O�J���<d�Z`�blE����"O��2�L��6t�4� _�-Pa"O,�k�DO�j��@ѥ*�=s����P"O����>�ڑIPJ��A�haPd"O�<�F�-�q��/n޼���"O�AQ��L�G�ʹ��/���v���"OL�aug�1�Ryi��R&�17"O@y����w:�ң́�Z�.u�5"O��c�ğO}��	��ʑd���zV"O��0E�<j\��3�W%Ia �Z�"O��+U{��ig�Nd�h@"O��W�~� 7`�F����"O���DR'|j��� �i+�<�"O�S�˞)��ma�.��)��� "O,�
!'�e`(�@bؚ�b%җ"Oztc�F�2���.0�j5Z�"O�\��NH�^`l��ޜ-�&�@"Oj����T5��D�w��}*�"OXXs�y��c c,!Y ��"O�X��jN%4
�ʱ��)_��"O�,���É"��"�+Vi2�"O4�Is��2�2�� )i�j�"O���b�	:X��T �!R�A� "Ol	[1��s��@�g�\*�D��"O��;�/Cs]�����
�>�x%"O��hR�6+NH!A�7@x�$i�"Od1��Ε�BТ�VU�cd���yR��?@r>���>�~hA��X�M�h�'79��"~nڔ%�H�r/���ec��ȍA��C�ɍ*�T5a�P񨤂��@���	�P@�%��*Y��zB�'KN%XV/�:/_� Ie�=Y���!��q `�B3O�)��$�:L(��ǣ��y�\L��94���c�����3���x�L�v:�	<u\ a�P-]�~���D�G\�'��9�F�͉o�X�ӌ��t�0�'�\����u�ayrn"��B`䀀U^(�+���ލ��G<� `�U��?�Rm=�')���]� Ŏu�LF�&�-9���3)TT���G(<aA��rCl)g֛X���Kl���W���vyv��Ջ�?u���jq�N.sBPY�'�Y��`�]���:L��)��̚%�@5�2LOxj$�}�����S�?:��2���# ����ܸ�><S�f̭OB8*��	�ڕ�����`哰g����%�A1HϞ%�0��2�x�O�-�`lُ6�l$#f�O\%���	���r��`���6,Xt�tl�,ܢ��'OܤP��Ҳ;�Pl���'��w�߬ j>z$�UO�M9a����R ���bIVpE�����O��0�n���� ���t�O�gU4]� k�$!��0ȈHe�B�I2v���G
	tŒ����(c� N?z���(�Ly>p��a��q���G�I	p��I'��-���w�	R�	ۻ:�����,�Gx�J��>��ٛ&�����5BS�o�F�pa臵��]�0��Y/*M���Ջ�jp�(Yuy�Z?S#�"��鍵T�z��eGM�������3�d������ҍM��t+E/�^z�\#+�9����-_�X�aA.̴\T� %!�=��92�faɗ�U��$�ቼ{�ft�DWS�ڙ���C�����gG4Mb�aU�<c*��૞�z�1�:��0K�~�j��ʐ38��*�Nթ1� �?A-!�$
�N���
[����	��1A�A�$M���I`잛g�Y c��M�䅛p�����=K��ջc쓠,�x;fe��RmR�0=)V�X��B<��mK�?�2��P��,����A�P`���R�� M�AS�O���|��'��!���t���[�F���Y�r�p`�6ȧ�'�tl�f��w�ډ���T�<����oy�h*�O���!�).(� bGH(<���O�Q�Ζ�QyazRI4F{N EK��k��	�r��i��XS�Q��Y���ޱ+�$����L5ǸOXX�;� �����ZnhM��MǾM[����6*���H
Ӣhr��̸o0BU2�`)+3�8�`�ʧeLȀ�&��$6 .��BS�'3%q���+?�����-V� �X�z�ܸɲUD
[�`0Z�n	�~���B�,+��� �Dp��ˁg ,$tՒ��'1<ai��$�H1/ք-�4���C�'dt�bR��M���E=[�|0�b>	)��y9�=ʧo�*����d�#D����E�<@T%ڃ�W-DuB$@�_�T �Cb?a*S���R��9�|8��Nd���u�҂9����"O��K:�A�A�,������򰤑cA݅h�������-�D�؇oF�L�"0����tl��3(���ѡLF'F���@wX\4��E�-A��mQ�ۊ�y�o�p��\� �Jj�h��bM��'�Z�9�(�[��EE��R9d���Y�D�7���y�ԗy��#��av����+*�@U`'��,=�'V�>�IlAQEm��7�z�V��9PB��Z�H�&K��c�|��RG�42����k�lxY�*	��=ɳЅ0%xL��H�=Y��`d�R|��г�a�C\8�듼id��Js�kr`,��Z��h��'����W�ߏ@ B��E��^�`t�«^�-�:5��\���:��i�.4*�z�*Ҽ-�z5����
�!�φ`<�a���p=8V��a��d(�����,�ɰ���a�j��s��@"�U*�JI����i�z�E D�d�� �!RJ���T���Id�ö�?��Dp�H]��HGP2�3�;A�y�OL(`?z\bꅶ��t���9G�Qa��?K0��YA���u�ΰ�6�c�(�$�'l
�ڦNz��-Y0�ȴWp 0��$ۻ;+������ħLJ��� "h[ ċ%�
��q�ȓ&�� ˗���NParpꔃ;j (�'�0)E)��V	䠥OQ>qZ���R�ԭP7���j%D��Y"ꛦj�ڑ�#�ҦM���+r�ƛ��%O�l�����L�3�	_T�ܪ�O�;Q ̔��B��N���\\���'Z�B��2�l�`e~%��hB�Nr�U8� j�-��)	[�:��U�
D��æ'ob!�ת�w���K��K�f�;ӳೳ�<D��W�F0ZHrHB�� !>�D)�n??����@xH�8J>���ħl��1�̜�x��ț�*L1T�ͅ��M���'JU@��Δ8k/��s�L�cf���*&O�p!a�օ7���5�U�:��AB��'��|P�͕�.��#��,m�h� �;D�đ�d�.Ml	y���R�VLQ �/D�4�2l��<|1���+hj|��-)D�`!dJ�*�qڱ�=mj*x��c&D�d���w���Qs�L' �~����$D�����*<�j�'�[qv�fd/D��;��J�[i6�9�n�6_-��gD8D��� �#S��R��-;�P��n7D�hC3�Κw(Zy�AkG������1D����ݔD�l��T�G�Tdz��D3D��g Q.ruV4�'�	�P��a'D��f���%�P�O
����_�N$!�� .�;�'18��53�@�	J�`@k"OhL�D'
'}��Z���9A+��A1"Oh,ۄ)�	��M���_�:QR"O1��eA��17��^��� "OR�뱡�`���`�.	n��t"O�4���9I���ܟ~����"O�Sg!��)�E8���~�L�"Ol�
��ɪU�)�;ج�X�"O"MA��7N�x�g�Fπ��f"Oa�D�Pv�4��&�D�U"�"O0y���F�c�H���Z�U)���"O�������@��\�0մK��+�"Ot���JKo��܉��!!D� �"O��!�%[p]��Ep�w"O2l��HZ����� ��9\!ct"OV�q���.n�Zs�'r��U"Ol�kN�
j���׮�8��A��"O�y����Y��ηP�B���q�<aDKCp������5w��yCA��o�<��C�0�jbɚ;@qz	�f�<!P�Z�Pgܳ��ѸN"�-QC�I�a�
�0�B�w+���E6++�B��k���ʑ�B�o�AH�iY(A�C䉋�F����`n� 	d	�74�NC�	�W��ɻ�
��.D�'oI�,�C�	7,X�!F�s���P�
KZ��B䉕o��r�-ۋV`!uD��xx�B�I�\�>8ط
4p���0���Q�hB�ɾp^��q ��4t����b��3�<B�ɦp�p��'xmʩ�7 #��B�	i6	!ԕ��I�A�
�B�ɗLIz�I�1�H�H@ �=1h~B�I �@��!-4i�T�j�'�FB�{���t�8	������<B�	�����6	 10��U�΢#B䉟8��U���J�S�}1����z�B��J�:y��'�E,$�����O�&B��	 X"	�*�� �rV�e��6D�hÔ�O�n�p�I���,�(���2D�h����`��(Ѳ)����7`1D�4��,��4F��I���k�0)#v,/D��ۃ��(Y��4�-� �Z�yb�!D��V*J��~i+�㖠'� dZE�>D�`��Ϭ{X����C5>;�x�O!D������5=ʴ�P�[�>��2e>D�|�H� �a����zsX��G�#D��x�悉Dz�}q�Gӎ~-�i��!D���H�.>��37l�T��@��#D�0a�!u;��0���h�#4D�0�T��{�\9�A�ȕn��e���4D�Բ$Z�C}����>qWֽ6J3D�8a���!s�hq��<�I��D2D��j��O���%���L�k���D�1D����#�R��������f�3�.D���RG��dP][�-F�Z}~@��i9D���۸<٘`zt�ge�*����y� ��5�,1��N�?'��i`���y�Ā:�y6��&�-"w�� �yR ��D�� �U9F��d��yB�/m�P�ӤE�<>c�\�Q�؄�yr$W{<kU� �P�qM���y" ��4�q�C�? >�@䓁�y���7iq�h[���p�8i� oC�yB#E�-�.T&�5�2M��[��y
� ht���L�bE��TL͛5�X���"O�����>#�ܜ´+(�;�"O^I��C�G�N)����! Y�"O�=��jdM�8!d� �9�mAT"O��yծG�81�Xq��ۂ9	��KP"Oj���犦&�<�3��p�ȑɂ"OʐI��K�0��i�$�4m���"O�a@r`/�,x�e�P�L/2Qhv"O��1�
&s^
�)2@�9c
��"OL��`S��M�G$�}�9�4D�t� �+%e������jR���m5D�8�uM�T��`�ΎT��I��3D���׃������ *b�<�2�b1D��a���b�%�_-%@i�'g/D��C��f�и���(,�Q��*D�h�UM�))���1Ζ'��Mja�4D��sҩɪzD�*�Յl�4h��>D� *�*ʺ_-8t��	��cZ�� ��0D�܊���!a�f��S�f砘��/D�� ��L=�*��S'7/N@SL/D��P�����dI0��k��.D�|�	�W����WL�T��;D���TE�)7D��ʂGۛ�z$�q�6D��b]�Mo��y'�Y�j&��� �:D���&$�R�T�W�fl3��6D�x��V�b"�)�SEP<#�<|�3�7D��:��G��J@ڑ��#H���@5D�@F�XM��:�bܞV(��3�6D��U��(��"K��IצD�F 5D���@]2&�r��U�&�ʈ��(0D�X�+D�>�~ejV��2l��Vg#D���=Ʈ5�/�N"��!N2D���D��d�a3��ҍa����>D���+^�(�Bęe��/�	�h?D�Ԑ�#(n^����a��MiQh&D�В h8�rMQ��H{���'D�, 5��� Fx\x���\ٔa��%3D�(�6d�:���z�fʵ5:\{�M7D�X�$L�@�*�k�g�?*�}[��2D�pA��00r�y�'M���a�*4D��狏9e�ܸ1�01S>a�"3D�쫶.�8\v��w��R����.D���H���EybcK5o&�X���/D�#��߂{�H���6- �*�*O�P#�cɤ3Huz1O2r�d�c"O�l�FBO(m҅2���n�(Q"O��k"M�-A�!���
� � E�D"OTHx5A�#3�����P>*��g"O򜀂
η	�I��M_9"�{"O���gZ�P�@�����\��"O$����X�j������b��S�"O����-�-r���3���lW$��"O0 *��?O^��ρ�jz�QC"O@�#Ą̡ ��Q����m��Z6"O���U�s����EH�+h�{�"O�-
�)(̀�Z��	>ʈA "O84���*Y��1Pwe�b��y5"OR��v�-� �˳bH�e�Ҵ"OLɹ���7��Y�0�<᪄"O��� �%7�@�H��I�D0�c�|ªɄE 4���>�\��V�] &�{N�"B.��C�5*��"��%
Va	�ɠg���e+��/p*C�ɧs�����0F��`���F<b��u2O���dAٍy�<��d�[��D)��QX��w	<Z��W�lւuÎ?�ڱ���v�,P�� h$ %��y�Z����(�x�G�@U�׬D�JUn�2��4  ��p�f�I�hƙ�bh��)U�B\�>��h�a ��P�7܂!�	IH*��cF�R��'d$陰���8Yb�'ȊaGB�$�N� 2�Bw�]�'�8��B��.��co�x�'s�}[',	p�(�3 �D�H$S��֭}����j�<�x"�N�:�B̻#a�T�TM���4␹�'���2e�y��9gM�c-���`�kyR6�J!��$pr1�T�Ā2;E���n���"�A�e 0;"�7�F���G�eή;��ð#= ,3,��j{��ƀ����āïK�
�	Đv�*Ԁ��)2Q����<�T<	�背:
��O�X4@�ʉ�g��A���m5�)(O�9:��4Jm��h'� O� ����_�~�t'߽Y�*�S��O��wCF�>���zש޻uit�|:��8rgPA�E��k�DcG��;3���.�p_P��t\- �K�<°ԉ� ֬K��m1'Q����3L�{
nъT�_�qP1��K�=���y��� �~Rq�B 8�X��"���?�6���fb0�'H�P ���2&�8iZ5�F�x��z�Ϧ�'��1�B��c>D��.��x��[*�P9bC3��b���)�l�#E�����J��		cA�=b��\��gK.��ɜz�<Y���'��Lq��.p��\��ы8@Z�{�{�H�%����4�
{�O]L���O':� i�g�&`v��J	�'���jP�R(TEY"	bA���@�� O a�J�D35�<�%�C�k6 0�B���	��m|�<�F��qҺ,�t�L%JM��3#�FjV�XX��J�I�\���'��Љ�R4"
~��	�>-���<��hX' ���I����t��F��i�n$T�  �+1rfd���/�!�$����E��a�<;W��Cf�0{����I6>J$KՀ�J��yWD�2oײ��d�X�'G~��g��y-�pp�t`����H��+�T�6 g͆5'��Ӱ�����S89j��Xch�pb���To�KHP��)|OҰ�D#*��H�4*���jȝ�(5�0���~�*E���|�1�B�5Üh�ՀY�m<N-�?Y�mG�>T��3�%�'9,�xqţ�?�`T����,^(��ȓEW�A��ժ:�"�����*4ps�7)�H����>���OD�:Gb�:0��X�3�ʦt����"O��S�i��Q
0����܆U���V�'�l�He�Ҋ��e��Vr��7,�+��������l����/CR�p���M���؜�La���E���Q�OVD�<�g�Z�[��8��� �pik �y��m��W/�4p�x1a�C�ʘOH�����(�����T:0�[�'Ř�ѓ-�v�zBϜ0yr��-)����ƈ�;|���7���?E��'=��bY�[\J�9�h�$y��	�';�i���#�>�� lT�A
0���c�Oj8R����Lm#��Û�����!�P᪐86�n8��m۲z���%�ԋ��Y�g�$�q ��%a&���caɿ\)����	�=�f�WoH� �JŐd��?�&��XQ�	q�4�L1C/.�����.g��m���sZ!�H33b���0AK-Q��ҧݸ>I�I�/�xtYfG�t��S�O,j�� �I<��Qz�@�,�zͱ
�'Ҩ���Ƃ#_�M��#J50Rx��s�:}�	��ol��P����{�낊/辱 S��3�dɣ������?��+��*��H�H��I���C��p2�=	#�[������} Zu�FXm{�i��лk0џx��T�bj��a�����ߞD=�sP�F�\��D։_��y��:>|�8�"̐8P��؅D���Ę#t�8ّ+=��	�a��6
��1�Ȕ4C䉰
X��q��ީF2�ՙ)W �V�H��뉀t�ax���/h�i�DT,Cʐ��4�?�y2�)Q�0$�JhZ��y�ʃ�- 1n��H�:��?�yBd �{GP����L� �����y��@�C>Ĺ ��T�>�}��ϔ��y���85�ʍH��45�j���y�V�4Dp`���W=7AV 9��yB%d����Q�z8��
�y���� ���ӿO�^,�ԥ� �y
� `-�`G�-_�˃C�Ts^�d"OH J�fT�}�	x!ポI��帱"O� bD�I�s2�9B�J!?4(3"O�����1Q��a
EL������"O��e/�	)��41�`t��"O���B��bI�o���E�5�y�U6�­!4�F1<�u�ө��y2L�'�đ��N
�܌�1+�9�y�
5b6�� ���,�AV���y"��'P,�k�C�t�u���y���{�4��Wj�9FO`m%o��y��*��#�#H�,�@Y��"	��yL��'��i��."�y6�/�yR�ѵ	�up˄�o��䀦O��y�L=�<�9F˼i��X�)M��y��Q����f	�i�$��	^��y"!�W���u�[;m <�R���y2�ȶG4� 	%�')����ױ�yRMS�1��ӧgJ�v�fU� 3�y��#f����A"��f9B4p�X��y�N�0� \�_P�¢�yOe�z���^  �p�xa�B!�yiW�eK&X0�/!N�Hа�]��yB([l0X9�C��!	f�I� ��>�y��9m���#����2B~�BcH�y�dP]�b�z7ҫX�B�g��yr/\M�z��Ń�-+��1�g����yR�R�Y�䬁�h<)a	;� [�y��wNrXaV'��]1V��,���y�ND(S���T��f�V5��h�y�,J�,�U8@5A�xe QF'�y���2<ߺ5� �-�\A���H��yDH0�`e{����^�i�h��y�+�ZIj��n���(����yR���w�˲�V�[��X6j��y�K�E�@i*q͑�#N)�e��0�yR��	T�-��e��.��i���y"��6=A2%J�,�/i�]�4+�)�y�� �B�R��$Ó�/�<x�����y��-[�����"<�D1SOJ��y�Ȟ~��A�mN�&�Hk�Μ�y�G�z�-h��@7NʱcqQ�<Ab�Gp�RXґ�	�p Ck��<�rŖ�g�꜃�5p	�峆I�o�<�dްA:)�6�U.I�� V��d�<���ZJ���/ ���xF\�<���;R�lEjr�p��HX��R_�<Y�)�	Sv��<_"�HR�W�<�
�s�5aL_� �T�L�<�T۰�F�(�"��WG\�1GH�<)�oԠX6Y1���;*ȊA�'LV]�<ٱݥ�B���^�	�Pa��n�w�<A"�$��H�QbY�F=�����l�<�cș3=\yh��-���H��i�<a�*K6^��s0ę�ʁQ �Q��X�E~��X�`,�&���,����U��yBˈ3S�����3*���G����yB�޳r�$`ǟj� a�D���y���"o*p��FB!Os�[���yr�\�LW%9�k
�N���p��y2���Q�4�"!I@v@TB!kS:�y�MߠJ�(�F��%d�#�p?!��V6�M��a�2|��]a �T�c�&�9�)j̓a�.���k>�2�ᛲ2tt1P�5���+������#��0d��T�lsN~�/�� 6�:C��%ېP�`ƃ��lJD�Ӯ1�z�	�	b4��0|j B�0Zފ��������$l��-��-m��?Z<�����^I�P���:V* P �G�dG�L��D
t}B �J:�5
çj�İ���/_�VL0�(�e^�шf\��{qA�j��i��O=�!j�\)>`�D���ӹF�n�'�B�!S����%Z7S�b>�A�X,�r)J�JC�e(Ì��S���Ń*����t�Z����S4��=���ް �*0/ЈQ5vT� ےh)��ʧc��>���ő�R0���T�eo)��˅(R9�R~��J�Qe��Y�P>�����@2Ȫra�5
�#�bN��ЀxA���(n=q = /����R:�(sEi��*��!��W�(��@�3U�~h�Q)��v�X��O͚Rj�:z���IA�G�*Tɗ,� W��q��IL�dZT-B�����'I��3���\����8�q���ޠ:g��ZOE.L����à�?F�dȅ	C��W޿+�69@B��^�	R!Bм�em?��O��`��MA *BÈ>_rpMȄ	�)��bO�%	$���6^6��R���yҢP�Ja6\�'�C[����Ԥ��y�ğl   ��   �	  �  �  �  V(  z1  ]<  hG  uR  �]  �h  .t  �  ��  �  �  ,�  �  m�  �  y�  ��  ��  E�  ��  ��  7�  x�  ��  *  �  d � � o& �, S3 �9 �? F �L �R ^Y %` �f �l �w � 7� �� � q� �� �� C� t�  x�y�C˸��%�RhO5d��p��'l(�I�By��@0�'�F��L��|�t���pd��46���jɿ���si��w�D�K2��I��99��ӻ8r��"��u'B�]��T�	�~����Ȳy$�2�]�zo�M����;|���� !cr��;��[Z���3�1��ݞB����M����'y��dT@F�){<��e��$�ZRD���	�*�&!P����Dڞ:��7�^3�Z���O����O��D٣[怵9�(_��k��p�����?����?i-O���?a���?Y7k�"��lȲ�1BX
  �fҡ�?1��%�'�B�'�H(��O���,3e�Sgg� ��(d���prC�I2e�Z|���	�*�"PYuj�� ��D�d-Se��**X���%�~R¤ƗLEzv�I6�$	�@��ə0#
9�4��Iѡ;���',��'��'���'�O���1���,�� ]B,~���'��7�ܦ!��46/�	 �Mc�O��Fd�>q��L;�x;Qm�+-ʡ�ە�hO�D��LǮiX�P+\��\�x'�ј��<����_<̣�mN-i1���爚FQ��)�' �%uG���,���û�>� +OP��D�=j�����o c���6��oDџ��'1�f)�K"d����Βo�XH��'ў"~��$�-Z���ng#�� �n��hO���@�?u���6�F��5J?R�%h���O��O���"�3}RD<��M3��ġX>��d�>�y�&Q��*\���G�>xx���y"2�F�:�k��CR0$� �D,�y"��;au.��B��3b�-I@�V���?���'R��N ��xR��	{d����d@>k�?Q!�]2~��j[U��Av�S����IT������(h��Z�&0�(��e(D�A`�ڱGZ�-c# �(Tt���+,D�<8��q�(
���
F��@�T�*D����*��Q+7/�'LV\!��*��U�>]�4"�+p��ĳSj&&�|3bF�O<E���i>�������'�d�{ӌ��Ÿ�%չS��U�	�'�9K 3H�v4��9L���'��#$��YT����IS&A����'��x;У��d2<KuL�.o9T���'9��p��A}6�C �
��(<x+O
 Fz��I�j .�R�I\�����5a�4/��I�6����ܟT&��>HPÄ%��VQ�G/r!��"ԋ�y�iA9o����@�[�`��*Q䉁�y���?TP�w�z@\Y���yBi�> �!�Ǌ�W�
)�Gˆ�y2�P!D�f�#S�Y,AX�Y{��$��>��OҔ �-�馹���$SR�<�`����ޡ�}��_���'�"�'����-.n��D�$ɥo�HeѕExr<'�-�ax"�5��䱈y��T�ȱX� �`O�(��:�0<iW�Eݟ�����I�h����n]�6��w��7+�.��'w���n�z4��)��.�h��1K�2���D���,S!�/nP��� �_J�����O(ʓu�������y�'qF܊�Y�p~��1�������V�'⡟'+H�]*�{��)��?V��v�٠f�D�5�3��#{��D�E�ᓒxr��@N҈�4��A��3X�H�!,%���X$?e�|��� [�tQ��81�}x��EC���T��ɖI}�d�Q)�'<��ihsB΁T��?!d�0i�	0l߰h���D(Ҏo��~y~�I���)�Ñ�?!���P��^yB(�Wn�p�aU i�ұ�5j�c.�'�T5hf�'�Bd�g�V�2��?�d�!qH�0T���7a&lHօA�g�Xmn�1��'
�\�Bި-j����"��ēy7���'5剞HH
ո�'W��UJ��M�fT\���I���':�1㥠 o"
=����(7l(��S����4,�6�|�O��tV��HV	
�f���DǪ 8B��v�!dؒ�؟���ßX&��O�n�
Rl�T��;�ϐ2IZT ��/�x"��f��=AqMY!=Q��dϜ%�"���'��=aQ	��/e�9��θ>fL�wb�.�?�	�'`�pc�U�Z����e�ĳ�'���a��=c̜�e+�3b�$��I>A��i��'���c��~r�븐��#D�oR��1�PG�����d�OX�$o>��Bɀ"�A�OX�Y�.�)� �K!��.�`���a�'O�L��f�'�@�8�%I'8|]��*�2�B(�X�x�dP�S������#�0<��*����	]~�N�v��LR�)U=�Via6*�����?�ӓ R�!��GB6W�@�ӲA6{�����4�?����d�x1b�C���~,������'9R���L~��
��Ov��M{��Zپ�ء�K6NDˡ@�\!�ԁ���?at�]-+f��v$O�tP�Q���	7"@�M1�926��45ʬ"���x~R	B�s�!&�ϱF��@R�3~r����ReX Q����1<�V�ɰ�	ҟ<G���'-"Y"���?`q�ֆ�.v�(s"O��b��K(	 ��q�GU�4������h��(�c����� VR@�/o�2렏�Ov�d[�!���m��?��	۟,�'��5�s���1o��p׈�7S���MP��F݉@�O��6� �1�1O�`�޴\��
��P;�*ܜ8���d+��?I[*v-�#�3�	�z>��bDƇ�S�y�t(ևr���$5?����(������?if�U�"����a��q�����L@B䉗8��0��r���1mZ=hʓ=đ�B�O ˓lL��c��F�3F�yV.ƹD�`�8�b$DțV��I���'��I��T�	�|R#��:"I�C�[���M#w����뚘3�x����I��A��#8�p��A�Q�w��0�K͇spa~���9'�ػ�iE�xM8���x������?����?�/O��8�I#QR*�1��Y�+#�E�)F!$���ca�TRѠ�"�>d�W
1�&��8ش�?AN>1��U����:/�]�$f����H��M�� e�x��q��ӟ���O�-8D�Щk!����Ί�u`�}��"O��犑f�(�%͆?x��9C6"O�T:ge׽T���!%�ƭJ��=�"O��uM��w�� ��"�u��'�|�D
k��T5v�H5a��b]ў��sk=�'5�\ӄ�5��(@�'��H����?��ln\<ف��=1���	@���v؇�*>�9B'K�i�������,�Շȓe�iשK��H�@�	�p��ȓ%vԕ�f��#k��)@cBS�F��$�'R�8�9&��_�ZH�K@> E��%͞"<ͧ�?1����B)�$��d\&��b�O{!��n��y�m�7:qȑ��^�D�!�$G:u� ���
i �j�Q!,!��K� |�T��ES7f7Dp��D��!���E�4�嚏����	ÿ4�	)�HOQ>m���C�n�����,$��Y����<!���?�����S�'1��G�
�����M�}L�Q��~���c���ڝ�r�2-�H��W��ٸs��t�4W&`�v ��r΍��O&���t��c��%�ȓ*����ӣ㌼��$�CZ��&�@z����R��WB�$���
2w@���kI�c,"�|��'L��3(�)�!B�<N2�(��XւɄȓyHLy8G.�2v܈��e�^h�!��r�D���]�hf���0jǐ#�`�ȓ�Ap��#��Z6�Z�����0�?��eӴ�^\c#o�0:�0EaT�'��"��I�r�d�)רHK��1��A�#[��D�OR����5�bU�/e~i#�l?դ���v�$�8��]V����.nY���6��p�Cf�2eZ��k���ȓ:$�H���	=�vTbtc��<�z�F��6ڧ ���3��Q�q�7���T�	��N�$"<ͧ�?������g���#�)[b��9�ӫ	R�!��+�"������H�� �jQ�!�Ğ�U� �Q�[�$X��X�~�!�D�� Ǣ8��ή�J��<�!��Бhj%#i_�~�(�B�U���I�HOQ>�Ӄ O0��3�N�4\�^8ȣ��<� ���?y����Sܧ-��t.��j��4xBBמy��S�? h�+sa�Z2l���'I� �"O�[àϡ"��YP��U�j�"OB\wGP�ӑo�<�)�"O� aj33���b�AB�?��#W�|B�=�{$6l�sӂ%�B@N�>\ ��C��9)���If������O\��T��,��R�^m�� Q"OR���M�GF �!@abF31"O�e����}2�xp� a�J��v"O���q��+|_ꍢ �Y'8K �� �'�R�D�z�q
�*S1{��xsD�{fўd*sO!�'����5 ƪO�Q"'�Ch]���?i	�gl���	�e�	��"E�W��ȓ-%t��$!"O0�xB$cBx����ȓt���� ��~(��)@K��ȓQ�tp5+Ӧy���c@��2���D".*ڧaJ������.l��� w���	C��#<�'�?������K�w�hx5�X?��(�C b!�䊫 ��a�
L���E�E��!���ML�y
$����tJCgP-�!��Y�;ָ��fݧ.�z���À�8�!��P�
���T�in��ǡ[�I��2�HOQ>m�E�ƒxJ��%͍$j��:�,�<�"�[(�?�����S�'3%���sƉ�.�T�R��/��`�ȓL��tkՕvnź���4itp����jũG�$�\�q���)*4��I�|�2%�״GJ-R��B�*���a9�%�s?*KpHbm@2u�X$������F+S�D�ac~�11-I8]M*x#���6b2�|��'��%Ӿ�H���-+[6h#��,vi�̇ȓF0�H��7�浱�C���ȓI,�q�3&̥tj��(E� �N8�P�ȓO��p5�7]�� s�lܠ����?q�*@��jt �������%
;ў�G�?�'x��T�E!��nt��/�Vl����?��Y���1��ݧLA��W�N4�"q���d��얞.R¤�X��<��'�1���A~l��g����]�ȓN4�Y�mύ,r����Q��G��6�'woF��
s�ʝh�C��,h��ɿ�"<ͧ�?9������/��#�Y�O����2�C1�!���h����)����.�pp!��W6���0C�LLF@hZ!kh!���.|3���>tܞ��A�j�!�I��,�BweV�N��+�iӰy��	*�HOQ>��6[�h��HIc��_�dS���<���R6�?�����S�'���  J2~��"*  d
�Յ� $bD�WM�t|���V�aĬ��[��̪�e^�!��i�$-2k�=��)2����˔<�nL2$E׫]��D�ȓ<@)���	<\F�y�.�t��a&� �����4 �D�vo��*H�a���b�U�3H�|r�'(�����*�H_!6���g���x=��5���R �0�� A�P:'�r|�ȓy�(�U��'�J�:� R(\L�ȓm_\Py&؊rܦP0��\����	�?��%B6K�:�lƕ}3�0x��d�'mL�r��	/;�DԱ � ����fkK&@+��D�O(��ė��v�0��@ѐ1"G�S�.�!�Ě81��P�<m:����eI!�HxP͓�C�K8�r���w8!�d�)4��@ȕ�$�1C�'	!џ09��i
�v@�,{�X.��|�4��I,�k�O���O�d<?Yu�	:ݎTYX�
����]�<�A W	e����J�)8��+E�S�<� �`��wZ��
��y�t�"�"Ob�:��'�~ AC'�z:��#"O0����~ĸ�B�ㆀrp]�\�����=)�1��e �L?�ŋe	K�(�2�~�� ���?IL>�}.]N�\3e��)i�x��E��z�HB�	�xm@Ifʃ*A>1�De$i��C�ɢLd  P�.܁�
����C䉝MP�`���%6���0TH� ��C�� p�:��QLӤ
� ��d��O�8G~��[��~"�B�D�i�W�f�x)�ק��?�L>������	6.��Э�M�$����#�LQ��'�,�,A�,ņL�7l_�C�>Pa�'�>�2�'AAqZ���*rvx�'Y�L�-�<~x`@h�;�X�J���K��Н�!���yv
��Cˆ�hO|� ���[�+�����	p�V �	�8��I( Ҍi
�!	.{� :�N�5�C�ɳ5V �r.�(+��	�� �-��C�	�d�1�
���8A��@V�B��+� SEKƱ
Ӱt���/n���?�퓍q�z`�v	���O)0���'�N�@��4���d�O�=�z��n��+`4LX&>&���^��,�Ŭ]�%4����<_�=�ȓ(�a��\H��X�B�פ=/��ȓ(�v�s�l%c�x���ǐ�"�f��ȓ5��F蛷E؃&G)�0��'!�"=E��gE?:���Ȕ+G+(�����ׅ��ČcR����OJ�Oq��y�֏@2�ɔD S�A��"O���,ޣY����7�n���"Omq��9��R�AN3JŮUA�"OV�jA�V�%*�e�F*�>�����"O�]�wmB�Z+�,0G�!�҅!��|��8�(<�� �T�1%E��Zo��avN�c��]�	Y�I����O
y���2��sp+ױ�)+Q"OjDq0��C}�=��V�<�KW"O��
�;4�E�U��#ko:0cw"O��T�� k�-��AY�4l�AT�'��Ē��~��Q"��-�ع���Uў�JS�<�i����-��gTd�S hL̜����?�	�
��P̝_H@7ƈ�o���ȓCX��֎՞0�<��@dR�j���Pyp����<�Z�4o�0/�ЅȓO|�yc���#Z����dW/a��!Db.ڧy9R����wt(y�Ef�b�h��	��&#<�'�?������ԑ�����Dj��@P��>X�!���0P �#�W�Q�H�*0��5&!���1�B��I�:*"�� ��J!!�Ę~�̲�j�]�"5x���F!���0zȦ���ϊ)�2��g"��	��HOQ>����47��0��&O���!�M�<	q,$�?����S�'`� ��;{��A���.}�8Ʌ�Q�&�A���.�椉тJ�c�$���a�U[�#Ԯ��BA
[��Q�ȓmR`�Ԥ*%��ÒnI S���ȓdq�B�M4a� �����}��$�0���Vy��dѣ �|���b�)m���✿-G2�|��''��8�f�9p)ĳ�B�b��S�N����ȓ/~�<�D#¿4R�y�*�*f~<��@F4�t �n����3�.���\
��#��||rU�F4N�>��I��?�c��8~��w��\c�kt&�P�'�����I�#��+�	E�?c.%z�āq�����Op���^;h���� �&*P4��O
�y�!�䄯g@�3&/UF��B�^$L�!�� ƍj���?l�hE/�/	H��Q�"O�<���/[B�H�n2��2���=�h�����ԗ[[p[�/�o��H���'2��B��4���d�O��7�rl1���V��#f�@�9�ȓF/@�{w���I
�y[�E� A��)�ȓ>C"}�����4-R 7g��Ć���B
?$�Yi������@�5D�43LQ�O�J������&o�<���)�'*�ґ!CA�(/V�;�KQ�Jl1�'\Bͣ��'%|���%�adBaS�_�����%Ӧ�yB�_x�`��f��P�])���<�y�̈́�;��h��F�v����yBi�J&d=Q@lR2Us!��y�+�(t
,Ic� �$���ҥEG���[p��)UL��j��X�NH�r'�]r���O�ґ|r�'���c*H�x�d�*f�Y:łͰ}	���2��8j�iR>Ml�<Z3䔬 P����6���$Ǒ?�2��7JU.A��E��jPD8RFXp7ёt���1��|��	��?����{"�H�b �">���%(Xs�'2�����Ɇ�{�H$���_+k��(�F������O����M|L�;4�°OZ ��&�̊sW!��[&3r�8pt㇟pYP�KG%H�:!��?!��q�Nˋ72�
,L!�d�'�Z �'�"l!�D9&��[�џ�����/dnx���? T�q妚+`�	Y(�O�	�O���/?a��A�a���i"�
<FV(�Yq�|�<Q�HU �0E�6�D�u�v�<�,�&��1���5# 1z΄F�<�]@	[��F�S��Pbf hR�!������CUJO���r,Zdkp��'��"=E�Ă�G�,9��đz��e�'a��2qO0��'TnYx���G�$�b� ����x��`(���V��'���'����1�[pu�YɅ���4�����Ϛ�~��m8
�^�L��5�I�f"����դ��ŸS�Qp��6yTTl����H�H�
W���O���&�'A2�iMpG̡T��G{��#"d�p��]����&/���Z���POK��q!%�OD�'A�{ׯ��Xc+�t}��B-O>XPT3O��6�s����#�J-��1a��	dA�"I���ɦ&(�c�`�`�`#QBW��?E��
��Ba�
%(�HY�A��yR��+Vt��᎐�-�45 ���'p� �2�H�i�����E�g��ɭ"h���O>�S�K~��!]�Q�	�A� �Ɲ�y���"�5+^�iS�
%�hO^D���*�"USB�P�)��!��o���'"*K�?c�6��Ol���Ob˓�?1�"H�i��ʷ@����V���sȡ��	�>0p�B�j��_��˟����J_3.��Z��3iN�t�&��"}�n�b��>[����|���g�'�h�35	�:����`X�:p���O�����?A���y�|h�@��u�؀)���kh�UR�!9D����ϟw!�����,wT�����OFz�O{rS�4!��eET�xR��i��%��'�:W��yZ޴e��8��?�/O����O瓿z��Z���2c���� ��%�% "G@G$�2��8��{�ҙ��OZ�óO"fa�ڑ��7r-8�m�$TE)�3膩>�2\�����%�
�G~�(I�?Q��@�w�Z��ŦG����񆛾�?ً�$/�DL���)��)����B�R�ȓ>2�|j�%HEMRt�d�Ks:1�'��6��O�ʓ,s�D�i�����'t�"t��]F�pE��+ϛy�ݖ'e��'r
O'$h�q{�@�1x9(E�F�O�I�'<�LH��Ѡ6�Iq��	}����eʋ?iƥ�g�+Ih�O���u��4�$�R�� +�p����d߷@���'1���� (�.'�P	g"�#R�mq�_���	I����G22����mA+}��إO?�O|�'p��&U�^n��v�n��ԬTj�sgdh9���O���
Z*�[V�-xj6��	�/	(�O�)�$f��NmJ��fW�^��h"O扑��	�m
E$U1"���J�"O� ����1U��!��؊ ����"OZ�Q���L�J��c�ɕaat�1�� ��|y#���<a㮙{d�U=4,Nha� H��O��)�O��,�	w�:)�$ �,��d�Eę?��C�	d�B��&×a���eMA�1�C� c�p�j&�@�2W��x���0{�C�	�Lq�I�`�x��]z�rC�+i�����N����>�_������	Vn�J㇓�?�<@�v��O���i�O���!��6.B����$q4%����C�ɥkBi���?���$�,EO�B�	�#7dd�P"�@�ڂ�1tC��58���q"����HI3�4"tC�ɛw��y#�է'�@H��#d�V�)`�O�0� Jئizg�Hȟ�ϧ8��i�C�Fc���t��]|��'Y��'BIĪIh�s#6�4�L��	�~0zM33hҖJ� x��I�	�r�@��r�'Z�SWꊉ'�L)��F�e�8G|�oK��?��?i����oŶA�١�!~cM�&����?��������uI3�B���#�a/1IN�G�%�O��'.L��Y���	���M��<@,O��O0�d>��f~�CJ�CK�Z;�u��X� X����I���?�r���M�]�e�/���v��M{M<) �7��I�D�Je�	*kzX���ѝ�~�TV�Đ��S��'��M* *F�"pxH��>mʄ�!��;�	5��Iqt�'���J\d�ˎ{B��b"+W5b־�3!�%��I/�~��s��0�٤�%៎sR�i4�9?�Q&�>QC�>�tUJ�D\P�4h�*h��qǃ�&0?h��L��?�f �b�����?A'ƈ�7Z��E��{��i�����T;�A*}b!0}�0{K��sܴ%Y�Z�%�*e��ԧ��h�~��'�l��M�	��	MbVxy��G�w�X)�Z>i�<��3�@�O�s� �$4?�bi��,"6�`�kS!��KD����*OH� ���|y�铞?Z�ّ��$$e*Htg�~�D����~2	A����?�	�Y�t�	�IF���ϝb*��X��\z�ĔӰ?�6(�kQb��(غ�69�iI�<)����=�Tx�*4Ls�|�D�I�����˟��'J�맖��M�mQ6��چjB0#'0�0�!��9�IV�	4���4��6e(\�b)��(@�q�a�ē�hO��v�����*J~�ׁW�Cw�1A�"O�����$T!�aa�+��@�"O�)8��$��X� l��S�"O�,)@Ӑ8��y���:j���S�"Oz�31��uB�e@� ȒPH�"O��ѳ�0ai��q�NN/~S�p�"O~5�P#��h: $u�V;����"O��{�EL���D���;)f��r"O�Iڡ����%E������'P
�9�m�j(:ˁ�ޡ^@���$�O ��O�D�O�A'��T�R% ����>�����ş�Q�	ɟ<��ӟ@�Iҟ���ԟP�I�L��[	�✋�iS�i~X� 5�i!��'�b�'"�'B2�'�b�'�X C0+�%p⎜��o b��a!h�p���O����O����OV�d�O��$�ODeJ�h_3,D����ݲF�x��&�Ц��I����IПH�I㟖�U��Ο\���f��d�2䇉W�PF� *��Tz�4�?���?)��?I���?)���?Y�DX2����u�TXI�.����iAB�'���'�R�'��'c��'�pq�R�I�TM�6��/>o�� dh���D�O��D�OF�d�O����Oj���O�Yz��Wg�Ƞe�e��-R$�����؟�������	��,��Ο����䫃$_H��x��՝�f1�*Ҧ�M���?Y���?���?9��?!��?�)�7'vX�@�]�V�*P��ǭ^��V�'��'�b�'x2�'���'���CMv:�A1GZl$���SG�7��O����O����O����O���O���L��L@񱋖i�:�A�Ć&{��lZ˟���柈�I�@����I֟���(� ���_l8$�@ ���~�-
�4��$�O�˓ш�,�!��Q�<�@�!��8>2<H�>1.O\��<�<�MC�'D\q��H�*Q� ͱ�i(��M����?��'��	w�OD�l�b?���Z%BT�p&ȒH�����d�`S�A���4<O���g�T�0������oNRi���'�IO���O��� �tP�遾�@��a)�nXZ��TA}��'�28Oʧ	MB���i�::u��W�,� 1�'��X���J�O�I[��?A��q��HF���	�0���%{��o�jyr_����j��~�d��RO�u���*G��>V���I���<�"�i6�O"��F)!���B$^5`�	�=r��d�O��D�O�%e'h�b���T������1�
I��,�$bb���M�Ȣ=)���6�S(9c����ݍr ��a~ʓcy�I~yR�'��vi�bAg%�)��Jc��k��Jd}��'�6O&#}��u�F��(�y�A�¹`"�iR� [~"�'�F��	6��'��ɰ=��A��\9=� �+#-IFbф�ɵ���f������wQ��)��2�u+���O�m�|��\J���poZ��?�$�*P��]E-ߏc"�  1��"|Z��n��<9� 2]�:��.Ot�ik�Y����%i�&����ސb8\���O��d�OX���O���O�"| *� pnP!ɴ�ŋ/����N���IП<��O\���OIn�A�Ju��T�ߑ#����IW�{3��$���I����	 7�ao�E~Zw�#�C�#ry��9��Á/E����B�"=��/��<�����m�q�9��ٷg�B�O�4�'�R�'�"�?-�t��xM���0�#
Ԫ��r�<�US�����p&��O���q�Έ�haE���ji���C+/����4m��i>Iٰ�OZ�O��I@��=@xe��fY�H��@�d�5�O
����($� �F#p�T�iP��)D0x��<A׶ip�OL��'��72/ֹ�v�� =�sˋ�V�n$oZ:�Mk�'ܶ�Ms�Oڱr����s�*�d$�|���C� x�>��ßd�'��'Jb�'8��'�7p^"�d%�D����A	�FH�'�r�'���d�'�\6Ma��R����O�2\[%/�
~8q��J覹�ݴՉ'��Ov4�	�i��d,y��ŋ5A�)v���JT��9�2��X��ɯD��'
�i>����)�t,��3퓎1��z3�꟠��şT�I`y��>���?��1"��� �G���2�V=<PUЉ��<y��Ms�|핼��q
�-�2%�HL���\���D6Eʢ)ڇ�v�i>-K��'�(Pϓ<wZH*�ȑM�Ѝ�����j~Q�	��0�I럄�	t�O��ĝa�~�Yֆ�?W��!jሌ�d��)�>9.O��o�g�����F�$Jd�㉀��X�c��	�?�R�i5>7���:7"�]�'"���F���?�sB�}��C��<=P,+[�Li�'<�	ڟ�����0�I؟`��R ʱ��~u��� ���C���'�f��?i���?YN~z�%���2B���v�� �ǝdeX̓�^��ܴ���,��CѬ��$�.F�,P����Y��aǫF/K��	)(H-�r�'�V=$�$�'�щ�- ./�m:bF%����q�'��' ��'��Y�$ �O������U�eN
:�(����*q����צ��?VU�`����tϓT$��+PB�!Gn"iq�BL' �rx����-�'� h˥�I�O��.̗h��T@A�.[QM d� ����'R"�'���'�r�S
e�L!�s�]������c�%�����O��$�K}�]>�Pߴ��'-�(�rT[01Y%M� h-XN>Y��?�͸ݴ��DX�/��D.ydz��OD7Xˢ�ے%�)& Y������4�����O��!,�)�3e�4�AK$�	�0���O��G$�������ោ�O��%8g�P���A�L:T?V��.Oܔ�'>¹iO��� ˺x�/�iV�8�"X�R��ٲ�W�e�"Pc ��L��3�2 �J�I�Q\�(�"C7�
��S�����	ߟL�	��T��m�ly��Of��`�'r��� ���,@,)!W�'	B�'\l7�%�������O�$�r-]�}������q��(��+�O��ě�x6)?��J�����O��>��*$oL�TV6`RQ���I���$�<���?Y��?����?aȟ� IF
�%Q���	Īۇ ��b�>����?a�����<q�i��R���Ը4-U8�td[���+�(�nӢ�&������sdpӜ�	�%S,���gG�R'�P/dP�DR�|��C��w�O��?���a\V��A���YF�q#�X�sD`����?��?�+O��'~"�'3��=`����Kr�I1
ҵg<�O�l�'b6mY���)J<���f�j���r3�X�o'���.O� �*ɗtB����&:��
�?��F{�Hа�Q�:��s�?$z�i �%�O����O���O�}2�'d0h���j���X�Κ�~�q��/ �IJy��mӬ�P��9�t�P��T_K��ږ'�n����ɫ�M��i��7-׶L6m4?��m\{�p�	��R|��0$�+\�	��Q�h�j��K>.O����OH�$�O����O�7��M�84���ur��(�<!�V���I����Ia����Z�+��$d���ߛftR-��
�=��d�O^�d(�4�����OT�enR�[����)�x�vD�!�ҽI�6�,?�A� L� �Ic�fy��ŤZ�Lq �
�I�|��)�ker�'�"�'�b�'�������O� ��0f�0<���˃*]���D�'S^7M#�I'��D�O���T����s��p���ՏK?�Ȋ�M�V��7�%?a#�S�l�b�|��wcz8��o�bH��#�X�&\�q���?i���?����?9���2)ӇX:��e-<����'��'����?������~v�*a�R���E�;�R\��|r�'�r�'��q��i���1\BĹԭ�+Ji�):��I()2�*G�0K��d1���<�'�?1��?���³",A{�kM�6�t���ꌛ�?�����DWx}�W����e�TE�;s��P��(&*���B�I��DA}��'.R�|J?�Q�����)a�dM:H�lpD��R�dL��jmӢ��'���C�]?QK>�!㒆b�v �d�83�Ri���O��?����?	��?	I~�*O���^[�����6+Qj�Z��E�R�x���O��香�?��Z���I?x<����s i���l� h��ܟ|�# ���e�'s8DAv�\E�Ww�-�/�_p�%Z���6¦8��Cy��'Ar�'7r�'��?��/J*s*yZ��ѽ���d�S}�'���'��O���g���I+P���xR�K$� �Br#�	~�����O��O䓟��R� q�n�I6]������S�K� 9AV��%Y
�d�,q��'�'��I��8�ɜ+����o��N�z��,Z1^<���Iݟ8�I˟��'\���?���?��/��j���/?ܽ3뀲��'�t��?��	>�''*��T��a�P$��(]CH �]�,B1��W5� �5?�'�d���y"�G0K�8� j�&3V<�ɐ�K��?y���?	��?ُ��w�"�ǽ',TQ�J<X^�)j�,�O,��'S��'7�"���?]h���8%!�1����lo�y���X�46��f{Ӹ�X�e�^�5��m;������H��:�h-ea�p� �^t�O���?���?���?���F���)~	l��֩֊L�6�R,O��'���'������'�xQREZl�s�
�>xr  �m�>a��i7M�@�)��a� �Uǈ���][�	��\�Rt���X��O�Ф(���O�|�I>!.OtTۢ(�u�f�s &\�&Y@�B�Ox�d�Oz�d�O��D�<�`]�����w$`��&şI�~Y��-�޼�I��M���O�<����M;��'g�ey���rv�-;�(��X*����M��O�8
gi����D4�����2S�ڸ����N�u 5�'8R�'br�'i�'�>����ui�1�O���J%A�!�O���O0�'
�'�6m!打��-��=;�e�v����6M�S��֟����?�hD����'��	p̎-���Ҧ��
<:�[�O�$����I)m��'��i>��	�,��?L�]�SJ=���HǄ��P�d���ןp�'s�듮?���?�ʟ����&�vi��p@G6c;l��W��R*On�$i�� '��Z� ݃1H-��KD2A��E	Ч	����@"?��'E��Ā��E#d p��'j�(�hTG)@<���?����?�����'��W۟��LV��u�G�)<G̀q��O��D�O��n�Y��	���+�M��Ψ3m����1�j3%,ۛ��m�VLc�.g�4�5o,�P���~�d(��ܑ_�<��E�-V���C�'��P�	۟4�I�$��S�D�^ '82����'s5�"��>�����ҟH%?�I��M��'� R��X�}�H �B�9�����?�O>�N~Z�E�Ms�'v8�`G�r*v�3� ��t���
��*����X$�����'�4��I�~\��x��M�v><qP�'���'O�P����O���O���Y�T�<8��$����� �����\j�O�<mZ��M�x�՚Z��fL#<4�T��.3f!�'h�\�c��'|��P!���V���P�<OPXht�ۡO0����,���I��'���'X��'��>���tI�����7�zh�#�,5)�m�I���d�<�2�i��O$�i�iT��o�)j�t8;��+EU��D�OV�$�O2��Ťx�����Պ�~چb�#PIk���t���H#)L��'����	⟬���h��$@��1ycc:ϬLJ���6>��4�'t��?A���?�I~�A6h�r��
v��9@G
��_�D�z�S���	ڟ�&��������
SD�q'�� ��J��V�4,ţR&[�%�'�Ҍ�T��X?�J>�.O���h�)z�ɕ%\�JB��R�Oz���O����O&��<Y7\�H�	((@�����qJ��	8b}�	-�M��'�>��?��'h�x�D	�_4x�5��Pkb�bH�0�M��OF��V�G��(�2�l��Q�fπg}f-*�`�!K\��O����Or�D�O���,�' 龕���@�%��b�i�Z�����ȟ �I ��D�<y�i�1OM�b�ވ`#�	:��F���S�|��'z��'��kD�i��I�@5�����@X�W��)%�U����\��"�Ī<�'�?���?!A�9�iPK "�� Qf՘�?�����J}2�'$��'#���/�b	1��R�>젶g�Y��˓���ԟx�In�)����Xy�����ٛ  ��4�����(��f����S�L��d%��M5D�,�;�"]�p����۬���$�OH���O��d2�)�<ѵ��� �x�s� �tȦ��&̢B�*�XF�'t��'��6-=�I�����O(��l�+J�,`�L6�R;A'�O&��S�R#�6-%?��J�*
^c?��UB>��=KfbL#,��ĩ J�Ox��?A��?1��?�����̩2���,�yPH�@g�I�P��?���?����o�b�ɬ?e<Y$j��� S�M,����OI%��&?-�tl������h��kG`� LBt��R�W�\�I�v^V��'p �%������'�V��
��mֆM��.Ňiu��J5�'���'��R��2�O����O���R�mEZ���j�Ŋ�rn��8تO��d�O��OZ�[�C�G^�ҒC�pV:Ua�M�<aa�F�/�f�ش#�OU�����y�Kءf��$P�+/	H�yק��<���?A��?)��i~�4@1���%/�ME�`;�`��kD���>	���?d�i]�O���˅]�&�����}�!@@� ���d�O��$�OHq��y�"�Ӻ�"������W�"�|2®� 4ܺɨ%�iB�'���Пd���$��ƟH��~�)(t`g$"4K�eXD�'9 ��?���?�H~�b��d�:]�Z��m 6#�P�`Q���	ݟ%�b>=!�S�f?��� ���\j�@v�lhV�:?��̋�$��������D
`��� p��!@MF��3h9h�n�D�O����Ot��O�˓R��	ǟ���]�H��i&n�!Rh�X�Y��� �4��'�^��?���y�k��;S�����ܘ<󜈹k�7c+� I�4���Z�jߎ�
�O1�OM�nD�9�@�
O���y�Re����?����?���?�������"�ō)�Ҝ٤�O��L-{��'�R�'�fꓧ�D�ئ�<	B^�U������7-�ЂA�IE�����şS�ϙ��q�u�D���n��A,� �B�Z�ܽM��P��O��O��?���?��r�*;��$MB�bvB`22!r��?.O���'b2�'�R�?�[�"/0�5�A��S�i���<AbP�P�	֟�$��O)�YX�i՟L���Y"�
Y�z�ЕK&��شr��I�?y:1�OT�O2���@�wz�րZ|�É�?����?���?9M~�,O���&!#���'��#�ʨ�%�@v��<�i��Oب�'���X�9�!@�60*dB`f�-R�2�'u�`�R�i��	g(|D�����" n�A"�@>�I��D���rR����۟�������ǟ��O�L�x@�q]��XT$_�S��B]����㟸�	_�s���ش�yү)Z��!5���T��LY��?����䓵�O?r���4�~bg�BVnM*׎М3���b���?9d%ڤc���w�qy�O2ə�6�:YA��O��ä��x<��'���'h�I�����O����O�a��X�b"�!��� �U+A�(������Ȧ�PܴCf�'����I�m���7 b���r�S����zߖ�S��.?ͧ6���$֝�y�f,*۔��&�Ǿ@ք�;�o9�?���?���?Y���c��Ӗ�D�&�����K1��S
�OL�'\��'��7�!�	�?=x� Kd��c�j)p�R����HП`���
�4n�h(ش���U�\�^a����u�.]�fN�\ö�Q�I�x�����+����d�O���O��d�O�ۀ(�l��SB;\�P	�gA�	�Tʓu��I柸��Ο'?��	�m��� @J�d�P��杼E)��O�$o��Mӧ�x����ڈqsnU9��ڑ|P̫�����]� ���D�']3���*�t�O�˓]0{2�ȘX���H��ߜa�Pu��?���?����?!(O\��'� Ħ.KiC4NW�C���w�U�O��q����O����O���	8;��]fo�U���Xt�X�;���7�t���c٦��&.�>5�;7R*IQD͂t�Q;������ԟ,�I�`�	��L��P�O8�q�S �.�6�z�ǔ(¤2���?��g��Ii�$oӌc�\�V#�FI�":E�8l���NE�	��M㤽i~�$�(e�����p��r|�� -�p�h2��T�`�&�1��'�b�$�ȕ���'���'UJ|���ŁR����A�8諐�'"\����O&��O�0u�Q�b�R��e	�=쌘����iy��>1���?IL>���a��)Q�)S`$��`Ӝ�R�鞽	������d�:��$3�D�%F����3��B�4"��95�����O8���OF�6��<Ʉ�'��e�!�S�%Ɋ�7�L�Ja��j��?I�����D}��'��1�t�!}�>�K`�En�I���'��D�	ϛV4O����1T��y�O?��?qiF\{qA���.���Z�l�6�Iuy��'�R�'���'"2�?�*�K�+_ώ�a�(�,\����y}B�'��'�� m��<a�퓞s@�+4��=%���h�����	y��_�5��l�R?iC'�b^�u��M��t%�����ܟ�*۔	���=�D�<�'�?	�\�P/�ę�D�}p��ǩ�?����?����VX}��'���'��81KտN�D�d��G�������v}2guӈ�n��ēY[n@����X2���+�x�L�����?!'C�8|��Ѕ��N~�O�����W�G)h��Yx�d˨0�Ʃ����1���'`B�'��S�<� p, ��x��Đ�,R)@1�q��'!���?���T9���|�'���bU17�te�5@�{�.�P$ώ={S`w�R�l��MFD��M��'�"��.E����07
4�;��]5R���*'������ĕ|[�t�I؟��	矀�	ܟ(#)]��n0H�$E�`W�1[�I���Ľ<i���'�?q�L�&fX��w���Q&�� ���4�M��i�`O���8��h�m�S�.L�[smڎEj��4,�&>|D˓k;FA�c�O��IM>Y-OP��E�V���Q��n?b���+�O����O|�$�O��<�$[��ɦ(�x ���$r�x-�$c�GZ������M�L>��	 ��:�Mc�i�����Md��3�ï ��y!�+�:4���i��D�Op���c��:'�<��'�yWg,]�����@�
fP��C�?����?���?����?���)��s$Ms�@��dNz�h���	 r�'2f�>!���?!�ig1O4����� ���bC&�����|�'F��'+ ���i��i�qqPf�s���h�eyu��V��������D�Ov���OH��E�c��p�q䁅_w�p)�	Ä!����O�ʓ]�IΟ��ٟ|�O`8[�!Ŋ;'x��3�D�}V��X+Or��'{��'hɧ��FZ��hFa�6V��K�(�T_�����3~3�7�FBy��OZ�����,�Ջ�Y�G�&�A5��\H�!���?I��?��������� ��C�8p=<d�����Z��1s ��O��cě���s}�'`�0��E�-#a�����.3�\�BŨΦa�ݴY��9s�4���-na�����1�H�'_�|����_DU8ԩ&٤2:Y��zyB�'���'�"�'2��?�*�i�Nd���L�&����]}R�'a��'���y�eu���ɪ[��XV WZ�3��)^ꀩnZ��M�x�O`���O˨���is�$ʳC~�Qd��'A����A�%��d����H��-ғO���?q��7+H���0i�L��vj�&B<����?1���?�.O`��'�"�'�iB�x�&��6l1��T����:Hc�O�U�'�i�ON����!+����T�`��4J��'o��>I���zU
�!���������F�X牐%�*��g�F��*T��22\�d�O"���O4��1�'�y�f�h�^@*7*_�.���!�?�'Z���'O�6-?�I�?�3����u��8 R�Z&k��eM�ݟ��I��	/k��l��<q��H�~-��~��N!Ue����&��:�pg�P[�Iyy��'���'�B�'u2��|x�MzC�ė$�<�a`��I�����<�����?��a� �0H�Q���̃�_lqdQ�X��4/țv�+���A�As���q��?
��M֬,i
غs��>�ɭY��t��'1|�'�p�'�8��O��F�<�S�LA6�Yq�'��' 2�'�^��p�O����6]#��І�̛oф��%��MZ��DRɦ��?��R��ݴb���O*M����v8�K����	�iS�N��V���;�E�K����ij�Z�%�10�����˜)�W��O����O��$�O ���O~"|B�G�3>�"��B]���)�7�M͟0�	̟<��Ol���O�Alb̓lze��R2s���iC�u��hH>q۴u�&�O����i���OX<�����\�x��A��ƀ��^ �.���B��O&��|���?�[���b���<񌕢��a�������?	+O��'�	֟�O%"	2kМA4l�9�
�,��)(O���'�R�'�ɧ��1p���%MQ!iuxl����1K��EA�"~ˤ�ƞ���ӄE�"�]O�M4,D�qN��O���̂>[r%������ƟT��v�My"��O�2&� RЩ��a��j!��'F��6�M�Ra�>Y�A\�+'�O �c�%�	|�����?�V#���M��O�B���|��W0/I�}�#�˩{�LP��й�?�*O��d�O��D�O����O��W5pPG�[l��K���T�&��O��d�O�$#�9O��nZ�<u��0c����Ճ �A��������	l��i�S�g��n�U?qs��hjthP!��[zZ�I�g��T�F@W��-��<i���?���~C��a*�@X�³���?y���?������PC}b�'V2�'���ز擁՜�ɇҢ1� ���v}��'U��|�F�i~Z���"��AK��Ѝ9�IOR�t�&�]٦��H~�T��l̓pY�Iyre�(*��ѥ�E�����ҟ��I؟t�IK�O5����<]@���(i���I5 AB�>i��?1ıi��O��iP�9�v02�MA�Xh���$d�d�O����OҙSt�m�|�Ӻ��CQ���4��/C� :�)�� ?�I	�@�(��':����\��៸��ş��ɖ3��<{d�C*&� �F6O�E�'b���?���?AJ~��� ���3 无%�.�Pd��a#BI��Z������ '�b>�HQ��5��X�p��&Iˈ=�ч�+|-�tl3���	�H�{�'W�'���X����%U&�e��-&\f������ޟ���ܟ��'S���?�X�T'��� ,�8��`�E*�?qòi�O@��'0�'e�Q(WY�e�ގPW�4�0 �9*��+��i%�	�xx�$c4ڟ������|
T�b��$L��B�G� x�d�O����O����O�D'�g�? 0d8�-� �a�S��+V�"h���'���'�T���ę����<Y�(�g�*	�F�5_��̹�A�ݟ��IΟ,�$[禍ϓ�?a�F]�1��K�+�T���Ǝx�����꾟\%�������'���'N\�s��)V� q)�b��-Њ��"�'�\��[�O���?�Οr�Pdլ<��]�uAV!_`p�cY�� �O~���O��O�65�����}wF�ha'	�e&$1j3�@GA��m�N~��OE����!W�x�U�U!@d�2E�6\�-j��?��?�����'��HƟ��Qd;��%�" L��H ��O$ʓc7���$O}R�'��X�D�%'Xبu���t���'r� ��af�V���qd	�0����@�l�%%Y�A��AN�J����'���ǟX�Iş��Iß��I���/V�	��>r�-��fܘ3f�	`y��'G�p�m��<�p�]�g�)�Oȇp匙c-�蟤��[��H��H��nz?�R朁Le�H�Pe�~^�YC���۟�4��=
S��:�$�<��km	$H�\8�$�{�UAc�]��?����?����ğa}[���I�q��8��N2A��i���T>ڬ�?�qP��IڟD&���G_3OLigAVQdh�2�\jy�	Y����U�i}�i>a��OP��#*���8��yc�jte ����O��O@��4ڧ�y��^�����O�a%Lt�6���?�4\� �I���Rݴ��'}�T	���8X�Ug���Qѭ�%|��'5�'ӘaR&�i��	�m^THcUY?��5� $�X�Af�2��Uztk:���<����?���?i��?�m�	58u*Q�	Ox�g(����r}2�'���'$��y���j�	k�];.�XYu�^<��듦?����S�'��y
���eJ�$<L�vp���M+�O6���4�~b�|�Y�\�@����,-�`${^�+��_���I˟<�I��x��wyb
�>���n��\sY	�u��.3�����۸�?Iw�i��ON��'�'�󤀁RT� �h�9u�tQP���
-Ď��4�iY�	�M��# ��)U+ue0��N�#��������I̟`��џ\�	� E�Ԏ�&�vQ{�eF�%?`<�Q��?A��?9W�$��ҟ���4��'ߌ!�h�+(�=ȁ�S�M�O>���?A�,d����4�y�֟P��}�5�#d� -�liA��)kTp#��O�O���?!���?1�@��IZT���Y��bo	�/������?Y+O��'���'\�?]�M̉#�n�k����NS�0QF�<ɗ^����ҟ�%��O���e ĕ^�l���ߝ5?aP��/Fѩ�4��I�?�p�O��On�Q��M�vW�E�t�>�0L���OD�$�O\���Oԓ��˓a=bk�#4��"p�f�v5J'���?a���?Yмi��O��'���K
-�vY�U�	�n�Z�ZX~�<*���?�v��4�M��O�.N��Sy�#�c@����G�G>^=c�X��?.O�d�Od���O���O��WW|5)F*��v��p�cḴTb�
�OR���O��D1���O�nZ�<	�aۦxj�qqO  �@@�g���ɓ�����`���4�~Bĵ_t�q�p�I�g��w��?�E�Ŗ��ې�䓆�4�B��T�"Ā�4mo���K�>\�����OB���O�˓��՟�Iޟ� aǒu~h��˒09�0@ a�W�a���,����5P�9�0��	?�P��Z3lS�5I*O�4xD`�&�fM�G���S
L1���<�H9?z���5��-/Z h�3�Q����	��������F��:OZD)jԄD�9�	ˬ&fh)�'����?9��y&��������	0&�=��\-ή�i�I�O���O��n�2;���o�u~�gC�(�˺k�&C�@�#2m�q\ZLAAy��ayR�'���'���'�; ��أ�A�JP8q��eR�e��ɤ����O����O`����) T����%J��|���^�ֽ�'f*7���K<�|��[@k`P)&f lЍZrX�dd����F�����!-E����͈�O�˓b��2�@s<<Dj�T�@�@!��?���?����?�-O��'�b��%
Z��ec�)M�u���{�J㟔��O"���O��	-6R�K���4"�pk�M��h��g���YV�5�R%+�'�y�e��g$�m�k��<�N�1U���?q���?���?���?���K���`*њfN9%l��ET�'��$�>�*O�n�S̓h�~��%Lѯ<����΃'��]$�����P�����l�|~Zw�~�s�O�o.�da�ɉ�U�(�@&����*���<���?����?��N�T�N-	�l�)�@�Ҡ(�9�?�����dq}�'�R�'�ӊ1���NI�v����ӮX�B����0�	q�)�t�R�a�65�գ�/2�9Z��R�����π�M�gU���*T}��+��U?<,pzE�S�<��YH�Z�	�O����O�D�O@���ʓ+M�uV�J@$J��C(��?y/O��o�]��N���՟����N��`Q�cܦmk\�A�ϟ\�IR��o��<��Oi�\Y�ӟ��-��M)��/X˦ٳ��ݛ[My:�����O����O��$�O���>� ��r��F�D@�)&�C+��ʣ>!���?����䧚?���i��D�8t؉v�ѝ<'�`5����y��'$�'���'l��.Z�?O>��s�V�l���1%��� ��OZ��M�~��|�S�d��͟�k�AW1/1TpiJT�_��Mhv,��P��ğ��	Wy��>�/O���[�9�Wd�ה��@̺�㟸�O^=nھ�MC��x��=Ϩ�8��Ǜ��}�q����䛏z7F̫�V?���r�������.�a�wL١v��ZeL�AS\���O���O��=ڧ�y���i��	��A��T����?��_��' 7M?�I�?� ��,	ф�j��8M?y�p���L����I�CD�Lo�g~RNӛ@�2��κ��AR��K5�̵A�W۞y��'��������x�����	d�d)�5P8i��={AJ,M���'�8��?����?1O~��B}P�QEC_��=���΃V���eW�|��ǟ�&�b>�:÷T�*���j�=����,�8i�DlC~rǹ�-�����$^�&�\�S�ʆ=7�����#�D�O
���Ox���O�ʓ#���� �Ƽe�(1Xa�.=�H�i�ן� �4��'����?����yr!U
.t�*��Dc�`�J͌�HOV��ڴ��4$��XP���o�A��� J�@�ↈ���Rt��OL��O���O���O�#|�`�I1�z��Y�8�J���e�H�	����O,�%�F��(~*�"F�v�84�C/K)Y��'�B�'���I� Y�F����!C���H�(|�u͊�p��ak��'D�%�p����'U2�'w�0)w�! *t8� �2�[2�'8�V���Ot���O�D!���[�
���0�EЁ0����Fpy��>Q��?	H>��VYW���
P�RA��*�!�QiU�u.�P3�������|��
�(�OK^�T�FIH%.uA��uk�&Q�'��'����P��p��?.i���C"j>\�4�1!b`�	fyRrӔ�l۬O���EB}R�j�,Mϲ5�Hͨd?j���O��Gt�0�S����'�����EE�05����B&Rz� *!�'P�ʟ��	ݟ|��ğ��	W�$[-����w"��
��*v���	���I�$?���M�'���c��3�`P
Z�*ㄘ#���?YI>!H~j��ڄ�M��'�I�S��"ZI:���	�́��<h)��OXA�I>-O�)�O��p
�.��(Z�Y+%F��9&/�O����O���<�S�8��՟��ɞ��j�X��1 �&�V��?��S��b۴/��V�'��P�/���!��Ҧ-�Â@ɓ\�J�I��i�4i�Ox�xI~��Or� �'����iъ#���c#��8�����?1���?	���h�*�I�4L�aa��>Q��)�%A4h����H}bU�T0ܴ��'��� õ3� ��K"uQ���͕��2i���l��M��с�M��O�0 �)X���v"O�S���SA0Y|xȔl�x?P�Ozʓ�?y��?����?I��
q�m;ҊH�n� ��b̒;j��hZ/O�m�'���'Kr���'��|8FbY [gXthÆ�/��5J��>9вi7-U|�)�S�B#�e��"��!�ɰ�D�~���8�(��>)�Q�'x���փ㟰@��|�S�x0�
�4zh����#�8_��iA��@�	ʟ��	ȟ��Icy2	�>���Eᾖs;0�ia�Y*�ᕨ�`jߴ��'V���?A���y�1�h��B�# �(�� �3X|�rڴ����Kθ�r��ޅ��Ǜ4����FZF��� �O|���O����O�x����%�'m�i��t���"d�)��d��ٟ�����d�<�5�i.1O� 9韧|��#��32�tu٥�,�D���]�ݴ�z�.V��Ms�'��㌶C��X�f�1(�䁒F�w5�}�bJ����|�R�@����	ş�U-�(&Ax����ä��aH�]�p��{y�>���?����IȘ6vT���@�-z.��կ��:Q�	�����O"��/��~:gf]A��m7gED�"��ڵsH�a�"O����'��TmK|?�K>�Ə�D�`�%� 8~�6h�
�?����?Y��?�N~�)O���ɝ~J��M
=7���a:I�h�d�O���Aڦ}�?&V����2)�"B��-�>�s)G u����I㟨y�]Ϧ��'�����ed�;��%2���z�X4�h��a	��	cy��'���'���'�2�?qa�ϰD�z�kU�WC���2cO�D}��'�2�'���yB�wӶ牽|�S��@��v����˦ 6����O�O���6����x�^�I���i�c�utp��H�?��P�!9B�'N�'$��ӟ��ɶټ�b��;p����2���Gx�5�����	��'�D��?���?��3Sd!����,P\-���=��'����?����3]�9PFʹ|KT�+���;��В-O�-!�n{�p7��n�Ǧ��Eh�
]T�yb�b�L:B!�yW>]8
�GNm��M��=(�@86fՈU��Lєa�v��z�#�U�=���	se����)��c�dl�@/^�.�9@����)�WL�R�pB4hT��y�*��w)�ĈEk
�s���Mޙ%�D���]��(�&���Ub�Q��O�?	-�]qT̋�w6����D�
��3��Iє�٧�r���I�K�.�)"臹Q�f$����iJ(�0�n7H��T�@/&0q;�%ƞ���֚E�6��񄑲{hh8l�=h����m�? ��sԨ��|�x!�2��0�0�⡦�1Y�"hk�=?)�c��+v�M3E�H�O����!�Y ���33�$r�qa�**i}��$���Z�V��'8RA�s/��2|�rw��Ӛ��e$̷8!뉄�q������]����2�I�@� �z�`���i�킛$���i׋��]�0 �%�P��1F@�M5��a���W0x6��w9�B��h��ؤ��,v/FQ��b�&za�q!f�ܗzt����Z�F[f�s��Q]���87�߮x� AD$F����'�����$�OГO���O�}�f�Z�^P�a�F�����c]�<	�ښd��D�Ov���O\����ӑh����� h��4�C7X��<�����?���;g�I�'�4*0* �f�h��I�)�ٚ&b��<���?y����'=��Sʟ�q�9VD 0��O�=����Ӡ�̟���k�̟����|�� �	m~��؁�����@I*1;���?����?�cK��<����I�OD�D�O��5�^� ��u04#z`��!�?��O��DG�B���d;�ԟ~ӑCC�Vڀ�� �3�Ј`��'����':Bam���d�O��D�O���'���Z@�ʫ,�>ɠ5bR��q�'���'�����|±�	�bu����,�,�1�ʫgF��{���?���?Y��?i������O���&�h�[��?3%4Eb�E,~��2Cx��y2�lϓ�?����7�1E�5�$��c�x��	ɟ���۟���`y2�'k��'����h+��
����	-�J�I��O*�+bK�O��B�7O:���Oh�D�wQh� W;/�e��N�&���d�Op���v}�W����G�Qj�Q�m�.쉡Dןx ��'��:�'����'s�'v�?�r��!U�(�S �W�%Kب�C&�O,�'��	ҟ�$���IҟȘ��[�;L�a�w@��.k4�yƎ��V.Z����Z�ԟ��ɟd&?ys��d�"%:gd�-f�lk�A�+c&�	cy��'G�'N��'����'���3m�E�Ju��	@%JH���Ӟ�y��'���'r�Ow�'�?�֮��	 �!�G�.ʔq�A���?�����?���O�ʀ�y���}�FHD?^8Z��π��?���?rLJ�<I�	���џ|�I�h��aNkOB��b�2qt5y�Jz�I�0�Ɇ=���?Y�O��a�������a���Q�9��͓�?9&�i�2�'
��'/ʓ%9P�X�G��L(caD���Iy��'���\>�e��	��4"��-i��̪V��1aN���㟸�޴�?i��?y�C҉���$S9Z��-)�!
9f[Ъ�L��?����?	����|�A
��<��s�x+�(#!8�M�F���q1|ð�io2�'�2�'�O���<��-��
�>���I/X����d��<�IL�	��tS,?+�Dp	A%��U6L�A(�$�("���O����OP˓���$�	8u��s���:`,�=�D��B.x&����<x����?��|��'%��QSdIg�X[�@pÖy�����$�O���2�	��TΓg�N�[���X����!���F���	z�`@z��#?Q��?ͧ��|>�16�K
��ת0D�c��=��I~��?�/Or0��ņ�H���$jU$%�u�6h�|�f��'�'�Y�$�Or(�y�ˍ@����=XP��6-�<	���o����t<
}S�ą�~�z����\??��'�B�$�y��'�맖?����y��%}�r�[�!�O��������O@��.�9O[v*J"\Q���3.H#+���R5��O\�9�
�<y��?����?	���ĕ��
 �!�]�#n��b���ji���O�˓qTXFx�Ou��KA�R(zD�@�5'	f�*�fKZ�	̟D�	�T�	��Ĕ���ȉN�n!� �ħ#�աS�<�m`p�Gx�O��y�'�.�&T�ș	���cf��87�GJ�t6m�OP���Of�DDN�)
�'�R��F��@_D��BjZ#1�)z��?L>	�k�̓�?��?����+P\�`���h�G�?���?��xʟ�O��;�"ќn0,la �ؾ"�$C֧%�$�O�ٸ!��0��韼��<Qr�L�y!z��C�R�kجm �oן�'�R�'�O(��c�PX���#g7H]ڣF�t�5y3N�O&ŉ�lB���OH���OJ���]�+���b�6z�\r�Ĝ��d��?I������4�<�N�>�d[���dF���(�p�|��<O^��OB�8�i�y��'a~Q Y�cO��8�!�1��D{�'p|\��S̟��O�ؘ$L�`�V�xwLV!e�����?���8����?�\?A�	�x�;2��ы��J1?Fԝ �4b�ֵ$���'.��'���yBO�	)���aҏ2ך%YD��?DQrU��y��'I>7-�O����O�$g}r�J[�΄��N�48��ڗO��\H��'���>��d�<�-�n�r�DQ�8�Є3�/pV]�!�_R1P�$�O,�n����Iʟ���;���<�2)� 	���{v*Z�K4�؊f�:�?��
O�<�����$�|B��S�|�#�v(K�/^�°����6� ��ǽiQr�'���'
�����O2�P�� `�(�'�Ui��M3A��˓��d��2���ѿ	p�	�O����O�P�2��,�0��K�~9@{�-�O����OJ��'q�I�ؖ�~�ɯظJh�O���P啄��
}c�d�*(�����O����|Γ�� ��1���.}��4@��@6.j��s�'�����$�O���?Y��?���-ȸ�)��w���r*B�׆��>.�s���?����?�'���?)S�.S�Pl�s�L�>5�4�6,�O"˓�?!+O �$�O��d�y����#`�Eㄩ��52�p%@SM�T�	�'���'S"����~R��0-���� 	��h�IVg�*��Ĉ��?�(O���O���NL��*?q]����$�&mW��S�;E"�'z���y��'*�'�?!��?��FC�%�tqh6N�G1ڭ��A*���O��OHm#u��8�'�	H"r���@ C�J��)Yx,��'	H8��'���jӸ�$�Ob���OT�'	�x��Z .Y���&*ѵp	 x��'���'�訜'�2[���O6r�[+Z"];L��t�ӿC�4��\�"�'|<7m�O���O���Pg}P����:'E���%�D0�4�%�ܟ�Y�k��$���O�>݉�'J�o�f7��@-	+~��@,�u��6��O���OH�$�P}B]����<�!��=?0�)�K�w�e�0�����IXy�*(�y� P�����'���'����B*[�V��͢q�P��>���'���'������Ox˓�ywZYbB	H��F��ٱ@%���"��$�*��d�O
�$�O.�'f7�Jċƅp��\:�肦2cX-�����<Q�����O6�d�O>��a,W�S�j�iqm%�&�!�e����d�%i(�$�O���Oz�'�?�S�Orx�b�R�~4j�a��
�Gi�Y/O����O<�O����OA���O�	x1a.a��ZV@�M�`M�7�C?�y��')��'��O�b�'�?��e�(P%~X���T�|���y���?	����?��� X�����H�{��許`F1%�tI���x��';�m�(�y��'~��'�?I���?1D_$'�A���'�ⅸ g"�䓍?��(���Gx�O |	զ��1C�<����z�m��.��̓�?���i���'b�'K�ʓ)7��9�Kҟ%xR��3�ǔC�P�Iޟ���A�H��e�IX���2y^,-��w��/���Ip�:]B�'�7��O��$�O��du�	ן�jl���6���7E6�h�+�����t'���O �$3�'��ʂ�p`���$����R�^��*6��O��D�O
��E��?�'@���Q�>$��J��<%b������0'��͓>4����?������V 3�dP��g� ���+酦�?��?AV�xr�'��|b��,C(�B3�T:i R���"�>W��I�`����	5��Iџ���ǟ��OU�p;�;R��h� �[q�y8��ʉ'+b�'��ǟ�����Ђ J�}rh�p�솞/� �O�/5��ɴ5���ɟ���ٟ�$?Y)��*�J�F�"=�D�Z"*?T[�Y���Iџ�$���	�<ɵ��������@Tz6#Ɗq�����Zs����T��͟<&?����O	,i)�m��@,�i�#�Ux����O�O����O�<�7Ov��,<"�eόW��<S� &�^Y�I����i�g9O����A��'��'��(�[.}t(x����d��|�'�r*�&�yb�|<��,�Uyh÷�H�Ddj6�'��`�'-b d�B�D�O&���O���'E�Y2� ��(ui�"�����?1��X\F�̓���򩃮iN�*�)Y�h��e�%ςX[� �O����֦5�	��$���pˊ}��@�MWށ�p�*%�l�7㒂&�b�A���|bU>�H��`����~Mz�%ȗ8����%�v��Q�4�?���?���M	���4������J,���Ů,�B�%�O����d�On�
P;O4�$�Oh�$ي؞�S�.�1��Р��'~�����O���WH�i>aFxR�ƪY'f�sG��]��4���Y����?�%��<���?�����O^V��֠ۑK��3d�F�� ����?Q����O��On�$r�|�d�\X�$j�l�6B�k�OX\2r�I����O��$�OҒ�6q���>�h0 �:v��=1 �F�F���D�O����O(�$)�I�xn�m͓�q��!�@�D��U��Q8��w�c���ğ��I�?u�O/��`�n�qJ%���܇@U���%��ԟt�Iv�ԟp�'���ZI�XiĎ��XG��[_����4��O`���OL8���Ol�ġ|��?���%:�bZ>E�	��h��dA$�I>�����5�����4
�HzPlX��17&F;�?QwT�<!��`�v�'�2�'d�o�>Y�ȋT�
�"wFļo����"R%��U\�����O�-�/h�:���us�\4�1`Fj�=�?���?����?����?���?i.�(A��-�SQN���A�n���'�HĪ��4��[tV�,��/��;�r�I�&���lh�E�1�ڙX��T�
Ѓ��YH����o_�9�~�	YO�r���O����*k�(�Kp�	? J��ֆZ*Ry�6M�Ǧ ���?����H~����yw�ϝ( ��w!
�}�4	�c�|��V�
�����:l�T{q B9Oe�ܨ�!5s�ycwBM�	;XDSˆTR�� �IG�lU�1�աx���fB�n�tj�k�MJ���`:l-AOJ�@xQ�ޫ
P�	��@�^y��;᠇3R�>���nS1w������&%a��
N��s�n�#1$�r"$��S�L�v̬��GjT?_�0�gÀ�y�E�!g�%��B�?q$��:�Y�1���['o�H����mW��[0#{3��RvA�1e�iz6��(�T����9�E�`H(xH؂�.@4ք(# fX,��ʢ�t�����O����<qߴ�\K��~t�d�&�=��
bN�.0@���QKiR���e�3�)� �a)�JS�}�bE���L=��5�S2����1�$p���E"m����',UbA�K�H��᩠�.��1G�4?�cAğ��Ie����G')	�у�F�v|lQQ`�y�<�D���8T��I�	�`IL5Quf�v?Y��)�*O�a2���n�֑�H�.rq (�m�t�o��������'���'���F�:�2# ��d�P�:�F�^���bR6#m� �w؞�%� ,������S"��[0+�Ψ	�K��/���3ۓ6�xl� ?�`q���8=x�T��-:	`��hO#=�c���8��$�#�@�L<$�S`��d�<���_+o���)�I�*/�|�g*d��Le}�[��J�ϙ��d�O�7mĽ^�M{���b�ء�9sF��'+��'�r��'V����QD�#R� PI���O�B\��icO�%�&!R��[,Ǒ����j�L����ݺ!��=�'`��<
��Q���@��=.$YE~��Q0�?����'uYl�!¦ -{���N^S��O���Y$V:5q�M	�^T�\@`ǂ+=�~B���K �Ҵ<�Tpjq�H�z�<��W����T$Sb�m������Y�Sßl��{7RAV Q,~o���B�Gf�@���iW�M�������|rI�	���h���2V�
̓��
���0W���WjS�o;����S�s�X��uf�5#JiPv��6T#��2����I�����~�����Q��&*�N=jE������ğ���	&o)�|p��8Oei�eH�h�Z�I� :b���ٴ�?��$�ڣh�ࠣ���6�:]Rq�0J��D�O,�B��mZ����	ɟ �'՛��J�_/��H�� ���ï��x*t���S�����S����L?Q ��� �"���#$;����5��P���\�uo�$�Sb��3[�t:P����4n(�'-z�9܎R�J�ȡ��	H+Ԣߦ��I�8��	�MS�'�?i���?���M2��6��	;S��y��c�S�<1t�+<���eCD%B>�|;u�P?���i�J6�'��[��[�P�q�0jކũ@�(-(u��B��4�?���?1)O����O��Ӝ0MJ7�@"!����$,�nd��,>a�㌚�?ѡ(� .q�)S�j�}:�Ȃ��=�O�K�i�	���1[��JS��5x���H/9$�<�5��=Q5�h�E�'�ȩ�Pa7D�`��i a�4aR�&�ְ�Q"(}�K!�ɬ0@�Zش�?����M��JM�Bc|�[� A�K���	�����	П�ja)����<�;|�E���_%"����gG�"��dD~��_��H�8����.I �\`C���r���6�	m�~�d!��`�A8�+އ4�H�!�K�>q�C�	
�z�J�Q����I-R����d�N?i%8hD$���eɰC�.�hbLGx�$[�*�Y�'t2��d�'A�fj�&�
��r-FU>	:�D�=o����R��� �A�3^X�����ʧ��'k��D�g��'2�X�`ݎZ���'��A8���2�6��"�/j)Q?�0Cɿ&�L���Z�~WH��#�>�W*ߟ<�IR~J~«O���UO�8��J�n�){�DL��y��ܺyvYA�D�
m���yq����O2PD�����(���b���b�6���'��5�����OV��7y��o�ߟ��Iߟ��'t��)ȬI��AY��<hȪY��'S2��Z�Hņ�	�|vx1�3�1*�qZ�� �nТO�����'�� ǅ�N!�8 e
M� �.�K<I �۟t��I������<8�0d����B�n4�-�F�N���؉i�����HO>eB��qnYI`�U�b� J�
K8e�^$ߴ�?!���?�/O����OJ�S�jCZ7���1���'t���� �_�B�a"��M�C�P,��p80G5M3x�łA؟l`f�.4J$gY�M�>ܨ���J���0q�fH<�Ai_1`�LC���F3@T@a^s�<I@(5 �kuJ�\���;ԅ�z��k�D�0�k�i��'��&T^���ˆ���5?�"4��s2`��?y��?% �?I�yZw*ް�F�U4X���,�9�1���M�p̑>��W�E3T�2(9I�fC���!7�B,����ԟd�Iğ�;t��x�ʀ?~���Ə�3�����?�����E�u�Ju�1dF+�&Uq�/�&G��~R&��D�d�Jo(h:0źz"-�BW��D^�7��lZ���Ix��ßDn�gT0ͻ!��d �lr��̀^`py�����E'J6P�ɧ��9�	^7S�yrnS�6q�0ͺN��ɄG�vű�lZ�)�g�? �����,����C��S�=��]�l��h�O��d�O���"ҧ0*�\��לs+�x��T6��i�OL��$lOFu:ƪNHv�E�"� HՄ���������1hR�ߊ!�8�e��Y�"��vɛß$�Iߟ(�QlJ��M���?�����wL�����YA�#H qu�!L<) �ʌz�nt��	��xƎ����pf K���'� Bѧ�Ԥ���	4^XMa�"Ǉw�Xi�4��8��p`���?Y窕��?��S�Y���ݦ����p�����F����?D�8��ؤwl�\�&E�%��b��@���4���$�<lX� �xt��!ל&��1J��^�x��"�i���'�^���	ٟ�'$�4�l����kX�r^j<i�)�
2l���N6P��n�����QA]��������6ϰ?�	�զy�p�̭S��kAB��p yy!��7��x�,��6��A��gS�0qc��A5�yb���}�4|���
�$���L٫��I��p>)d�D[$�Xッ�hN�)`7�F�<q�D�!��D�ck��r�RE�ȑ8��c�MO.Z��Q2�ł�@���-C4gc�U� !�x�(Q��X
�!�¿\����G�
��Ȕ�,x�!�Ę�D�vP�,��,��4iV`��$�!�D	
,�����l�4m$`!�$H[K�ԙ�n�t����m*�!��5�V��k�KR�A4���!��
wT$R�Cʹ<����C�r�!���[�hqy1���  �p���<%�!��0k�����B-{4t�2ddܼu�!�D363��UAW�����Ƥ.q!�d��1-~�XA�_�O	tPC7A kO!�D��i&�xd�ק8���@��#H�!�E<�"`�D *_Zi�с�E�!�������H�kN��!6雕S�!���4!�	�.�pG~T�"���!�D <j#��]88�U���F.�!�#2�*2W���3�K��-�!�DG�\������9�wj�2�!�I���R���wx0�B��]�Y�!���I��1p�%X:(z,\T	�<QE!�$�	9[fd�`+T rVq"�ٗJ!���=��FD�1AZ��c�UO!����u�U�@�mIʽ�:2!�$�0g��P��+a&(�QKC!�D��~dl]
��I�!���*O"!��<A�\!��*baX3Ț�!��	.�ꥹ��͟V pCp���P!�%Z��r�nM7B�;va�!�$��U}C�/�9��{�F�]�!��Z�FT�p���U��%ɷΊ�1�!����t!ATgv�K-�\!�$�0M�H]J�N�2D�a�Mƾ0]!��G�z�n�B��+R$%� �-7!�$��@�|	�P�K�cs,Pd��!��� ~Y椃F;QT��&J�VW!�\7d�fq
ե�jS�Q�C�R!�_�4Gʅ�R�"SB޹臂�!�9�H�s��k?L�t�H@!�䒻?w���<����,-!���VpqɁcǜ(���g�,	!�d
��ʸ��E�`�el��;!�d&T�X!�PCZ+�j�q�&�![�!�>�� +&�S�~%�dI;N!�ę�.���-�
%�|9A�ā"!��`�r���7�.�`��Y6~ !�$�����E#^�b�=!,�c!�F�-��Y(3�À=�HKA���!�� �`�D`i��!�gX00V�2�"OUS�BE��I�,�1 �Q�p"O��1��f���V�����"O��`lʡ&���Ö�?(����B"O�]�7�,U��B���0Uʆ���"O��ہ�[E�5HюU/��c�"O�I��J׀cǨ�"�$0��3"O���Ä�h���c�L��;��b�"Od1БP&O�\��jJ"��Y�"O����ũ|k0!@�I�\��h6"O�Ai�̭m8�mR�#����"OX��CJS�n|�"DJ=<���Q"O���߃�	���K��A�1"O���3K�"��X���<.��2�"O�l�"�.(<�Q�D ��!�"O��T@˘G�j��&���Q�"OX%��+L4Q�^��Ԧ� �:1�!�I+D�z#~b��Y"`#0XЃ%	�9᪑PQ�S�<ŀE�&0� x��C�Ќr��U@�<�D�6=ZuClW'T�(���hOC�<q�DS,���7��#	�I:s�UV�<I�l��b�� CQ�r�r śi�<1�*g8D�걁Q-)��3�FY�<#�O8,Pp���_Mb���.�Y�&��zrNI,i��%`Ix29�#���xbniӸtȠ�Lҵa��W�<�q��'Bh*��MKܓ�li'�Ġ3�(��E@��n���EB�=ڧ	
��)�$D�H���o\�-�`�'�a
�
�ptɧ(��1���e0�aD%�5z�U;��'�,h���
F�	�ӲXJ6dVt�L����ٳG��tym�eBfQQ���)�!K4(,Fx�jQ�'���+0d�32���pn���f,n�1�r�~�P�ـ,�])��(������G	����k�L�B)�hiv�8����c�	Pԅ�v�B/M�Ȣ���+%����>�e�˸T	Fn讴3�m��X�4��%9WN ;��l" 3a�S�yf�!��0f�n��>�%�~���X5;��7sM޼�ӊ���%���T�s�Ycwd(<���QKސ@��>���bkNXJ��x)2�k4c�]��I
	�DEV�+Q�!���'���HċSJ3���N/P���8�P�8�Đ25�ъ4BD	�������'y�l���50�� ��NL6Pc�Od\)�D (��x�N��'/��D�6���hq�ّl^������W���SW��*��];`JZ����=����o~BDӟ	PB�2g��4o��ku�N
	C>��'�(��6�Ԋ<':�4����p-��o�V��#����'`L3WV`reF��i4Yq�%!�O^yiP��5���r�X�kVp�O0�X � (�.����aā��3񏄲��(�2(�I�'X��x���0��Ԥ�wx���w��⟼���Ӟ!�}8�i	C��I�L�l��c�P�$ƮXZ1�ؓ)V,0WM�*9� uH",J$D�)�� �r�h���%��O��q�@2[�&�)&G .M.}w=O4�e,ӝgz�����W?i޴Y�,�96�OL*m9'�ͨй7���[�|�g� T�Jj��'��(��hG/{qa|�>O�\}(��Ŝ1f<Q�/�
d����-�iC��~,R({�K'B�<ر�N�5�� ��������<-jI@�6�` ��Lf�'a0�r�}RO͙I���J1B�G�� ����x���ō�v&�1�'.�y�SJ�5n
ґD�G�4~�Z���"Ψ&� �H���?鷌�Hܓ<��3�E'tB˓0O����Ѐ<dD��7@ܤ}٠bU�:%�#&�O�1�F/'���5��		Լ��7Oh�r���_�Fp�(OzX�q� 
icf�;I~z��/gK�� lD�R�������Ă�o�������a��\��O@�����/�((��Gۜ|����uw̃1Zr���wP��Y�.�+Gfx� ⓷Hڄ��):O^=:�8?�$�Z7�: �C�ʋO���D���=>�슣���&sh���5��O ���cx�����>{�Z��x¡��$оg�r��M?�b�@�!��!i�!�?$��(�oY9;|n�+u�Y��"���Me� ��/���b휁fc��;��O�4⤉@?�'bb�H�8H`���/( �Nm���I{�O�N���̩=�):g,�H���h޴p_6�m�o�����Rr���"6p�ɺ$$��8ꓦhO���,KC�z�n�"E�cX<�#���Q�Fe��X_�t�Ҩ��,��
��X,E$4($�,��E%6,Dxʟ� �9�R��.���P�JL�^�8�0*O2�B��`?vmك-��`�
�Q���41qOȠ��!��
c?��
j�q�E�l~��s6�0�ax��l y�E ^�]]�(���L8c��,�6��6Y�%��*}���1�ŕ��m&P���@�8Lx"f����'r"=E����.%Zf�rcR��,l��Z>�y�%�"0(Y 	�=�y���
�|XS�Y�?�n�c0o��<�e�}���<�%�,r4�0��QwBP�JAp��B�$Ք*c�'CR�ڒKpB�d�Eȑ`p�L	D�6-���7�x2(��iWj9�����O�W#�	]�Z�&�6d>�<�� S�ay���O~b�<K�'����@jPgD �l�s��U�v{rdz�+̧pN��'���Q	�,7��ɟ�dF�Y�͜H�"����'�#6�$��8� 8���'0n�`�4\���P�bͮH��'�#U���d.�Ī� �p(B�@�(QS����E���Bٻw�r=	D���#���u�V�ZR�k���' +��+GjE�$AS@ꌌ>�N9Ԏ_�)�\�2��x�/��cv�I"�?��:ō�#���g�%"����.R�$6��O�6M�~n6j��+K�u���І}�Ҁ�-2����dc�j���%�΄�r�6U�J��a-��9"� �$cL)+��U;e�Һ��3�OHQ����q-�ݘ�m̜DL�W�2�o��`�jqKZ2���D|�j�O�����؍P$za��V0��-�T-|ZT��z����$�U������&u�ؓ��^&8���'�V~�)���A�+�@������e�d����^�~�ik^�s�VJt�)!�@(�J����F\:��w �CE�Ճէ-Mf���Yr"�'�2"}�'��B�`�	~�
�����*a�.4  �����h�!C�W�0} ��	#�g(>���+�F��b�kȱsۛƌE1�`���� rx�d��,�8X	j��4�$�!�Y�qbM�#%�#p&��CH��a�=1�i�}�(�@+�O6�r#�L,
�2����ޔ
�����'edA ��׬Z��h�EѴZ�r��3c�R�֘���U"T�b"΁H2qO%��g�'�ʄr��IM�L��L�`\�}�d%Z�" L���8u��
,D�F�&��0i\+�����ί̆s�b��,���9�KJ�=��̺`��1��	�H��ɴ*<�q�`ңH��" N�/j�`�Ñ"6%R�$L ,�<�2F+�@�)%���.[�yb�5��"L�7�ı]��M���O��<���0/�:� ��E�P٪M���qsXx�B��W�J(Z��:��X�{���}{�����[֟xjg� �pBܭ:B%S/���8O�Q�*�<|�X� Ҁڑ`��+��/� ��WG� :6D��윃��'<��[��>;_?��E��IjD�F
B���#��6}b�ԄZ:��yƄگW�di�c	M�Oٌ�bp��}i�iB -�*��!��H/e|%�=E��'A�`h�B���{G	��#��=r�5&0��a���� "��""C�hx��B��'����l/F�3v�[�%��y˅�K�,ּC≋P8f����:%��RëNm;�!z�#�;�~�(�_w`�X�l�����'D��b�G���CƬ+1��#��Er�><OĨ;��!��Uj�G���M[�� |bdQ��ݖy��fcS�<ɷ�Ɨfy�q��
1��<1͝9*MD�E��:e�q����s�2�HPҌوh���;a�Q�0�X1�ЉkP�U��ԥ�����桘�g_���x�a��_b���eµwǆ=P��C Z���u &�$��.��3K��t���j��G}N�(5b	�7_�y�G�7iC�	 -�愓p]�WJ`=sa��]V���/O��e+դVCy��9O�ș֨U%;�dµ�F�(��%v"O�x0)��,�n�J�#�0 �19O�4�v-���G� �4��Ϭ�&iqc-ӏ|�:!K��;�a|�ٳ[=��tgWK��8p��2P*X�	p/��d�kh<��N?8z<�����|�0��k�c�'rvB�]�}w�l���H
`�R�J]�Z�H��f��d!����\R� 70�4�`5�Q8d�Po��7x`S�>E���Iv����ý5�c@EȲ;YR��6	�)"%f9\��0C�+��N��'���Ǚ_��z�Ә:q�9d%.RL�`�5�E�y"J� RX�
��S�=��I�
W��yF
�`@�ȤL!��X�t��y��,dƄ)�e�HG�$�[�X��yr�Ɗ~��MjVe�l�"�d!�?�y����\T�=���[k�1��L�y�j�2��ڱ���;|��R��	�y҈��6 ��(��/4E�LY��y�(ܹA� �z6)D#Ǔ�!�� 6%�GY.S�Tx�f��=I�| �"O���5��?�v�� ��O7 ���"O���sfO�x)�`-�] �2"OFL�r�N�С��kûotQ�$"OJ� C�H������J_(w�*Yz�"O�dᔯЃ[��0K�hW-2��h�"O:la�i��2���h�0t9�"O\���$��8��8�EG4R l���"OU�2M��Lap矗r#����"O�(�玌�Z�JT��h��Q/F}B�"O>���U*�<cF�B�u��9g"Oh�s��EZ��GG*��q �"OV,Y�eK=�ڼ�B]�8Q2"O�ŀ�7�dY��h1	�)��"Ox�9 �Ǜ,`�(��X����V"O`���I͢Tՠ�*�'M7��q �"O��,��U�	��hL����"O��Rf)�?*�\�Q�o��+s"O��!@�#�°睯0#Ҩ��"O��Àa@�:	�\�5,�f�5�"O�p(��A�peТM0B�'W�����F�T �!�:4Ӝ=��@/��F�ݎ��- �ev�<�P�Z3/�ް���H��	 ���r�<I�I��^�,x�dE�pp4T���j�<����)A`�I"�\��d�	G.}�<Y�e�")W�(�D(Y�JT@�	$@w�<��ԲC�lz�+ȋ<6bݐ'�u�<�P�]��T|y���r��&�W�<q2�G���;7�oƮ%�#�V�<Q�拉x�~L�2��6��w��{�<�r��4�`���_HId�O�<qC�.^%��rA�ӄ	���##r�<�25w�Nx�`Xǆ|r��[n�<�U/�=�,���ZSڱ�b�\^�<9��F,u��������nf5âo�A�<�7�A�<K�l�"́���2A�w�<�E����\�Ӎ���T�	v�<��mδ2J֥���A ��y��DW�<�G�U�:��EH�JK)�HI��� Q�<Ѥi��y�	9gKùwr@a"##Qe�<��/k�@UFR!R�ԕ	q�Y�<�榚* B`�p�~�U���9T����;A���P��ʒe����N7D�$����0hj�@�t'H�I���b��3D��y6��(�V�#!��p�U��(2D��ǯO7־yRࣆ�z@�`1��<D�j�eL��H��ڷ�T�� D�4X �x��Cw�_Z(m�2D�$9�o��� Cb*� .&��sa�.D�AR��vr�Q��Ն3����-D�h���){y(
G��)2~Z�;b�,D�P)A��8��hÃ��V��a��+D���t�������t�@wh)D��:E#��pĢ��]�pè�{��*D���3��$M���(�F%O����l5D�����,W���ĭ3�VQ�H3D�p�F�HZ���b �^��9��%D�D*�$�9���G�_�>�HD�(D���2�4TFL���[=~�Ñ(D�̐���FI��yөX�Q���;��'D����Ӯ3(� v�V� (�y�%D�xIZj$|jA�d���2�#n�!򤛌Q a�`FZ��E�&���A�!�$Kwg"p2AEO���I@�(���!�� "�30)���(��.����"G"O8�؇�(CVF,zBn�2%jH�qd"O��K�%	�.�n��-TXA�F"O�|9bԕ8�x�"�L���F��u"O�5��b2y`<�D�V2�����"OJ�
1Ð�d+D8�B�8`�	H7"O>R��ۻ>���  � Hh�"O@)��X��e�0�Ddn���"Oh���/
�\D��Z�n��"���
 "Ox-���?f���⇚[r����"O�!Qh=E�l���B@�U�� $"OB-C$�W�q����cV�Ufya7�'�
�@�-���}��F�S�N�J�I��6�|B�ɓ2�m{�@C��: �@eP0P�f�|�U@4�+�)§X�4HS�L70Ldl8�b	�B�8Q�ȓ.T�0�����M0�h�D�!�RE�<)4D�%�B�񤇲1�*Lो� �(�$�J��!𤆰5�p���Ӑӥ�Ё�,����Sa��L�r*�	���ݎgE��0˕>#��`��I=s3�5!�{RCU(�h)�l�m`����H��y��YR0��ەi�ҥ!gn���yBǺUW&q��*
|�4P�Ś�y2�Y{��%R @M���Hzc����y��S�����D+V2�b�LU��y��3ؘ�GȊ ��QB�͓��y�G�>i<T����L�NA!� ���yrnJ' S|(���[�m��st���y��L'V_��@����B��.��c	�'?@���Ť^�a�*ѿ7�d!	�'�p��G�Ùu���Ve�4[ ��'O,�'�B�r8ҁ��M0%[��#
�'I���&�C�r�,y��(�f�0 ��'´3��'G6�
��
�7٠�@N[�z� �'�ў�'=q|訩O$��/�:���R�c�4���"O�x$FD1�ة�N\~َ�A�P���O� 3�h�q���	�Fդ0bz��r�Rb4Ǎ�A �s�E��[{)	�*y8��{�,�Ld�s烈�}R �&n�H���b%֬=�ȻQ'*b��c�l[l�b�Hԋ��_��3�	p��[p"�.&f@rJ�#GSx㟈x�`J`.5ӳ�T��>�����':%�F
P��H�:zAr�k@o�p�A"���az��HU�%�"�5;!P�e�<=��p�P�O�jrXPQ�K "�M���/�ɶ���N�iE�(��c�==ZD(�-�J�!�D'�)r�ǒ�
��yѥ�l.azb�H�&o��PgWZ��:��r��(��ȃ^���O�ǰ<Q�ˁ'm����Q��"4�G��t��$h���5>(����+�1O(����A}(�H`Z�vZxlR��d�$!�����;��i�ä�&&|�'�\�B�Y���͘ �y|�C�}BB�i΄� j�Z��dCY�b�����\L"Fi���E�0=)�펳M�  #E��'QXB`c��ĐRZ�9ٰ�x	ߓ?T%ٗ��iz=�A�ڑt����G�@r���ܚi~��h�A�[����Ra|�$�"M���f��L]��D,t�Z��k�;L>�8i	�P1�ih_�Yn0�R��ע��S�^�s��H(!!��i�1�ɠz��4����2gv�TJ���'����B͉�l�ʰp��8�޵�O��c5�\p�iqGǾШ8ӐE,���\�	��悋lی@��Z�}C����X�.�ʲ��k��$�3�'y��2��	�8J`��KE0%��/��a��R���D��{T.�0D�Q`��F�ѐ4@��T!U�$Ⱥ6l�[A�yWg�q�ȈSۓvo��'�91�\H�q�J +d�8�T�6�VjV��@��x�,C@���YU�I5F� ���|�%��ĝ"h�A2B��HR�i�<A6J����h�#c@�H݋%�Vx�~Ԓd���Ŭ���Y�kY�)�1�O��!��ǒxӘ`��J��X�����ǞF����<�Ր�V�l_<�o�1:���A3m����'Z �i���"#�J�1�*�m�4���R�f;�,0���8s/�zZc���(��&�=�2�9$�|�
�'��qy'k��A=��5�ǻ@����j�n~�j�s�qO��1�כ v���b��72&تufڻH��Č����h��',�� 6n�C�a�N�禼� ����	�;FOPV�T�=����>9����,��T34NU�~�2 z���`��.r
��ϊu�������F�Xx�O\�Ӈ��ox���M^bc�[��|RM_f��E�R��-p��)��@�'�T� L�h^���L��0>I�/�nZ�Z f�>T�]�ꘂT|B]"宕�E�V���p*�(J�V�J�,O��8�=Hw!�	ɸ��a�M2�eQa
O��$î?!L�iD\-C/�,�Ħ��fB0���'\��rtR���i&�5����Wۖx`�LL�|�c�^�_#��ÓG�=l���;&P8���_>Ew��0������Sc�$D=��ks�T��CNM38�$}��C1I
d`�5�Wh��Ң=�D¬&�I�Dԝ��{Ħ�D≈{��3�]�I��I����I�������K�Z�"���bD�T��,.�Lq��E�p?7Æ�_���ra-�m��%�!CɈ1�ly���	WV�iҒ�OR}b���'\����;f�J�FjǩV�B�
��Q:9Ҁ�Ɠ!�~4�㉜�9N �S�ٛ"n�5�C�O#��I�"M�sǥ�>"����@�ȼ� ��B���n�X� k�6HKp��3);<OX�"c��p��7!$m��)7 ]�?3Ɣ㴤��hNŊ���2�R���oU*��9�>)�kި\���<S��@`���5>�� ��Tf��~���"��D�q�*-2,�~��\���<2��d�<��H��"./�̲�%	�I����/O���˛� HazB�ktz�:�6Pl�!�U*��Th��B����``��"{咩IG�8��T?�h@TF<PxksΘ:=G�����!U�	��D�<��)5��J��)	d�܃��Տ�bQr3�Q�dB��(^���g!S���H���	��䞇8T`� �Q#�98�&E�n��љu"O켒,̸y�6�0��CC+�Ujf��IR��f�;'c�%2�J�<	5bF�-挬�<�"�I�$(��E�t�ԓ�jGV8����H�'�P<�TCF�}ٶI��inV�aG.
$G�pc�F2#d.˓,4�<IC�Xz���K%�əv�R�:�Ɨ �����ɶ<IE�z��!	�;(�Hqv��٦�?y"�C�
ɂ`�`m��Q���'�.D��� �M5\�A�͔� 98͘��S�q����R��;$[L�
��˼Y��L�$��!��T��R]�w�*8����>�O�"ǁ��ؠ�4˘�O
�hE�ġz���s�:*sx��4Z-h�����>��FH�+�z�ⵧ��џ��R@�+A�.���Ϯr����t�Vz`k�}�	�M�Y�C�I%2$L���O\��i@Oˢm�|�Lx0CՌ��%:��B���:�L�g�7N�4x��K�puRC�ɚ���b@`7m ^9����A��j6�Y}����UN������{���l� �:���"C *��?A���6���p�*L�,��3f��,X�P�R>o���(52y��'LqvB�����
���ÓSJĵ�"B,P�Ic� �Q���+�4!j��=ps��
4��x�N�r��)�@��{������Y!���؝m62����%}"h��c>�{0?��a7.	��,X�h2D�ࡐf�H��R�	*Z"�K����'D�H��:G�R�> ����Ë+�� vF����5�8�p��*~SLI[�E�9p�&�է�(��y��ԥ�p<!�,�o�bdk%HJ�s��<K��Uvx�di#��p���r�E'�^Pp�ɛ!�!��$e������͕S-�����V�ee�'���Ey���* �2�P&��[[>���$��y�#�
��8! �!P.���a�/�y�BL#UO���⁙J;@Æ�N��y���|��ˤ`�-�Dx3O���M����y���1�x���i�P��wk�8<MH�aBP�Z�:q�'<H��u�y�r�qPCO*]�h\��X��㍁rB�z��'�b5�M�,��Y��}���'�}��R�\E��K��\�!�̌
P\�-��EUih<YE���%{�Ԓ�k̒N�����g�'M,��CFɐ9qz���4��)���ʧ�%hD�a��c�<1����� �Ph�9��i �`��q�	"�F@�K<E�D�����
D�7PMs��0�!�dE+��`(؃C���� m�!��4?�>�+�Ɓ�u␥� ��i!���4-�$[�nۙ`ɂ`����,�!�$˲D��0�J�5Y@ �'b�!��̀���� ��쐕��e� 9�!򄙱-N$��e,�|���8�O!/�!�� @��g,΃҈��h3�0��D"O��ŏ�>n��y��~���c�"O�܉s
V�B�.�0���jӼ�*�"O�l��i\�-�4X1��T�hĔ�ID"O��Q�����U�`_�Z�ܘ�"O(-�d��RMz ��	)h�*�r�"O�PpD0�|�`��8�n��c"Ob-P��V*+c�X�L���"O��f�9TQr�Y��20`U��"O�m�`F;ArP�+��&�E"Ot�x1kZ�
cfY�R+�?�tRF"OС񤤆�:���XP+Z^$[�"Oʔ�5����APu+�#Iq�"ON�c���6�6��	 �l��"O0Q��S�����V��(O��p1�"O(����(H�$T)g�A�-z�T�E"O��kv �>e^�{ �ۑ	m�(0R"O�=�w�T���!ӌ	
Z�BIa�"O�Q0b	3�:�ؑ�T%�D�4"O>@�nI�-A"]#�ɟ�΀��S"O�s�����j��Խs����"O��Xvʍ1Xtz��<!�r]@6"O2$ѷ��
a�m�d�͜����"O�@���)� S$풬)����e"O���׆Y<�a@��R��H
p"O*	a���)2��Q�7}�=�1"O��("�@1fH���E�(x�p{�"O�H���Pp��1-ΑUe�,��"O`�b�	.�.};S�E�JT8a��"O��᳆I�	fqA7 �7*W(�X�"O�%���o	x�BQ4/�.�K�"O�J���#������#BF��"O��*���o���rSY����2"O�,���r�����kےa�4�H�"O.!�1��/�(U2�J��t�h99W"Ot�0E��4'�D聿�^�"O���!L
0��=8u�_9"�T8��"O�a%�,Z�.%�;R�l���"OH��c���]o������|@"OpE8��]�����5���0�*hZg"O:=�d�^7~kȀ��Q$�$�Z�"O&k�OT�bT(9����Y�̭��"O¼��(.8`x�S�ʗQ��(P$"O��X� E	X�2�peV $���:�"O�H�P�E}f�q�c�g�l���"O�B�m@�+=�a��G(�*���"O��:@:}t�e
7�KF��1!"OFl��nH�\@SScӍ0��5"O�Hy'�Z�	d�����M-�X	�"O�|Xd�	��i�V?#�b�)"O0!��	��>GnH9CƔ���(�"O��.\	T�,<#gd�>�Xٵ"O���g��� �$��r�zU�W"O�Ͱ -�s8t8�▕mҞ�E"O�cg�В$�o�{�da�"O�}�cG<�bwѨi����U"O�B�	K�Qά<�Y��nR"O2E�T�VJF�{T���1�|��!"O���b@���s�Ά�=��[�"O�p�+^-AnPc��� q�D��"O���F�@�|�DB��ԩ.U���0"O�ƀA%��|BX�f-����"O�9[�i�V���C��M�c����"O*t�t �?J�ԁS����l]0"O� (Mb�/5wʔ܂���z���S"O^@2��4X�`Q�+ގpm��;�"ON�4��:�z���`[<7��J�"Ot��� O������:7�L͑q"O�K�|(iɐ$�%#��HH%"Ox��rk� i:�t�c�P�D�fP�"O܁S��E枽��C��F��"O��k�E��J�DH�웝:�`���"Oz��!�*<�������7�,�Q�"Oz<�1�A�fdk�qzV���y2m :�T�`iC�ET�1�NO/�y�DH0l�y@��E��iA���
�y2	��z��IFIŢ�<�	�a���y��$B�
P��	��d*k���y�o��l1� ���	��	.Y((1��S�����c�d�% 1	Ě<Y��ȓy���B2*��ˀu�7�F�ȓx������ĮbX��;e�ύ�����0����č16�0ek��S�y��9�ȓ!�R\���ܼ	��`��
�jr���VƐ�%F�n��ˢ�@'}�&��ȓ_G��A^8LKh�g���k��l�ȓK���3��_�5`xdP��
�J��ȓ��`��l���N9x"�H�0��>�����ڲgUzܫ G&D�ȓ�f�  >f�F�.hl������SW��9�|˔N�+/rt��#����)71�C�(=�f�ȓt`�SЏԬG.<͂�o�(4;&��ȓ7�@`�L-��*gk 1�nM��+�T(F�ͅ6�`�"��9Pp4�ȓI���#@�
&�:��נ7e\���R|H	�H�T۸$���	'k`j��ȓa��{f�V��AQ�V:Cḵ�ȓQ-�����o�����2T����ȓW�`̺B-J�sE!\�pW8�y�dK��l�x,�|F ��u
��yRN�J,���[�}�>���y��)W����[w��t���:�y���C&�ؤ���y (�!��T�y!�!ظ��C�o�Hٲpǟ�y",�+{jXM�N��[�|K%���y2���Y[�k���d�j]r2���K	�jS�+~��G`ˏT~B��ȓC����!F�cm�e8��
D�~q��4�y����XhXt�*m��ȓ"A(��)�2`���'�:Z�,������f̍V�2�CC�1#���B��]�q&��sMR��gc��$���	6���(X�@��RB�H!�L��r4L=�C�.z����p���w�y��IɔA��ׄn����S)�Vԅȓw���"����Z.1��p��)��Tz�R�`]'|̂���ID5M&��ȓCq>"r�E� ��d���I.H��ȓ$G���3.��7�Zh�Eӄd��Ʉ�7"�P!���:X��:�N�����%,:i�,M�|L��Z�r��(��%�<����L<n�4R��0LuJ�ȓu��	*�ʽ}��� f�#����,�<�9��P�d&<����L��<NP2�i;uRd��']
��=�ȓ.6A`N�=h��&�J ����o.��g�Oa��������9,
5��S�? ���� X�4��5v~�p"O� ���?����Y =(�aas"O����kn$A��7	���)�"O����%�S����b��-?��a"O�]��@˃G��@BeLE�"�B"O&�"�j��86��6�þS2<K�"O��Y ��4ӘU��F��֤Х"O�!�@� c�lЃ��3C�L�R"O���ĜPv 5#��E/��ȳ"OHQ�̝��&���a�X���&"O�bU��(b`D�( ���`�R�"O��� �!�P�8���l=��{�"O�ӷ��$Y���ȅԹ�"O��iߞ1𚌸�.�j�6���"OTI��b Nԣ�m��
�"O|I���l$�L�I�"O��C���,7`���IW�^`�=��"O��b٧C&��造qU$\r"O|@�NX���r�]4�d`"7"O
��dM�颽��g�aI�}�!�Dڏk�\�Dhθw*��IQI�(�!�d Iu݀��I� ��(˴ʞ�$�!�E�PNl�j�	QF�:��X�!�T*%�ʉ2��C�TC�yГǓ�n�!�䉠9I�Ea�X,}��@KD�=~�!�O�_O,e�"�:wnSEe��?t!�d<}���4E�;ezF�q6��~q!�V�r�:� ��_�,�e+��[m!�dX�FhV|���GN��		�MR!�$�S�hi�CbZ=:0�!+f�T� 6!�$v�p���AJ�$x��<!!��Q�.N`�K�bPoQ���ѭҼ{�!�$�G�$�iĈ�M����,*O�!�D[�&y.u2F�'7��W˄�;�a}2�>��Eˇ��5#g��!��9��|�<�����5F )srB1� (��`x�<	���j̈�Q��ՁX�
�`�c�M�<)A�	���X(G�O�J]Z1x���m�<9��)N�4y��O�j��]�G�l�<���Q�1�#�O�x��AXb�<�2���0r#NZ+E�� �F�_�<y��3� �
�k��bU-�^�<�*ЂZ<B�a7.� -��x�!C�R�<!7�M���v�	?g�
 ��I�S�<��+Z0���8nƾ*J��C��K�<��O<
��x��!�<5?��y�#MK�<AQ�V�>�J�:RƜ�[ި���"Sm�<1���D~v	���h��:�!D�<�u䒫[���ʹʨU�T�|�<�����iǪ�/8�\xᲮ�w�<!F�/D=pBدE\��0M�q�<�s��'�P�T�-PF�PA�)�G�<�W���qئ5`�C�'1���W��N�<��݅w�V���f�$$v$]+@C�_�<ф�	 �*uš	$,w\$s� �Y�<Aw�N*i�T��F��:+ިh�Q|�<�F�M�R�����%@��0��x�<A��$$5���Q
F��ș�D_�<�ta>Kmf��T+
r%0�eMO�<ׯ	o&X���W�~�4a�&��I�<	2D0bɔ�a�`�1
N:��f��A�<q%��2�N�)0�E&g��De�F�<ـ�ί%�F(�4�.I�؜� W�<���]�5�y��cޫR�lQy3P�<� ����BP2N  �bfc�(\K�0	R"O�0�SŒ
D�޹��!W0��a�"O�\Y�a[�Z���A!��ʒ"O0dh�)JW�L!������P"O�����S)��A���$=��]�e"O:�h�a�2�HU ��w�f<K�"O-�0���H�ҕ
է
�.$��"Ou�F�Ϧ9k��s�Ѵ+H��z&"O4�耝>���wd��S5<d�U"OZ��RD�6L�5X�LM�	4�SC"O�9�D�=<�r0��](��kV"O���O�~�6t+n:�M
�"O�����gX��a�$�3���`"Oބ�vj^9\�R�D)ontQu"O>��$�]�"Y�����`�:q"O��+$N�{bu�����;_(y�Q"ONXN��^.���&B�(PH��"O��y�!��H��ӁcCؚ9x "O��Qԭj�Ԭ8+Ɨal�x��+D�IF�׸E�VИ�.�-@���s�D)D�ĩa�<�lk��e���$.=D���ӡG �LEi�g9$|A��O-D�`Y�Lݧ_B���׈Oْ�AB(*D�t0dĐ<�ސ@�	E�&-)Ԧ'D�4 �%Q����e�F$8���C&D�Q��5�>`�Gf�>o��Xa�%2D�P�U" 5(�T;��	%����¥.D�,��D6'O�����K��;r�+D��r��e���C��x���!��6D�����F�@\���5)T(}�8D�C� D�����Ż0�P�a��R�?f41��>D� iS�!�ʍ���T�|��I��<D��j��u XI��ӱnr�a!j9D��j�q�H���R���Ů+D��B�懂mq�x�r�O�BFeb�.D���`�ڶ�X��#i%Vt鳄F(D� C,�<u�l�Ã	�HǸ��6H(D�X�M���I��2_B��r+%D��(��:~�L�oƕh�b�*A*$D��yu�=�,��B�5IY|��t@&D���t!Oa�U؆�_:2m^��@�8D�4:E��
%k�����݉h�z���C6D�P�unD�RD��e��F�>���3D���Uj��H*�3�c(	�j�" �7D�((�&��	�� ʺb�:-ڀ�4D��� M6G�xs�5$"6!�2N-D�@4k/E�B9�S�j6� �&!D����E#Ub��c'@C*c] �A��1D���!*d���oN�o��!��(0D����䆕�
��cB�>d���J"D�L��mJ0�lI ���2�L�˶K+D�(�D����Q���"b�9i�E?D�²�΂xgԉY��	B����@9D��xCIA
 �j�Qb�� '��ht�:D�4���܂E� f��tZmb�"4D�pq�X
�h�S�ɮ���,0D��1��ܫnP8s�(�x�y��9D����!�w���
AR�����J7D�x���&��-K%��:�pIС�5D�p��Ԡ}��bY�Sfe��O'D�P�V}�	�%[�H�(�q �*D���4�h�Mj�������(D��q��Z2������:����G�+D��)'KQ_F�Ыr��S�L�)D�� ��c��F�%��,Pv�	"���[v"O��X��=���2��f��5d"O~�I��Th�bA.K�dt�"O�	J�J4<\���J"p�:4�P"O��x�	�%�N�{��P&(!��p�"O�9pd*��*��`��z<=�"O��Te�wd����F��\�
S"O���q�:5�%X�&��Q�"O����E,\0��*�;OW�[�"O�A�E�@��9�%c�.r<�(�p"Ob�Ip⍢|H�!HW��< �Y��"O�<Sw�2@�ZS��R�L�(�"O���Q��)0,+�M�	<g�� �"Oz��$Ё���b,	�`e`'"O�s����̹g#֦4j��:�"O��p��ğf�$"�˄lT�Ԑ�"O� �ʙ0���������"O�u:Ӈ��	�>p�!,�b�:��"O��p�-T�\ς�
g��?Co�T�`"O<Ar�ZQ ��%FGn�,�Q6�'�Ope0n�T+��s�%܏]��8��"O�I�4b�<�ܣ�o�)F�
��q"O�a�!�<%��@PA�d���0�"O��$��w��1�ޖ�(���"O�`�.LY�NT8���;���a"O+e�U����\%��|��"O�%��4u�$ ����&-2p"O���P.x��RѨܮW��A A"Oƌ�1���B�i��F�:���y"O�ĘT��8hHT܉�˗�r�ؓ"O4M�䂈=�@�� KB�@ Ae"O�5sÎ-�2d�gHĜa��0�`"Od�x��م/��)q4%�<pu20�"O M,t��2	�{�vD���	4U!�j�2�zʃ�l����a���!��MLR�I��Q�H���j�H�t�!�%�����%T���X��+�!�d�b�5H��c��e9�Z�5q!��q<@�F�����pH�k�!�d؃�)Jw��{5b��4�F:T!�U�.~�$�kē+^�K��]�n�!�pQ����];(���C$g�!��7XnѢ.{BmRE$�3�!�D݀T�j�����ai�=�� �C�!򄕳N�,�Uk��xQ�1�f��LC�I��TE�WC�JFr�b�1+C�	�V�l!�Ul��xל�P���>o�*B�I?��5#Ӧ��%��5�t�D�S�JC�ɠ]��#MM�<�v]��+�	i�"C䉪2΢��S�&|��ަt�B�	
W(h@I5�
M�>a��Pi��B䉅4z�q0aJ�~x4g��AJB�ɹK@6ts0���G+�M��a\:Q B�ɢc�H�]�_/.� �Ǵ<3�C�� ��1���6q�h��1��XЦC�	"af�6>�01�'��4R�;B"O\i�ʟ}a7��7���>I
�&�R�AF��d��(A�ͻlʬ܆ȓkbP�S!ת6YD�0�A�7Eᢸ��p	HX���Y-�ň5J�E�����	Vy����� 
K�8��ȫ��Y��b7D�ȫd��Q�2���)�sfΕ�4��[���Oj��I䃐Fa|��R(U0�EK�':��ЃC:h�i+R�πljx
��� �ٰ��}c$��+�ܐa�"ODP��I�<qj�B�>"�䪶"O�Tre�Ke��96!����yy2"OH0"˾c�h!V:��1"O��6�G�2
ت�k05��ę�"O����:d��I�%�z��"OuZ�/�+)B�5�S�T�@��Hk�"O"�#�N�N?�B�+��Ʉu+R"O���%ś<���a��P}P�"O��"��t~l �� �5�2pS�"ON�vG���:� ��סh(NP��"O�Hs3�R�����ɍZ(����ibў"~n� \�љ�� 
�|���"8xC�	�	�ĩ)�H#1V�q!�"�&j�pC䉉u�\D�sjͰ%���	�	_�tPJ���2}R �)����̫����뉰�yrC�*�@�iЩ��Ȉ���y��R�/�({gٽO6����y� <z���I�$	u*8�fOF$�y��F>vX���� ��u��,˒	�y�_��0�o��j~����2�y��27ְ��V��<d35/P��y�-�1�tūZe�(�@T,T�5C�	�\�Ĵq�m�W4�i����A	�B�	]�
Y�vB �r �Y��&�vCC�I?�|�X�)�D*�����:F$�C�I!/���@/�QXY�'�(t��C�I8$om�q�R��V8\G�C䉣5����FL~\ca��F��C�ɩP�(h�ƖFu��!���VݬC��*0���1 �"24��3�(<�rC�	�L�	��]�;�EId�ջ>�C䉯c�r��/f4��d���.T�B��@�x���Ԝc��Yu)�8+�NB�Ik�����k�� B��P�J#D��kǧ��J~^
h�"��IR#"D���'�F�2ʄ��P�\,�ޑQ'�>D���s�y<̓�I�$T0���H>D�0�"c�F�-
U̘�a���V�;D���X:Z۞�6��[�ęSA�,��hO�S�R�ڭ�D��\�@E'O�B�	�J��� �*���%B�$"?I�����L-H����"E+&&�(e�!�d�K���-\�h��ī�B* ��D{��`�J��r[�l�%JC iG&c�'��H�$L�A�?V�����k֕�|���'����%���&��g M�/����'X8���?zܚ�6n�#��\3�'>9y*K ��Iqm$��,J�'�n0i7�N�#Z�(�l�q�\[�'�2IQ��[#$����ڎl�� 8�'`��S���p����C�پk��|��'`Z����(�츲��>di�!��'�`�xpf���zE�UD	US6X��'�l��#(� k*�	�&�0A�TH0�'=�E�a��V�h�� �݇��y�j�2E��j���.b���F�[�y��5��9�`O*:��Y�c엑�ybY�qą��F��>�yBAG/�� ��N�0��u�UI�+�y�  �t�G
��"B�X�,��'s�y��͆@�.Y ��h^5
�'��y�GK�8�<���3}/H�
�'� H��ĻB}�8q*;+�.����� REy4E=^��MCg��8&�h	�"O���3��x6���0&�b:�"Op�Zr��{��X�NվA����"O4��c�V�j��� �B�=B1�4iP"O��T"�k�&	J��X?�x�j�"OL��fE��n$��O�vݺ�"OikӀ^ r��`$�!]e�	i�"O>j恁`(�0�A��
M� �"O�T�E$�(?�ƥ	�0�8���"O��L�y�LLä�(,Ҿ�r"O��ڂϖ"T�Aq��!�>ȹ"O�x85'��R��ţc���ٱ(��yrnQx��G⟮\I�I���y"�Av�as�j��J�,D������y��	 �(5;7m�=_B���%��y���!f�"���/L�>}­D-�yB	��#��њP�O0d�-�D �y�.�-�bx˵W�l�{�D���y�Ģ00�0�	��T��(��yb��;V�R��g��� ��Ơ���y��,U��P UҖr�l;a/;�Py��5~ة:$M��&���0��p�<	A'�2+<�y�O�E�JБS�Hl�<y��}�ʙR��ǃB�lq��Ua�<q�$BDK8zS�cF�p�MI�<a`��n� A�'�)1/��BI�<)�kI�v��C�dF�.g�x;0�,T���q��2��u�b-�����$i8D��AaߢLV����+il&���5D�Dy�H
=V�#���g����K%D��$��5*V���f@�.�,S" D��KC(��#��P�$���	!M<D��Y�ǞT 䝱$�y�v�3�.��<i!+��zD�����W�>�4xe�Ht�<�bڼK-DM�a,R��o�l�<!���{��h�2@� Y>Uc��i�<T��	�����?X���Ik�<Q	��1�����=Pjܸ�AN�<q ��)̨��R ;gDԙP3�Pp�<y���'I�THӓ�:>��X0q#�o�<���XxA��	T�G�A`�(ZG�<Pן}�r�;'�̈́?�軇�}�<itdÀm�,�+�Ղ?;0�)�n�A�<�%�3u�f�Q`K̿Mw^�ф/�R�<q�+�W�D@���46̽�c�J�<����/&j��@.@�Y&����Fq�<	�j�1$�<�ퟲ/&�0�Tj�v�<��*L�}�q��h�.>�<�@�[�<���� gܺu��I�Gb
 #��S�<�r��1�t��w.ǳ���ʖɑi�<a��)~H��g�����&��f�<9-�=�qmC+y��Z�'z�<̚��Œ���*Z����A��u�<ٖ�>D|�)� ��-Vj�s`HY�<yqLR-DZ����Τ3�ΘSVE�o�<)V��e88-�pJą#`<���Ah�<��g[��p�*ف1S����Pb�<!�@Q>0����T$��
���dj�r�<��ʦox��R��7�Fc�t�<	�dGE��[ǆWM��E�
q�<A%-U'���Ҋ��8W|)+Cc�<q/$ �*-�VϜ8K��Wɐ_�<1׫�[[�AZwn�Z�Ezw�Pc�<�܋i��96� � e�4r���d�<� �适�;dGf);e��9o:�[�"O����0�(9)ޞ�$e�$"O���#������P�׸=N���"O&d ׇ��R��9)��ߨ4I�a�u"O���"�ƘN����B�\;R|�"O�a���N&y���bd���"O����O��D�R��CF�x ��f"O�Qs"�ED���D�vѸ�8"O���'D��3/ϣ3��a��"OJ��	0
�.��� �B�a��`�ȓX{�<iU-�*!��!Cq��1P_��ȓ���d�ʯl�H�r�/a��L��>��L#CN+G�̬�b._v���}�"m�G����0@�'�� �ȓ*G ͣ��U������,[7�u�ȓ/n�I1�*��RN���5�͏C�2l��QP(� �O1om`�
O�#�����B���h�J-��8���j�Ʌȓ$"6qFG	�Br03��E�&�ȓo��"	̕j�T�R�k�Z�~��8^@��0Oj}j�J��_kL��EPu��q�"	�c�fKl��'�p�A r�X[eA�!�I��) �Pr�b��L󄢍)2�$��ȓ���"r��3" ����-D����ȓh� ,�R�)����)sl
`��&[�`ka���V�۳ ڣg�)��(jx�2��Ό���3�Q4:�4݅�t�TH��^� ���t��R0�ȓp4���U"��&tjM��㓅d�����(4��&�Ք���sC��d��ȓ|��q%cwj�X{�L=� ��>*$=1�a�=JlУ
�a$�ȓ!���@��nx���#GȧbДl�ȓ;#lxɖ�xf��s��AV��d��%��4�V�$�,�{'hL/*��Y��`S<A��-�PT�[�C�^ܔ��g�C0� +d����I�>���#�tE[��G4]~� u眻&�Ї�B�8�iӥ����܋"%�;D$dY�ȓ��M��mϣ/7�K��O;A
�̄ȓd{T��d��U{��3�0!��r�lY�b������O�Y{��v��La#"���̠�EN m�ȓ�"��d�O��� �W�J�L|����h1U�D1n�t����(]�Y�ȓ"�$$9W��-X�|�îP�xP����ʰ, ��_�M'���#�Yl����ȓme����_�[`����N�{�Ȅ�4R��3 c /gĈܪD!�<+����ȓ\�N5����T�x|���ָ-�t�ȓ�\e9wF;�,�%�Y2wi���aD�HB�� ,����N,K�q��S`����BӚh��2N#2����-=.���/�	U��u��"ڨp�ȓd�^|���/X��,�&D`j���L�l����g��� ��'B��؅�=!�%�v��.��A8rn$O���ȓ!�X@[ �U�z��j�'�Bw&����\ �u�iOdR�+�"�:��ȓ3���j0yFb4��?�&|��v�"*���@]�u�V��{�P�ȓ|ގ��ʘ�F�1�h���<�ȓU�1���6B�Q�@j��D��S�? P��LB]TPh��c1@E�LAv"O�%�G螲@�0�RU�>���"O�(�d��U=q��ī)�5:�"O���B ĬxS���#4���"OM���"ϊC��G����"Ox�rGB&�*et ۿL�4��"O���Ć�!ɲuR��3��<#6"O:ظ�	��5B]�D�6�p�PE"O�+ʎ���2�b�j��k�'K���*�tt�9�cу0]��'�D���%�.-0�MJ�gG�e���'?:��g�<n�hqEE�w7���'l�����o�8����߅!���'o�X@��Y�'~�HA����]��'�İ#�јH>�U*�f[��3�'d�E�gA:r�0 y��ݚs~�p�'�-��F:*<�$�1|�P(�	�'��y2$¿0�Y���H��*	�'�(�T>4����I
$i����',���hD�a�10�<Z�2��'���;��C��B�{�G&O��R�'D�AB%��~�E)�G<QF�(�'D�,��^�,��iA�FŇ2m>�
�'V���*�T���ye.N9~8�J�'�@�6�R 7�`���
zbN��'�j�A6/U���fвo@Zt2�'��MĮG.�^���I�Q%��؏�$�O��}���5=Ȇ<h#IMd+e��y�<qCK�8K��jUB8p�F�B�Is�<�b!˯�̐�UiF�L^���l�p�<y�Ғ&���;�/@ 3.�)JDl�<!A�>W�`ࣙV>��k�d�<Y!B7V�p�#��A��Z��$Ēy�<y�F}���T`\��4#�C|�<��^�(Y��PwX������u��E{�U�m�I�"F� �ѩ��ǝ�y���4!�D�HS	�����Ɨ�y"�Ա6�\ B�A� I�ɚb���y�%<ޞq�g�À-�Y�m�yb��-v����ĉ'B$ZE�ٕ�y���3(n��E N9'Ģ�1�k�5�y��./>bd{U��3�(5�$c�0<9��1�h;�'\N�#������{�IG���T�!np����cOB��G�<�ybMR�u�Uх�ߦ0����(�D"O`�bԄ�]����rd��L\�Z�"OZ �W��	��#��'uxt#�"O2\8P�0]������Z�0��h"Od�����J��χN.�St�П�D�4��-%Z���,��p��Cɧ��d�<1H>���h�je�H���	�c*�]CrA���y"̓<#�ȼ*SއRdDs6f%�y2@��|n��!g,�G� ܩ��	��y���B�|0��2F~�XYw	̎�y"�D�p0Dc��ln��B&!���y���~2���v���k�v�u���0=a��υ@n�tLQ�c��i���<��'�ўb>%���Y f{.��f����&0��h9D�x��H#-G\�)�U:fx	�1D���c�	T�z�e�}�ܥ;� ;D���#�T���!��x���y��F{ʟb�O��3jBY����0��u��0��"Oa�,�H���@@�P���"O�(�MȮv�H[e� �^�p<;�"O� 4d�⛳	��97�Q�4J�"Oh�ɷ�ړV�
Ź���} ���a"OF}ȁ��]b���Í��[6��"OL�To�,
�MyQ慭.j�+�"O�uɺN�z��cd��zV\��Q"O��B!���V4)�Yh1NȒd"O��3BD�w�^��t�<$ ���WO2����&݌ܢ�+Ǧ �v\"dNP:9�!�dE�x�0�гA�p�k��\�!��*Dժ��#�8!�V����&�!��~�,�@�B�8@�E8
�,F��lI3���bf+�gİ�X���y2�+[P�)�ge]hN��Bc���0?�*O�<�.��˾U��L��`y`��&O\�d:.(��fǣ=��
��V�:��B��

��;5�Љ�eK/�PؚC�IT��貑��5-Z�@���;z�B�	4e��M�go�1p2j)犀(B�B䉜d�����
/)�B8�NLm�B������l�.��2�@�~�1�������l��!d0��Z�Yq�e�ȓ>�8��I�#)QT0,L9��	�'��P"3�W6E��ӆ��"z�v=��'���b�j��[���'I�t��u��'9@9
a���V�A�EǌH�J�'کi��tv�`�mO3{�H4(�'L�x���_"%�����(�h;ӓ�?)L>!�J�Zʐ��+C8�RQ T!�_�<Aa,ܸ��C�	ޱ5���(�l�u�<�E��"�ZA)u���D�Y�n�p�<i�(ӷZ��1��-k�4��&�k�<�1腾)��3�R	� �`]@�<9Q�/ְ��i�i����y�<-Bh$x�BX"�	#l^SP�B�ɣ8Ւ��R�ƈK�����Z�zR�B䉔ap���oP�z�l���;m��"<	ϓ(lDP�"��DL��%��{_(݅ȓZ�| i��$s�mKc�������9�Z�#���}���d�#aQXń�	yy����bƁ'm$�:���G�rY����d�&P�����;\�;G�+]!򤔂�2��Ћٝ4 ;U&<N]!�DJW��}���KtL��O�'8?!�G'z>��h�=-�������Y�!��I\���'*	f�+��%H�!�Z%��X�*@U��Be�T|ra|b]���ɿ:�����f5���1I��B���������j�<-b���U�(R��^h<��'ћS"R���d��2X�S�V�<Y�"
�~eb$�J+r\����	]Z�<��{e���q���c�L���JX�<9�ׂ]<J�����_���WK�P�<�4)�'���ދ���1�I�<��M�I>�˱b�c�����F�B�<	�HF3x ��L� ��R�*�|�'iў�pn�)�K�,@FIP4���P��5��۰g�:~h���6q�ȓG�xQA�(�)4zF5h�dD'k�4Ԇ�t^J�'�:x��������B���% ��)���-B[`
c�q~��ȓg/�\@���~�Q�+�<��D�ȓ7s^k'�Au$ȑ�y'@�ȓk��r0lr�`hIv�U>��L�'�ў"|"G�&��@V	aHХ���W�<� ����FLp`�s%�
���U"O��ūL�8!*���oۆXK�"O�c	�b�}��"�/\��!�"Ot���ӗ}������.k�0���' �O�`��=�P��`���U�4�Şu��E�aE��и#KΝm�H��
����A�0�U�7ǉ�`�R���bQ\h��b�2W:h*�`V2v̕�ȓ=���)�iF5Yf�r��<Ѕȓ6��t���I%4�f
�Ʉ�=��хȓc�|
���S!f�(֮�X�B%��IX�'���׏9q���Y#�AO����'� �;�A3c'�<�Bύ�I�@�(�'�f��P�J5z�H�&G�Glp��
�'^�bA�Ǯ@�:�1��.\��
�'u2D���ߪWW�8`E�Y^�M�	�'yu�
�|��� ��"Z3DL��'�pI"Ԣ�)�fI#�e+g��Ͱ	�'� �I��4�!�,��Y���'����A_D��ʃXK�`a�'��93�+S�?Ո��#	�)9�Ԅ8�Oأ=E�t����f�3����;�8���-��y2�{�lA#�]-DM^ru+R�ybk?@�x�p�OL:(����Bҝ�y�j�
�L��Ȋ4�P�[�� �yb�R�B�Ɋ���"L,`��9�yr�E�7^@���/ ���C;�y"��F�M���Ę� q
�B�/z�IF�)��<�և��<���#`�,8�*x���T�<ɖ`�3�b���Aѩ/�����$Y�<AcC�iܔ�t,�(P����V�W�<a�On�PċF�!>�J��$�@���x")%1�����:`쐒E���yB�݇c���󲢊�-�5z�`���yR�H>_'^��&E/R`�����&�y��Q�\��Y(BR-y�01jCfK6�y��]+SK��[�蕼d]H�I0�Կ�yBg\�a@�%���O�`v1��e�[1ў"~�)|�9IT�0�2�z��F;e���ȓ`Q=6��D&����8!�hH��? Iz�H[:E�-(���;"w�ńȓ~�$`1�R�o�J u��9L�"�ȓ.$��r�;F�
(�th3h\ą�
o��R׬��`,qӕ0+8}��YpEq1�_"J�*�� A7;4�Da��4���<�	-u���	B(5��#"-�fB�	x���iu:Q��\jR��4E��B�	5�|֍�V��t�V"V6X�����>ړ_���*�2
a�(��J*=�E��K$���v�K1<Ɍ�[� �"�p��ȓ�R "���^|x��ҡV�F��ȓ%���8���!l,҈C��aD)�<q���dX.4�ĥ�G��Kr�4!�k@�Q�!�$�bAXa���^�m|�P�̔(�!�_�v,TX�)I�14�= ��Y(5���G{ʟ�cvM�/f���瀚�+=t�2�"Op@�0��6.�HD�
��
T�S"O�Y:sKF9N� q�/߶J:�m��"O���ĥ�
"F )�-J�Q{��j�"OLP1c6;��xCÚ:��H�"O���c�D���bR" ~�R���"O�h�dn^n��t�B �Ec�h���U�O�v�qTK�?&�E����5 ���x�'/�ic	O0#�h!xǧ��Y�py��� B�h`�Z<�Υ�tNV�q�z�b�"O2�a��Q$)�`9d�ڱ(��(�"O�M�S�V�Z#�`�y�:�4"Oд��]=e)*����R�H�`1�"O�0��N�8Y��t����+��Yq"O���	�<�ƙ��A�>+bFp9�"O��s!��s����!`��s��P"O^p"��L-,1biZ�/�2"��d�"O����`���@�7���"O�؊ &�)dQ�����[bd��!"O��h��}�|�ä�*B��SF"Oj���(r ��#c�1J���#�"O�Xj�O�	��:�l�4�8Ò"Ob8۱q�
ћ�j�c�H4B�"Oȝ��(��������<z�Hz�"OD��£�/!-��"�)TP�MA�"O&�Rta[�2eR]pB�+ZU�v"O�q���0Z��!$@'Es���D"Ol���ǣ\��m�p��i6�'"ODra�G�s�xݳ�e�rА"O
mɀ�D�Q2��w�ӂ��jt"O��a�Ž��h��O�"�ڴ�"O:ԀG 8 )P�;vO߭U�ʬS"OZU��]:p�hY�� ڪ2�`���"O��7o����Uj�=�u�r"O2���ի[&��#jE�_�nXb�"O:�Q⇋#:�%KFBW�i�D�{v"O
q0��,ު3b
�=��$3T"O�;U��_da����;8�U�"OR�)A���g*�0
ǃ<d6d��"OƠ ��
[P���d���C,�Cs"O��p�ģ����hE�cT8�"O^���ƖI��,z@'��l�h(�Q�'~�I m����@�jl�R�dސAfC䉞|��9RԫK�0x���Q�F�dC�	?1)%$�Y$�1�9/ �B�����Ҕ0�YX`�٪+N�l�C&D�$�g�fɾ��%4Qv�� �?D�$Ӓ$��Y*P��h��}
v�9D���&�8'�T:�i��=�8�Z�f8�OV�O��*��_61���j�Eq���a"O��%�Z
+��۶^�g�C"O
�ǍD"z�;�l� X>l�"ON\���
�0�:��A�ӗb���'"O�TR�m���U8�*K�$g����"O����EN,D�`��e�_��ʲ"O�!�e#m�e"EA������'�剷3����йk���A��0(�C�ɬcQ�m�D��h��!��m)�B��3�@��@YB�h[���jj�B䉲l<*9�U&g�j�z�I�j�TB�I�*\�4��W.@��:Y�Գ�l D��	�9`�1��.Q-�:aP�'4D�<!Ą
�H��ч�ϩ8������=?Q���%7��" �U
:��\���X!Y�B�ɀx���Bp%Q9b���k�V�|$B�I" ��J@�W�Z�]h��׿p�@C�ɳM�x�	"���DT�%'W�$��C��:e=��5�
�v�ç��5��C�	�8��i��׾<M��鎅ۼC��|K:D#�������*�>��C�66r�6	��K$ً'�I
S�C�I��Ό���7i��,�CD	|�B䉣[�H�fn��������'�B�)� �4��ȟ2����5r��2"O�lɅ�Jf���$냇N�2x	�"O��R�P�A*���"�Z>�
m�b"O��q0��e�D�����IB�"O3	Srhzt�0FX���qK>�!��l�Ӆ��3��ȑ��.]�!��G24�`{�Ȓ�>����'@,�!�DU�!�����6�&��1A��r�!�䏻rUV8Y塄-���	4�_Y|!��\�G���*�	i���I� h!���}ұ�R�ņ_��I�E�q_!����0Y�@��6�(	e�Z"f�!�D��]F��M����q���� h�!�d�'*��FȉU �hkP�C�!��O(J���ʒQ�ZyA#Ǝ�!��̔Uيi�F� N��R��u�!�d �JRH� ��	E8R1�U(^�y�!�dYl�����7�ęʄ猦u�!�Ć�-�]��b��]�X�w��l�!��(:
1�e��=fLE#��t!�D�m�0ǁT�昢v ԝ'�!�䚣"T���ĵ��)��9g>!�$�y������
�F�jХC��!��1j$� [�kT�[��@�g�!�D����G	��	�C-�w�!��]�E pb"쒔)PV ��NQ�+N!�h&���E�F+@<�I�_E!�d�>ANn!����h"�wd�1!�䘨q�Jp�@��B� �P�bĈ]�!���<r�4	�Nށi�F�K���U�!�dùk���qa,4s�����	i!�$�4,bz�҆��C{�I�@���Yk!�,hYR�(� ]��jpf��2�O��R7 �3iP�(i��ߩ�B%X�"O��+�Iڷ;�Fu��c�	0pQ�"O6$q�ΎGԆ<q�AG�/�|!�U"OΜ�G�H#|�:)�ĠT��F��"O\$p���oДK#e��E�����"Od-��fD`���w�I*M���xd"O��� ƚ)5���t@W�Ԝ�b"Ol�ˡjG�]w>���O;=�4�I�"Ot�1⃫lz����̷e���	�"Ov�k���s�(	�7�ߤ�x�d"Of�!%��<M�8��#B�f@����"O���Ec�dQ��a?�U�"O8�8��l�d���K�9'���p"O�e��M<G�2��nW�@� �"O��bN�ecнۂ�V�\��D"OB�!�gP�br�9ԬK�B��H:"OT�S�Xx�X�Дl�W��W��yR�S��]	�ϨF�R���K\��y"�/�h5��E��>��}�G��yo�/KkxIC��_
$�jm�q�*�y҉ȹ�Q�EU>�	�P�M��y�.Ԉl_2B��~Y�u��}�<I �5���D&߽�68�i�H�<���>��%�#(z��"�#��y��Y,)�Z�����s�~�2�O�"�yaǛc||@�3/�s�XY)�y��N&�&5pR���r��&Y�y�d����5l�j+�Y���<�yr��m�Q"�aH�]��Q�TdD8�yR��+���hc�E�����ǽ�y����9 ��KQl��f!��J ���y
� �Q���E�m��<z���9����"Oz�
�>��`Pƃ|���c"O�0ɠ�H�	B,����
'y\��`�"O�e�@!�(������r� W"O`��qg�,u�Ī$!�-����c"O�8�C΄!4VuJ`]�i����3"O��I�!��2��0dI0(��"O����J� @�AB�Dg��T"O�J�A\/g42�a'oV�9���C"O�8�挀)N$N9�ҀD�*ڎ��2"OX�B�@��.�����0�q"O~�!�L-RH���r�P5�"O�us�F�5o-h4�7�2 �P��"Oj(��ϲ1��l����-!���x�"O��S�׋]O�iQS<蚑�"O,j��?ef9`D����D:�"OD��k[Z��5�� ^�v�$h��"O�Ր�c��{X��`�o�$A�p�sW"O ,�d�Ba�jt
c�pg�%�"O��g�
�c�	�~T�Y0"OR(A3��*���s��rG�xA7"O��4Kܯm�L-���Ȝ|�DmYq"O�����J6�F�H��D�ft��"O��a��A3�<�f��l����"O`܉Fmѕzv*�3���'	�Zi�"O\��!f�/X�'���4� �YT"O@�܃M�6z=J�X׌��Ba�l�<���p�.�:"�A�̰��<�y� �T�D�*�G,f���bk�4�yb����i��BNY�:upċ�(�y2�� C�8Ru&H�n��4��y��ۂ;���I�	�B%+�,���y��v�&�I�F040�JU/�yΒ|��R��sAr�$��y� B+󴁰�@R�-&}��o�y��F0��(�sC�^Fx�7�2�yr���UܠI����_��E $�@1�yBF̦/i����8Q�V�p�J�yRᙶc�0S�G�n��[�#��yRK7F�4�&�4�ؒ#X��y�i]�"ؐ�@[�*e��F��y��3��9��R�}��0rG�Ѱ�y�n_L���(v5�l�e����yBÖ5.6-zB �X�01��ȫ�y�.	#
�R�a�G��RE�,o���yRK���n�#$�`;J�I���y"�|�T�b>�v=�����N-lr�E�Fo�)�,�ȓ.\��"rK�!��Y#��bn��5e����鍶kڍI*^
�a��Iqz�B�E�$��%��M� \هȓhA&��B*I���@���\5&5t܇�h��0�c�5xzmK0�0El����a_\�BWf��DV�Z�d��͔��Q�&	S�	���B4�ҩ7� �ȓWްH�F�db�0�CX�-�ZЄȓ",lI8��Zq��y�ē�K����yC�Q����
~��t �F5^��ȓ
K\����G�y*�`h@�ДZDA�ȓ,������=ҊU��K�b����!�r���@@�)��OX�G�
��ȓBN�4�F���]��
r�|`��w�^�I ���*Т�aS�T�ȓ+�l�����@4:I�cnLs(�ȓl-;�DS�jV TG��3D���S�? �1"�Բb�Na�����&C��1"Oʤ���g�J����ɓ	^���"Ob�kH+9o.5��N�U�Az""O@�uϏ��0���氫c"O��Ȃ��>"�4��v�	Z֔�S"O�8 ��Hh�R�iÉ�h/@!b"O�\���X�j�&U# #g�5B#"O��p��0h]�2K]�nX��"O��G1b�)ѷ�6S�đ "O ����k2�ŉiݜWv,�1�"OLl[�JAc�<�Q���Q[tIy�"O��GaR�A�z ��%_�#�$;%"O�@��-w��BӤǞ��E�5"O�3��Ӏ>�T"��zNM�"O����,@<��k������'=ўx��D��_"����nS0��� �f D�d��C:B�h�r�/������+D����:<x����v� Ui+D�LhE!�#a	cF���P8i��)D�QK�5'`���K���&г�j:D�(��@�#!
d�0��qTm4D�PF+�!c��@f�Z"	F��#3?����h�  C4�7{��ua	�%�b��E{���
_������_X�����ɂ��y���3S�:�`椊�z��hC��_ �y�̟2d�I��\,!W:�ᕭ��y��� E��T�֎$�5*�y�A"O�t�Ƭ�;9��q���1�yb �o
�xɑ���>��B�*��OZ�=�O�xd�Fʜ
4����i>4�y��'�����'��t�T���ےs�¸��'Π�C��к+����3-׽qu��'I�`q��<f�\U;��T�k��Ԩ�'���=L��N	a�*}z�'%��s��$�r��#M��C9<�
�'0���`���{��t��/J����O�=���KG,���I�16|tQ��>��O��3?��)�:�����,h�����TH�<�F������O56��%h�G�B�I)@���R����NsH]8�Փt��C�I7
]�	(b�Ƀ�2�R2�..w�C�I+3C|	��̈��ʈ"�g�A?�B�I1�¡XWC� K���P�'KtC�=w:p��$#�td��+�M:%b�G{��9O�) ��&��&dF�d�,s�"Ox�KQS��:��V� =?�0l""OX�)�U6T��qʒ�"Ip�mxp"Oʰ�C� ����[�V�t�V�I "OLX�@b�;�V��cF�2��l�F"O�z�BQ 
��3�S�Md"܁"Ob���Xc��@S7�ǀuV 8�b���DQ�8��p��t(p�IF�R�H
�b��C䉡2j$Qe
J �ѳ��'n,vC䉫P�$䙤����@��f��� t�C䉾a�������=\�(i�D�\s��C�	<�(u�7I,r[�v�X�*=C䉮��D��C*y��������K��">��Iǲ=�����đ�uT9$��W���sx�hR _�A0�!���	*�ĭ��2D��`C��>x��9��kf�H]���0D�ԩ�c�J/V}���ݸ|rFE{6/D�\34��E�t��Q���N�$�1c D�D�Eb*=6��h�%E*w�\���f1��hO�ӭT����eY��D���>��G�)� f��3Y	���2a ��lp<�(�"O\İ�mD�5��9qA�I/�|�Qv�d$|O�P�T��.���� �v���S"O�$ʶ��(aR.Ѣ�m
*~H �:4"O�9�َU�jiD���=5|��"O]��� �()׮�$(�E���	{���郣�T��E¢)��Ur@�I?�!���l�E���-�6����|��d,�S�O
�V�Y����y����N����'>\Hx���$Z\�)%�Z�IW|�'�
�)���n_�	���K;,����$ ��Se�f��9�R�C7�\��*�c��v2`y��/Ɠ�t�Fx��)�$�X��8x��n ��y"�Ed�<�cU�?��� ��kY��Ѓ�v�`��_��Ev0- EU%&�𑳦%L��ȓ.}VH	%J_�R0\�­Y\٘��ȓe�t��A�W�
-�V��?H�l���?!A��7QM���G̟�3�f)��v�<PfK3q��������E"�x�<��U-L��q`!|�6��F�v�<�Q���!���k�%�9nF,�"cdW[̓��+��vAVP��	]��0kE)%)�v��ȓd������(tQ{��H;r���2�p��d��?:�מQn���I���I�Qy�,���Z�D���ƪ�FΰB�I+5��-��+K�s�4��g�R�u�x"<Y
ϓR<�W烐T{l�t$��
�xل�v��YJ�C�>&�ȰB�dQ�����'(�'��?Q@�H"-� Xy0�^NE���%D��e듟yR��p3Ď�X(���r�&D�@�"I	�`8��n��j:,\;Si#D����h��-�-ys�q���%H"D����	�b�`�FK[�a���Q6`<O��=)4cя�T\�q��F�p C���p�<�!��Z�4A≉�=��
U�3�hO?�I��|8S����
hSa�`�C�	�|���r��޷:��mu���c�C�ɲ?<0��假
[�ԍ+��+O�XC�I�o�,���LQ�x��E,^[�&C�I�{��Eb�oՀJ�Z��ܠ]����(��Vd&����M�v����!�H�bB�ɸx����@�D4nNѻdεV1zC�QU�B�"C�ny|�3ɋLYDC�I�.�P�:��3
���d�T�C�#}� ����_,������(L�B䉅c�8u0�ʄ�iBn�X�獒(��B�ɀy5�z��03�tg"r/�B�	�FC
��g`ɠ5f�V��ʎb���	Oy"S��&���DGH�5[�-���`ǘdq׊'?I�oe�EVh<2�,]1S�D�Q,P؄ȓ�x��J�#\�th��"
^�h5��wT�t��Q�*`QXr ��
I��=T08 D��6� H�S U
-��ć�Z�&��i�vV����+I�x ���ȓf*�X�U)ԇ;h8��D!�	b\�A���I�O��	�t�*5��h�C�=
���_⼬�w�:�L�e6;c�y�ȓfEu�C튓HN �J�̖6y�u�ȓa�*L����&7��8�W%U/�%�ȓl9�����(��1��P]���ȓX���i��3 �������2����Wi(L���66��E�@BH�^vp�ȓ=֠嘶�H#5`�6J��H��S�? P0��ʖd��,���L�q���ȗ"O�@����pFM�C�T;���z'"O ��OI����W*
eQ[١"O�e"fB:wXt(ɖɛ-A?d��"OT��� �=5&(yQ#�� +^ ��"OLh���6�p��D\�m� �#q"O^�׈��]Ur|�1���h��"O�L�q�C�,nL�8b�n%H�S��O�<�p��H�	�"�
��'O�<t꟣0d2��Ά�<h�d3D�ı�Ł$D4��D�ΩN� �0D�@K������"�May�hI3H1D�Kf�][Nj|+3�G<E�^(Ʈ0D�Pd��>'�4�$� ��4X��:D�D���"x��-�&�7:=��r�;D��׀���7eZ0�T�qצ8D�H�6KG`:1�N�<���;D�X����@6��(��V #^�t(XM�����$� H� �@C)�����g z�!��{&���N�aP4G\+8�X�D3�)�@�	�Y�.��j	�6f%
#�
�s��B�	����ӆ� ǼѢR�ۣ!�B�	�Mp���wG�%u���!B���B䉜zǪ��0/��=D](�-ϲ�yRcH{ڬ<����R��y�5
�y��F4O�@l���ӥV.8u@��y�H��'�: a��"/pDI��?�y��)�'z�D��Dr:H)�T�Sj�Ȅȓ~h�` 瑄:�� ��GՑI��=��4����4[%"�(�A�3c� �ȓ4�ā%��)���k�FH�I�n��ȓk��RqH�b������+Wg���
����R�ZCf����FI<B	�ه�`��!��e�j�Ag��!,QP-�'GR��(�S�r	�({�U�/���``F8Bi�C�I$)5(8z��_6 ��zĪH�~�2C�		8w6]���N���"���%�PB�	2t��%[����U��Ti���7YL�C䉁YU�4���9v�,��P3qB�	:2̨�oȒO����e��}]�C䉣b�>E��Ɏ9�v��Wl�i1B�I�_��-�!X4 4�J�咂[��C�I9]2��*T�
�Li�� ��W��C�	>�Ĩ�d�Q��"}��KݻP��C�>4�t��_�)���q%n�-�!���(I�$P�#�0a�u��Դ7|!�E��%��c�,mv`��� qO!�d��av<��KF�-�Jܹu@V�{�!�3�>*2��2zB]�qfX�Dt!�d�� �i��D"R� ���#rm!�D�2^�B����D=�z�E�>WR!�d_�Co�)���8D�A�ׯ�!��+Y��Q��1k>)�e�ޞo�!�dW�+���A�#!�rQ�b%�q�!���tY��G1,��D�'o!��F�JDa��ٿ`�b�ZvC�a!�$��z���Ч��x����ߤ^!�Ă�/�V�����(զ;w�&!!�B?eĞ�X2蜬!�Б�g�-p!�AT1*��k���y��4�!��̦�
�á�\!���Ñ
+�!�d�B�ʥj/Bx�E�f;L��"O�	�ϒ\�H8%e�%#��U�3"O��:$�ԴF����Oϛ^@��"O� �J=�j`b3���fC��"O���-�?O9�0$j4w�
���"O�D��Ď� ����a�=I��5D����@�)�*����O�/lf��W�1D���S����kի��8��=�v*+D���L��W�f�D�j��@,(D�xb@n�Y�L��L8u㾠:2�'D�(�	.3S$�I��?pܪ�K$D�t���H�X� ����6C�LlX�"D� [U�ݥOH��s��]�k�\iz�h>D�dY�2�ڴ��X�V'�P�E:D� BqFگ\<�p��%��T�1(9D�Ě��W7�,l؃�����[��6D�Q1-";�*�zUo�nފ�*�l5D����E��p��e^��V�bpJ!D�|���<jU\�;��40�2��6�2D�X���},*5�S� _�.�6 &D������D"v(�K؀Ln��v�.D���#@�A	�����'��X-D�P��(%m�� ��:5����*D�T���S��)���X�t��/.D�Ã�7jZH���D�x0n�0��-D��2���*>����7-Ƕ\C`i#s�0D�(�Hڇ##N䫆GoC~	Z��,D���E���q�1s�U9d6�!,D���C���GS<=�c�S#r8 �i(D��k��'IZa���0m�,��4�%D����l��D� -���;8�����!D��A`�TM� ��PN��y|�Qѓ�?D�X@3� "bP�C����Az��>D�P���2��S4FI'M6l|�U�:D�̘n��]�2�s�HF�\����T�8D��8#�E?��9�*�	bik%6D��cO�/���3� ��>)a�2D��Z��\`\�+���t��g/D�X�V-F��I�VM��4x��B�.D���̌�]*ʭ���0�L<��&+D��c�
[D9�}K�&�-e��I�T�4D��2@����d�ȆAȦՒ��$D��p�C�J@��p��۔�Nu�w�$D�|Q�B�T���卛���u7D��
�/
%4���ɇ��.ؠ SJ8D�t���о@o��bA�L�/`�jw�5D�,y����u�&D	,E��Cs�5D��*���E2f�B`*��t�hD2��.D��P��_%7��Q'���ql�hP.9D�$���%=ي��2��0��*��7D�$�AN�o@֐:R#_C�"�p�%3D���c�3-\��g�\}U�r�<D�DGJ�Onz�#f#,Ru��s�C9D� ҬC*Lt���BK�1��(q�)D� �(M�N��-��#r�\9��;D��@��۵,��� S�Ll��u���:D�1v�ܳg�R9*"
� w�Eh��5D��2휴b8vU��d D�����'D�|����?'����@ 3��c�!D�LPe�(r�8���<�by��l9D���
ǎu�h�: ���;� [�-D�$hQ��&E:�� #?��$�,D�#�d�2��H�l֢�bU.,D�(򭜅
d�j�R\�l@S�(D��A*�@�Ψ*B��:a�v)k��2D�x����8F��!ΔB�L=�$�<D�T���P�;/ y����f@�5(.D�� � )%۰i�&`2����p�s"O�8y�-K)z�aJ��F��a8�"O"�A���� �� ��%��`��"O:k3����b(�5!�H�Z"O��Q�l�^b�Zf@�l� �� "O���ㇾg���8��܈YU�ɢ�"O��2�k��1lJ�S�H��[$	J"O֥��菛^X�sw.��1L �C"O
��3B�1 
��ML6�``�"Ol�sW�<�b<@&lM/#���ڦ"O�k�e�^"a8�$�p���u"OL��V�L$��q��!��Z�R�(�"O�3V���b��T�AX�Z�:�:R"O�����}4b݊��!c�T<ر"O�=hA%�!���"AF���P
P"OrXa�M� Y$��$�j�@� �"O��'�'R��0r��6�
]��"O�I���R�e&X	zG��Xw�Ps7"O4�A6�b9,	B�`��f�qXE"O�m��lV?L&V���o��q��"O|,�a`�$n���ᶀ�X����"O�ѻ��72�PD�e�â?H�z"OF1���${�:�PmTP 1B�"OB��w�М	֬ل8E�W"O����΋X�V�zG�3�%��"O�h��U�4�(���
;�]R�"O���7J���)�04��1	t팑^)!�:�N�2���J�B	��	��o�!�$�m������4PWHI�sI�+By!�[�30�9	�L�<vK�xzU�!��B�	?�X0"�˶7 ]xs�W� 
�C�I4E��l�s��*GF1���uI�"O����"�'�[W�̆+>��Y"Ot9Z�ԗ /�<!���T�2`p�"Ovɘ����:�D���	�7]X�qD"O���u
�_n�i2�UP���"O*�0§B?B�rH�C� (��0�"O��X� E�7�P� @�
��G"O��2����ћ@o]��1��"OhT�TG�N̤x��ը"wp�"S"O$�(EL1q̐�#��(�Nx�"O`I%��GDP�!��D7z*�z@"O�IѶk�E�n�3�&�	x�w"Op-Q�۪%�J�q�K�rO 5�"O� ``���'��p��+
���l�"OtAgj�7��E��&����"O�$�S�B�t:DJ�o�t��"O��2���1-U�)&+� K[��X�"O�Q��J	a0���@�/���C"O�R㮋+2�d�ǭQ�9�ni��"OH�Z�.�2^�t93"��X@"OL�C�P�IH�0��Z��B:�"O����MAsH�@uaF� ��]��"O
9A���$	����Ӡ�o���2�"O��W�83K�DZ�ł?f0!�$"O��k�:\HL%�u�ֶn_�:Q"O:P� m�B��h�2d؏����"O�}���ց!C�p�
H"M� ��C"O(�꠫=3�񡠩t(�r3"OJ$�u�:Dl����x��|�6C��.v�C�&��� U�W"�
j��B�ɚt.����� �4��UCH�~�B�	'r�*� �RH�Zk�o��B�	�e%Ze��랶��1[L^9ΘB�)� ``XU�K�'�,���ぁ G(�2"O�����؀~\ܸ�e��S��yh�"O0����)x0��W�?ai���'"O̍
���+愠X�bƔP��J�"O�0����� ��ק����[�"O<Z��M�l�4Z�,@�q�����"O<0뗅�0a\d�[��� T��"Oe1c�l�:�E��4�0�"O�q�k�8�0�x k{r$�z�"O�Ԡ5�ĊBs�$����L3~,�B"O6�1S�+�b(ca��n}�]�"Or�p��KP�)�?okbpv"OΜ+r�ճp��eD�&H��|�3"Ov��咨5J�I�ȏ���g"O,��Ƴz�*���gD�o@:T"O�AA`�ѵ|��x��$&h̐��"Of�
 h�>k0s2�W>a�P�"O*	�%��[� [mثa�ԡYu"O�<�b'W�U t�b��,C�QIs"O��#I�6yՀ)�	H� u�v"O�0��,ۇ^�.%y��G�EW�0:g"O"��/�H��� &��0��"O�̺"J�Z�i�U���A�ӕ"O�(�'�էPu$��ЧK�)��� 6"O�u��60��A���V���{�"O�-{+E�|KX�j�(t�ZU"O����δ��I���=X��0"O������,y	PY*�.ԉR�%K�"O�����Y�J�0�s��Y4`�p�"OJ�觎U��lr`��
Qb"O�� C �/��Q�ETs���"O����NJ�R�>��&�Qe��p'"Ov�R��H ��-G�3ch!�G"O���%��%�蘂���J��e"O��r'��4m�*�ȏe (��"O8�!ț�n%ЀK��	x��5�b"O�������Va
%�h"Od(��-ZX��P���8��<�B"OV��j� 6��!Q	�s��q�"O(aTG7@aV H.�����Y�"O�5�pa�(>��Ѓ-�>V�6��"Or���ˋ�N���Q �W�"��Q1�"O�ҧGU_6Z���I��Mc�m�C"O�@2!J�&F�r��t���.y�az�"O> �$#IdP�Rl�d��;�"O^,h�C"_Z ��>���
�"O쨑�P�b��i 6=+�"OTБA�t�B��WC��8�$�D"Ob��"�f��9�ƈ�8�)g"OZ�� L�-󺽋���gp"U��"O��dY������@��!��"Oq�e��&��!�'NS���"O�d�s	�aԹ�֦_�J�Vpp�"O(I���=�����C���!�"O2 �#�N�i�=	�
N�|����'"O��
�#��@r�����p{�H"A"OT婥n�g�H����x�(�y�"O
��фU�*�T�����Wd�̓�"O�� 'ފh���)Lh����TT�<Y#,�l�x@Q1�X�B��S�<����_�0|��+U*/xZUm�w�<ѡ��J*訙e����DRP"�<ѲY $����BJ�tը8�a�[}�<9N�L�`���qchE�;�!�� �iI��O8�� ��K�_���s�iϡ�ă)D�\��!��9�'�X�1��zb���1�P���g�&]�c�	(�!�@nH�Yc( :��[Ì�)J�!��!n����ȑ|�~�kckÀ=�!��M2>�)sBCαtrp)����!�Ǳֈ�����a�A�=�!�Go�(���3	H6�Qr�,l�!���9|:¼���̬YF,�c%��{!��H"\�=�8O��� (��r\!�$��FTcRh�t�I�rԿ7B!�D�>,���J�s��L�񏞴@�!���K �p4͟	=j����Ճ/n�	x���@�
;\�H��cZ�%v���D,�OZ�'�fl;1jM&X�$���	.U_0$ïO"���I�q|�@��_.����'�Q��Exҙ~�҃����`�.Ât��ͩV^�<iV@��J���[5A̻L\AJtF\��M�O�4���%-��� ���Yٚ|��X�<Y�G[<�j���?��a��Y�E�Q�lE��'W�5;���nPj���Xn��]h�')�0B�\�z6��aGM�Hoj��'h���I"}:t��	�B�<RK��i	�'W���LۣPE����a��|���'���"P��#�@���u�]�(OD�=E���Њ3�T�S�C.�l1�
Ɗ�y"l�.vFT 7'�0q	�(�B`ي�yR�K�w�<1�T�@�ʖ�-�yR�ܢ~H��1���s_���"@��y��a�:lxr��p/F���P�y�\�=:H�#���nXtM�g�A��y"P�{4,I
d�Z�6v�	'e͎�yrL��P>����aHDa�HR��yr�:g��y���]���i�o��yr���kB�+tD�>J섣B���>)B�<A�� n�*[�Ù^��8��As�<��Z�$4��t��az�AMZm�<��E��5���U$>���i2��j�<��B9��£(�Dq�g͗�<����Ec0�+vZ����wB�^B�(L颦�6hӊ�����;�rb����;x�l�cA�.��-��{�nB�8_Ĕ��}��qe�4ɔC�I�Yi�9�fņ&�č	�ו	�xC�I�&z��n��p�� �[nVXC��67Ƅ�x#��"bg��03Jؠ} C�	.5*I�E9E܌c4+X�!�B����A��b��1/�)c!àF�B�	�� !�$ő�Y��A&a�;tB�	�c����a�ئ�8�6��,,PB��؎�G�\�p:r��p`Di�B�I-|�B���!��}�����#/J�C�I<�潰��Tc���a��yC�I�H�HI���ǡW8��è  ֺC�	���I @W��p��6`��m�v7�$�S��M���-v���U�Ήm��l�,�o�<�7�ɐ[m�!��N؈I��`�Êi�<�3/@�R���`ցH]&�c�n8��&�����7�	��h&B����*D�32�2����M(��cr�<�R���)J gPސ"�ٴ�L�K[M�!��]a���pN�"-��H7".!���&ز�{��܏F�XQ0�O=$*!�dB�\�Đ[�ȓ���h���T�D!�� ��&�[�D�8RG�'(]j��q"O&@��K0r�&���1d�RaJ�"O�U���~��,����CҖ9y�"O�9��.ЩKEv%j�A�n��"O��#���&0��"7aI�Fe�]`"O�Y�&�,��I9>N���"O��ŉ́F��eΙ 2/D�0S"O�@׭k�j��-�-v�x�S�"OB�r�̶r�vg#�~�{�"O �aR�$S����B_Ryړ"O�}�Ĕ7�*�9��aABI��"ON���U4
����g�C�l'���"O<��1D��Вt��/8�\�"O.0�,������uLe�����"O��`��� ?(�Q��y��
d!��]�|�r!�6��J=L5�O4�!���5rB��7HPt�=�!�u�!���k���j�c37ǘT��-Fw7!�ñS��i��I�+LվQȇǗ�"7!�d�5Rp�p�7e�pK1�-+�!�/U6��e��GP|�'�B(!��
�n��i�y9l%��刡P'!�ăhS$���	��G6�hc�$K!�dW=��ؚq�/::}���-�!�$gH�ՙ���=dq T!R�f!��%M.��T!��w	�H�@��ag!�d�\p����KT�	���u���}!�+]�|{"	HV�AH��Śp`!��Ğj����W��&�!�/���!���QK�9Eo��u"8BƯB�?�!�dݨ-��u��j@�\ч	�!��,|��P0sƁ
1���8s&�H!!�Ɛw1�1�wEĴ`��%��J!�ĔG����JUn(�щ1�F�!�D�~tR�rS�^g�����&�!��Y碙��X�[��X�ǯ��!�dJLTz���G�X� �RX�!�B#1"���∀�Ջ\�,�!򄆩�	� B
~� �V�!���0�\D(p'8<�-��C�"O&8�F7�l|'N�#J����"O�p�С]��2�`�-�Qc\�"OP�0-�	��1uk�~X���"O0!�T"��/	��)p	�	V>�1 "O�QA��H�����_]��I��"OT��L"w��P�fP�����"O����9$�(R�HBȽR1"OZ�$�6w.��fUC�X��"O��1�@S /BQ��j΁C�ʑ�b"OLh�e���ưi����C�$I��"O��� I��
}�(\"m`u�v"OT�)Â׳r����8MZ���"O��9���L��<Y�!L� ־�"&"O�&S�!"5;��ϣ�̠��"O��z��S�hk��B�/�9u�C�"OD�Id�@/�V�PF��rl�J6"O.�@a������ӏD &�Sg"O>|�r���xZ�å��wu(勴"O~��b�(w*4��#��Kq�p�"OH���Ğ8��������6')D����OA ,��]Gn��_��R6�+D������D��ػ�m�2Al:!'/D�H8E/I�w�,P` `@Em�M��L8D��#n�S��}1��+�Ι��2D�� �����r״�jU'� I�䅳�"O�� `���k�rd��&A3o��"O�r��ND#�#Є@�{zx�(F"O��X$T8j�@�#A�1%��,A6"O���j�<(�ɺ&`!1w^�)&"O����
��cELfD��"O�-��h���e��L&v���w"O�\�3	Z4t��0#	[�\$9�"O����C�@�І��r��
3"Of���ظ:AIp��0!�X�*"Ov� .޻z�V�I��] ��y��"O�W�?�n�s��a2
��aMs�<�(X�9���QQ�Λ>����&HH�<y��|k�P�r�ٽ<�F�mC�<9�.�z�s��9 >4�&f }�<�S��#�uu!T�Pˤl�$�Iq�<�e�.@ZDQ���[�J�ty�C�F�<�F�y���V)N�I�H*0��D�<��ˎW�x,��t�!w�DC�<	�J^:y�����n��>T:᫇��@�<ag�*j�LE�և¼|�\�{�ŘQ�< �SU��pj��7��r�E�xy�'�2�kMP`0Q�f-�9cƅr�'DB)Hu-ҐW�~S�F83��ٙ���?O�C����W���@eJı`?��{�"OL�!�o��`�,m�cT�oӔB�I�t�`���e sa�Y"@\�B�0hj��e�
=�{1(���B�	KX��)�QOYB6�~Q�B�	5�*�;c�)� ���I�P�|B�	
50��R!	��F��" Ե~�DB�ɓjm4�ʱ��OVƬ
�f�$J�RC�	8Ђa�#,��nƮ`�a�M.\zN7�V0��?�C�U�v�(��֑VB��h2eSh����<�'��+K�My'�5�ڽPs@�d�<����5�X����|��d�ck�b�H���ǫ��
��2w�Jtj.,O��<��A�0PeN�6�ԿP��HҦ�V�'�x�m�!#`P��M���`H�E���yb�կ!ȶdJaJǩ�	R%J��y�E:��d*�b[<�4��/���?�'�n���Lȡ9�&e�W�A�r���'��X	IH�$��^�?R�d�A�>D��y�m;t���Rc��=�� ��;D�tJ�B�y�4 k��.-}�)2�:D�L�be߯bs*��0Y!!���w�:D��p1���PuF�[$j��Y慪�,D��	�jY�J��t�%C�8F<��qg(<D�4 ��A4d�,S�	J-sH"!a,D�tS��O�0��`�⁀�+�<���S�?��%s m� w�EA�kV�$9bB�	�u<���J,���թ�s��B�I�SB��Ū�p��|��DH;h�$C�ɦ=�A/�P�oM�`�׏1�O�O������6)h�x8Be�;";4�Q��'���,����h�J�P£�f�X�� -ʓ�hO�S�O�FlJ�n� g�A����@;|B�	bN�J�BU>h��˟�S�@B�	`B�I�^Ў���ޢO�(B�i�5ҐDE/ ���j���(Tѹ�'N���o����#��3�r���<D��a�N����qAU4tK�:D����$&G���@���cf�Z�,:D�$[ӍCQ�F=�U���r�(�'H9��6�S�g�? �谳F�	=�$��T�=n����"O,�K'��9�p�n^>S��p��"O|L��j��h�.����H2E��:�"O�S��Sv��"G��9+���`"O �x1'JZ���!e"Y?L�u�V"O�`�$��V�D�C��K����R"O����g�88I��R�Ozh��|��)�d� !�T+O�p�p��ǿk C䉁> �$�@�OYY�T��C�I�@F�mA��V���̑��D���mK���)q��SQ��'1[ƹ����oR:p)7'�<i�w���{���qfh�F��ȓh�&�I��Qas\���	6w�`��<	��)�rx�ݲ�J�n�0C^ ��c��E{����F�&���E�({~l�"��4��'	r���	�j�r҄�lu��#'l-K��B�	�^��'G� ���cɛ��6�2�Izx���MP�``��&h�v�T�>D�t
$�3s�|+��Gq5���Q��y�'�ў�'_�	p���*@�T��S,X���Y"�
�k�8ɩ&^?:Jmࣣ�%�hO?�D�?7� �cI�4#�1�V�R$D��y��	�u
T�ԣ�D���7�^1\�C�IP�.,"�K�.��\8E��˓�(O�b��$_�*v��p˄��g.'!��xB�>��O�y��Y5+rH3V"�&�~�C��:�S����Ev��c�8��*S"*!���������_�02J�,<!��1����⚘t[]KFc��!�D��3�&��B�S�?�b]�e؃k�!��t�ܚ�Q�|��P���+,�!�d�:́kժʵ7��`F�%�!�$�-~(qT
Q�!$��:�!���H�����+L��ɳ�c°B�!�d�=h�����N�'����'i!�$�-�.��ύ&P�� GrqO8�=aN<Q��D�)��t�2(��x@�o�]�<)f��8Y��X���2%ȵ�XY�<�҃\B����f�S�E��#!�O~B�'�,y�f���z�*� ��N1�@�
�'e�-�-I�|�hh�$��,�bA
�'ɊYB��=!�Y����Y�V��	�'�DHj!���o�,4ˇ�֥QA�``�'+��ㄫ�n�y��	@�|��'4 ��ش+�duI2��2��X�'�$B@�ݤ"�V����[ W�&y �'W� ���O�.r.����S�M.e��'4�lDy��I��{N�P!F0 ܀�3	�9�!��:�y��'\#5�H�`��P��	m��H����̱~�h�2�S�M� @�"O
|��˄�^�@��ӯ9֦=zƒx��'2��V`����� �ѼX&���'�]����(�<�c��"�nai�'�X�B�2��M�#���fa�y�O���"�)E;�Q`�#��Xu/ۥ 	�C�	�>s��S�^�b�8R�F�i��#=I��T?��5���1H�P�"�NZ���5D��8�*Ùd�2�gG�2u���f3D��{��P	UE�d"v�لU�(�iЮ3D�hJ�!Έ+��!X.41��*r2D����ގP��ј��ӝ;��IA�b��&���	.�J Rũ���#��J
<��Gzb��$�V�J^�P��,�7�b��#M8k��O���5� He@�)m`���gY�(.u���xܓ���� NP�q��w����Hԅ>�>��a"OZ�qT�����g�o��	h��$4?����>-�����@�M
�!��"
hH�l˰3�)�A|ax�I�f��
W�P�GID. ����*ʓ�H�`dÎ6v��<�6�A�Y�쨕'�ў�|BCn�U."����	-gpڅ��Y�[���O��x�L�x���1pC�J��2�yr�'����v*A1I"��b�&< ��'C���7gćdZ�Z��J?)��H�
�'{�0���شIi"T�F-@'���
�'�q�Ѯ�6 jA�� �Ď_�'�ў��h�c���0�޸
ԁ�}��H��.����X�J����܇]�h,��a�>��b�[#r���㍆D>���F�"�qwAE�9�Ν��Le���E|��ӪL� 9h'�Qj�q����V$�B�	&0͊@��cW�(RH�A7hث_�f�ɷ<�Q��}�W�Ǳ,�^@@�-�R<r|��s�<�FB�/f���� Vx%V%AW*�g�<9�D�C��	�4��*93Úg�<Ip���\��h*A�\ �(@�}�<�%�$�	3�	.���r.
n�<ɑ�F6Z��Y�o\�F��S��m�<9䑞"�<�â�O" �����j�<хFK9_�n(��N��#�+F�_�<Yu�ۤK � 9�O��^e(�pf$e�<Ն\3�����D��I3ՎOi�<)�@�]P�=i�F׿"ɒ�
!Hg�<Ag�N$,����n��J��tR�b�f�<�+��Ik�D/Y2�9��ۦ@r C�I�4�"��pEO-��(�DT�7r�C�	�@bp0[�����x�E�Y.�C�	�+6
\���O��\�T�K,(C�I��0��%De�����lKZ�B�I�)<�D�;v�`�#LƜ9��C�	�'G���F�	�8�(���'p�C�	�S(
�� �Vw��T�"�V,�
C�B:�B���5�3Ҿh��B�D+�cd�t�f�ԪPߤC�	*,	�` =dq�t� �NK�B�ɶ	��A;sA�$Zf>5�0��$l)�B䉿-W�����2Q
lQ[Sj޻��C�I��x0���q�|�vA�5��C�I�8UPH���Y71����nu`bC䉐j���A�gJn��Po��,��B�I0c��L ǉ0:�:]#���r10C�$�p����h��o��3*C�ɀ��1�JTw����
X�B�	�(d!I����(e�K�#�xC䉐��T`3�H�u��{#c�/>ĨC�I�B�lp��I�*a�ɳ ��C�	1uP.��&Q*�"C�C�I*`j:��e[
|,�����C�"\�m��W�p�����ѨAd6C�ɟ;�NT;bH�)���jV6?`B�H,V���ʹ��3�Iq
���ɼKu"����+�8�QT����`��G�Nf`Q�C�!\E��'��,	C"�k��[#�1Loب��'½Q��13��|���ŹA9��
�'�Ą�K^eb�j�k�>&H�)
�'�ڹ�2'GYaؔ��M9�⥋	�'�*�3�mM}̖�j`�E%Vmd\�
�'���I�.ٻ1��b-L&I@j�	
��� R9Fڹn4��W�A�����"O�12̓�ajX�B"XMg��b "O�x�k�$���)��{Z,L"&"Ov8���۶kh�ī�cʖ4ʭ��"O��&��}k��k�CѴ ��8�"O�AY�����A��<�y��"O];�,�tJ�h�W�rR�B"O��a�"7���xDg�7&H���"OZ���J԰b�t�j�l^�G~�"O�郖�+YPp;C,�9�|`��"OfL�悮�X8H0E� z6�8!�"O����	>S2�����uJ���R"O�р�F�$;��b�3Ax��#"OZ�:d�e�&L��I�22Α@"Oʔt�" 4r�"\�-+T%�p"O�x�a�+dQ2����%/��u"O�e3��װDb�O	�/	Ze8w"O���J�-61Zs�SWL���"O6U��$^D�B�0��(%KB�{"O&\�E
F�Ȉw���w?2�ʰ"Oڝ�$��5b`��Ó�ˉ�� "O�E*q�A_��!t��oz^Ų�"O�p57l��a��N
}O�)ҧ"O:��i�1)
�&��V|��"O�ͺ��Q(LT�'G���D�R"O���j̓+.�(�qHT�	 �}ɠ"Ox��璮O, �3�B85����v"O�����K�d�x��`i�4N�x��U"O6ݠbƁ-7
��dg��+���e"O�Ea��ܙ'-H��+@u�Da�"O��j�IDJ������.e���"O�����85�&�b3��,O^��9�"O�xS�$ˍ���a�>2�0��5"O�[TJS�ڥaJ apM+�"O�����C�5ΨJE�K�6ḵZ�"O�2��!��0�0	MSZ|`ہ"O�i����36�i�������"O>Ѩ`Ô|��01�J@�p�	S"O� ���!h�$p���9��BF"Ol�IV��r�8�	���{�Ry�F"O�챷GRV�n`f ח�Ƅ�%"O��˵�V>$�J�s�R�S��	��"Oz��IH)�a!d�9�����"O�EӲ�h��%4MZ�Y*�J�"O�D���Q=,6eZFC�=�����"O��8�ˬ3���Y���D��"Or-�⢃�>�2���w�f���"OBŃ�t
���ʹl2~�y"O0�qjқ?jve��'�+wO&IR@"O����;%��q(N6<,���"O�:5m�SfLa��uA�"O쀻t�Co~:lK@�W��)�"OnI�$Q>M}���v��V�D���"ON����'��H���
"q02"O 43Da
?ix�2gJJ�s�=�@"O8��� �: �8$b��L�4�l �f"OP�8P��E/���'�O	=�J`B�I��#~�Ǩ��P-����FL̙�@�m�<)��G~��`�b��G��<ӗ�Th�<��N�/m,�@{�(��=�$����q�<Yv��$A��}� �g��Qs��V�<�2iI9pt*!N��w/���'�L�<�&�(qzF82&�>,���B�M�<�0��a�v�7$D�y3z�P�+�a���z
� �0Q 8l0���8$�LLz�O�o��je�'�U5܁�C�l���K< lD���{�	�,J����f��o��סL���O*�G�tc�w Q�v郦Y��sC����D[��p� /��S�
��@4�$U1V<k`B͐1���DD=I�f�pN>A�D˷>v�i��e^ xw�D�AՆTL�t�Cg��|]��g��S^e��O�Q@6���n�'B&Hđ>�7M;�DH>�OC"`�a)��s'��
|lR���� *��s��9tFL�藆��HH<�Ɂ"G��;T���lN�LX%D�5#��'��:*BA��M	%z�ߢO�uS�Eª!�	�]�I�����IL?A��Pf��"L{`c����T?��KJ�N#����L9np��H�g�(���BXi	ؼ��G��A~�`!"A�O/���6�)��7�`��U�U�n6UI�:u��m��	-0��s�"M�$��U�V+O�M" 8�0 �3r�XXq�I\�l���󄂃	�C�i�T��g��d 
1�fK"���k�v���'�+E��Y�$�� �>�O�:���N�U8-[�P�X<�P'ǝpA��C�U�!�I��Prx�E{B���DK[4����N�4�|�;f�X�C��С-O���!e�5�G�es>�3�M����16�Q#���d`I���𢃯�Gj8�ӄ�Q����DҀ&Qd�!O"E�h�q#� \N�&׳Y�$�W22(Х�Лd�d�šO#��O�0�3 ���,S��c���<�Z䱴��!��?�G��� ^��Y��װp{��Vlm"�䁍9d��tꌚP
� �'qK��CI�C���!��Phe*�'9f�⟜��*�x��b�ؔ �o�؈!��;d&����I��~��ir�3�B��� �ϟ.�p�0�GG�GzXm`#�\�"����OvLX�'�4p���䆗~�BM�+��e92�%d�u�l�I=Y�-�!�/%՜�f�˿f�"ԃ5a���Rb�I:�y����
���Eg�)	�$0B�F��HO�[���M?�����L�_!Lő�
�����G�}��P�-O&(v.I	����dܶK���K��Ȓ9Vv\[ �0���:��'�A�$�\�B�ĕ':n����ӳ�Ґ �͊7@�dPK���^6��э�I�������SЬq��G�N��k��{�H� �2�n��^���u���3f��ӱ��(_.����
OpX���-�y2�͞9�� Z�KP{- X#&N���D��_�h�3�i �2s��Ӻ�<��9+O�	c �3jn�5�6hƸ��'��U�`����PDڱ�|��G�:A*��խבC���Åg~�+ۮ'���3�U�'�@뱏�/X.��֨Y&D�$�1N<!�s~�G>G�d�����gʘ$�N	���+:9b�
5m�su\�z�J���?�FG�Y�&R�)B(Y�� {��$�O�����Y����jȱ��RU`��t�R�Pd�'sQ?��e�	��crh16B���}ӎ�I#�i���c̍E�S�O��ea��J
��(���R|½��O��=�'"���O��`T��!�M6h�o�<D�r"O�����Y�Ba$��? ��ܙW�x�O�ؑG�)�E��6���F���L�n͉@�d�<��$��˔���$��mMXDq'�#hO��p�{���4&[X�H���wZ�T�A���7(�1
1������0<����O\S���9(�d��n�
�
��g��h"����>�Om(��H|�	�:��|���PO:t"H͕dL��j���"|�v*R=o6xqtn�&�ZY�%��<�FC �D�xP���<�Vć�U����B�8�X�� &�i�8�Z��i�9�V���fL�nMpX�ԅJ�O؝sb��(�Jp�+ǁ�x¥J/O�L��g �a 0�:"��?����į{�'�j1`&i�
Y�xk��d�w���7"�+ ($Z�6n��	�w�'WB�6�I>_�ơ0�Eo$t�a3 \�n����]'�"a�Z_g�I�_�­(�k�n&v��<���*���*.�m�Z�P-u�ӟ�XK<�El�(&�z���f�*kr�7�[�Y
��X��"[��U�M��Fd&�@r%�Rp*����x�n=pf>$A��і��C�9�'I����l�2�S@/�O���np�Xkd��{�aP�lQ�@��A�
tPJ|:� 04�$q$����F)rYz��+ГDe�͹!m��>Y��W(�Ms��M+����W��yG�5j0�D���&��eAP�p>1ܴ�R�ڵJ�8�n�֚�(����>@8�d`@u�l��P-Ɉ`�l��j�7c��hKD KG+�!��ر/&�H�H�"'�-P ����3�j�Y �E�  44Bbݰa�Z�#�F�#M������Bc7�ѡ�%�>q��E�^���$,$�Q3�|J?�X��O�N�>�{CL�5�ɒͨ�pnZ�6�ʌb��@)Қ�4%�L�:��B5',z�HUB�b�&|��W�ڌVu�ܚW,ԥ��I��H���?L P�F�`��`�3J�9Tԣ���'@~�#�H	;�މy$�SV�	�X� )�Q�Yt$I��[�+f.6m!F0^s�K���<�"�T`�? Q3�D.Y���A���*}��c�Q0�T��%��F͋��=|��u�#.ު���ߏo����v(m@��Y:�0<q�`�/P����3�Ɓi�o�pV�lc��0=(�e�
V(�{���*�����X�Os�}+Q瀽)( i:�'��Ԓ���OR�$,O"T�;G�ϴj-��%%��%m��8ۥ��:��Q��>*k\A��X��y�OҬF��OpQ2��J ��\؀/Up�^�"h&U��,���R� G)�F�1�P�O��9��q؈ 8N͹h�m���R�D�A'�	�0����\S����e���B]l d� '~ୂ6舾X�%pd�G�D�@h�'>�	�i%(�c�U�@F2�,�%�`��f'H�b��p<��m����7{�X�F7r�ܱ�
�,��IAEW�i�v��zw-��j��E�$l��!1x��M,8@4ʁF���I�Ys�|2��2zE��d�Əb�>��f�GN[�!���A�$�P���H���qO?�ɥs�ȡ�5ɝ�,\݈f �A
DWh��\��I�r�'T�P$@�r�̩�%Y>�	��yw�+S�!���9z� �'����xr�
X���0���K��=Ӗ	\�`|��뽟X�Տ6��d֮u5���vAR.��'��}[qk%n��׃�l�N��ϓn����n�H����|��A"q�J�����.N�))�2�8O�\�`mN0{��̳��1<O�t�5ܻ��A�>�V����$
P(L��D�S/���?�B��#�M�\wJ9Be͍;���S�
�E`��44�(�C��:� �ٖ��-M�µ	db�?%ڥ�K<yC(<#sP�#�^%��'�yw�_�TղUɓ�A�Y��"Ɋ7�yDϜ&Ǥ�B�ȃg�D|�eHŏ~C��9��˫3�(�X6Z�"~��@Q2�l�9%�ܭ��l2�0A��M{�u�pNm�)����\8iϓ�L�&J��
�R��	ϓV��H��/�b���q���jQ����	~ix|�R��)^Z,���C��	��Hb�FM�P�nh<a�I�G�� Ar�[ ���e�X�'�"��S���Q��ɔ�1����_jH�,c��׉wh!�d��Z�����:"��@!M)R�ܺ�X��ܠ��>E���q8X�Y"BӒ-����ҊZ	Mc�цʓ\@b� �(�Q#
Q0gK§���O͐*�!�n��́,�b�3gӾr����@��"�!�$͔n�X!G�D�c��H`��3@}!���_-����	N�/p�xN�F!��!����F�&_�D�@��E!��3T���BkKAwDR�`/8!�d΄o.�C�R�z��@�O�.)�!򄟗Q#�!�p��0/��Q�6 ��V!�$JaR@t�MQ��A��
$5!�ޏ9y����/X�`iflK�.U�G!�d2.���*gK�0sZzD�g��'*!�D��R�}:e�A�������F!�ŵ�.1�4f*�*��Sc>]!�d�3���o�,�t��#O�1�!�d3M��8�+3Y��-
�'�G5!��n�i�(Z�F�}1�S�^�!�*gB��q��C 0p3�h@�!�D�U�LJ7�T2`8�S%�Q�!�D�%��I��BS >���+ߖ7!�B?pQ|`S��@�r����e�5�!��HR����j��)֠���K�!��!Kǂ\�p�	��{�CQ!��Lv�����E���PC���&ں��5l�8v����c�	�y"���e�H}�g��R�H�����yr�E�{��P�dQ�K�e!��y"@��c�4��i��EB���S�yҠÕO1|)�`�+`e��["��8�y���>Ev���r �HF��J&X��yb��5=���q4=�L��`�U�<qTY� $��
�K�XFH�Y�<)S�7y�4%+�;lz�2�EW�<t�Y-�43�y/@�� �P�<��
g8��F���Kȥ���S�<� ����"3}�\�g#�8{�q��"O؅PG)�7v,B����	��+�"O �Zy@a�ׁ޾ ���"OJ00GӇ\2��!oI%CŶ*t"O�p2�
h^�rP.�V�B4"OF���B�V/�P�sm�5`���u"O"��`͑*V���zf��0i�)��"OL���>s0��#+�![>DZ&"O<|�%P)^�l$1֔zA��"Oh��J�$pR�)zC$��"O���-�=zN����H5-bD�R"O�����ߒLt�y9���7j4{�"O܁ρ("P��#�չG,� �"O<2���Y�@�Qo�� H�"O�TF�'t����D�Qi"O�}qBH���ҹB�'�!8� �"O�h�7�K�A��ň��/�x �"O���gg݀by��ifŉ4	�9�"Olx�0b�jֹR`���b"����"Op��� �Ј��/<@��"Ota7��%��B�*�]Rȥr"O\�Ypg��$dEY#j
"2�! "O���&��i׫O�%"�QE"O��a�EB|��,�8���"ODh"t�X�D�j\@c��>8�0��"O"��@�S�<�݃��"O;���7 �(�����Fla!"O�tR�B�Zޔ����v��8d"O�M��lYCdp 2���cDq�d"O�C&iA�R�����E<�|���"O!Ka%@4t��X� �8-�p���"OJ6�P(%,��^ؤ@[�-\:==!� =�rYV��u(`��a�Xt!��
/�Hme��12$��%��l!��`J�|a�	X	Ar��2k�!�
�I�"�pGM �9��)q�C��
!�dچD�����V[1.��h�* w!��/:��DI��' 4dy*��7�!�ė�2A�G�I q�H%���?W!���0��t���}��.��H�!�$t" -� �.C�FT����f�!�Dׇg��aC��Ә��H2G������q�v�)C��K[�mJ#,�5Z�FY��+Ԫ���*�r�h-�ꁳJSpe��Wٮm�a�.P��j`*Y�����	Y�i�䍇�V��<r�c�&C��ȓR������ ��	�`!/z����y�(M+��Й_
(��ӧ�t���<�qW�O�2�ؕ3�'ɝ�0���	:�:í�)`\X��ǘ� ���:X����D���R��<xd�ȓD�f��pjO9�Z���JG4Hf�ȓ����GE�%piʕ�U�J���~��V._�F�<�ĢO	V
VهȓL�@�3)��z�����(� .n1��>���0K�1�x�dʏ;&���'�4�qC��.�,�!K�2�F���Gt��2�d��3��R��(:)����Kz|L��/0���"$�L�oJA����4S7)�*\����� ��ȓfjnp���2.* ]�GJ<~�m����0����Tz�Cc��'��	�ȓo3�R2�[�$���*�ʆE�r ����!�E_�i�b-+Vg�zK�̄�S�? `a�6�eZ�Y JTJ�(hA"O�a�#�ɩT(��	�㔲4n��"O|-�s�P�>>L� RBϤ|?$Ց�"O���'E����r��{���+d"O`d)TH���^��o�g���`"O�PpJO���$ '�E�(bz�%�'{Ġ�dAy�zezE;�BH�G۠䡅�l��%��F��Q);_��Aƌu��ݖ'��l���2.ɧ(��dc �
%Kr���GHp�[��'��l#�ON�ɻ@ ����)l�hW"�;-[D��!D �Z����f@�'r"L���$Fx�*8.j�y�%�[#�8(5����I�	B�%X*FX�~"���"��"�ɟb�޼�7H�'|��a�M ?���	Vj�z���y
�Y��=j��F%C�'ްp�"�-Wf�~M�y�v�?[��=f�$�6�C�%ܲp�����"��F�TE�� K��m�T
�+ ���Y?�obp��
�g!p@9Ə�׼���F��g��y@F��f�,��qM
��O5���Bi�$,^�
� 1.��k&O84YQ�ܻV���I�TX���N���f����e��$��P����0lZ�`I��]IX�ti���*U�HP���6�_�o���@�??�ō��zИ��ъ;}�����!Jڽ^�>1����82�����%�	������@�4��k=R�8��|�~���A�iK2H;��
AД�'��<� �@�241��_�t	Y��Z��Ĺa�1������S�����t�8�ca,I0H��~LR�2b��P̒q �5cC�R�aȪ�YE�fhxsVD G��Z�.��Q��a &��X0)u���#˿t�lu �"�[�
�E|2�<�tx��R�EX@�'I�D�"�?^;�E�Qn^1&A��!ψC*�����_��	SBDA��L��O:�Q�?��A�N��l�TL�Sږ���o��<��i̔N�p)���>>��{��x���?��ώ�j`S�7��3瀈
5f���.���|cP�_�q
����TUZ�Ц�eC2x�0'�o���6�V!B�R=��h�揪+��T`�͕3"&e�LA6i���et.X�3�V#4�D����Va~"�.R���`�'�(\!�fE����jp��KLĕ'c�Z��@�?�&)DRc� ��a�h K���hK��On�*ġU5
}�)O䑑ˑ�%��҄Bɧs�b2%D�?-\�9��-��?)E�M�i� va<���s�ǔ�<�V!�g���i�<q�چA)�u��G/�i��R4iA�g�51c��ʄ��!��7.Ir�L�!~I� �H�/��	�g|�R�1G�x��u��P�'�l�QT�|�M�'6B%ِᛍ3|���2�;�O�ۦ�566~�4�K�8�l`�����N�\6|�Uz��D��=�h�?�px�1�����f[���5@�h�'�x�����~�d_(!��8�%�D�v0Z4ǈ7 ~i��*Yh�A�@�hj&��.V�`��7�r�FB虱AzZ�H��i���!��͔K�B���-
|�!�I��bh�JT8Q�].B��I$��`4��S����A�Ř�1� @��fm�"C�I-]� �XѬ�(s��pbܘC0C�%">H�b�M�9n½aT�ܽB8���^6#�BxC1@�	�0 ��\�!�R2	F�!a�e��)_�uJ��_:����At�@"�NIK�O��CfcQ>aI`<{�+��R�bp��'�~ً���P�~�R�!�ft�S��n�,�v�ZN�"~�I=I,xJ�41�LH0JP�S�B��)!�R<�CC�r�����扣48�QPǟ�M���	���asg�9	��!���.r��D_L�X�0C]�p�DhRe�D�T�f,k�l�p�<�ҳ $4��s(��Y-��z5�V-yڱ�d'?�w���sgQ�T������K����UaHe��0AwI��y�Ɔi5��:qŊ�Q~رA��
6SfpȖ�.[�2�Q�"~�q��I�b�1o�uzת=)&@X��V����Ǐ1t�P"⊔en�5�
y~�x�G	&D*�\Iϓq:���ϼr�4E 6�!-�Ԅ�+B� 9!�G:��Y Ō�DJ����o���`��\h<��CM�uR���E�(iQR$Q�'K���eG�-�\���iNk� �ܼg���QuÌ�E!�D�Z,pLp����q�&B��5#�5�����eYD���>%?a�&j�DӍ+P�[�)�V�V�@��TG!�d]�� �	BM
z��)��g=�	kP����	��,��ތ��S�� �����(�a�fBب��hT"O�����ޠ������	?�`b�dJ��� 
;}�)�g}��,i�M�� W&2�R�����y�#�1hi��S�HT� ̓�xf��m1jo��"Hռ*�{�OM�D6Д��"�> �d5k����=�W�W�J�~j�/�O ���W8Ϭ�B��C�: \�B"O��D-�5@:�X��Z w,�2����H��|Y��P��h� D{#Y"}�<]��LC'����"OL|B���=x�V �'�n��H�$D%"Ǥ���,%}��)�g}RE��j�T�[ w!��RN)~s$C䉢O���F،=�������,g�27흴3� �1GP��=�Qρ)9,�U��'�����f�f؞��"P=}9�����'�R�`F	iJ���A�r��!�'��s6>>�� $chԵp�M�;�< ���S�i�J)jBK�*\� ��٨/Q~C�I/j�����@)yW�t���ڤJ ��N��YqO?�I�
h�ƪ[u�N�	�B�6b�b#=�7kҎ�dk���4L����aĀIz>!C��!��	N��%X���(��h����K$^��jgJ�I��>E���+���f��
/`�����dh���H!�1�I6��A���a{����Y�K���)ϓopf�S񥊞fU�÷�5Y
������A5<5�1� �M �Ha2옳S'�1��sh<Y��U$���6��/��3�@�'t-Pp�H�D����iN�J?�A��.L�(�������Y�!�$�-L �d�ʋ5��@�ٍƖ��A�L	���C�<E��'�ܱ�&_�4�r��gM�L�T���'�����˺8�\��cF�F����'��#H�:=jthA4�';4���_�l��cE���U�B,nMp��ê��B7�
�t��:7`N/$,pɉ?��xr.�7`"Ѣ���bS29r����Or\�4��]h�\�e�?�ӡg
,���h&�����H8B�I��X}��"yL|Q)�OX�>����=-�����7}���'J8k�/�<U���c�a��'pH��(X
�Z���AP ^�mq�OX(���>� ������:���4x���R��9�!��i�L�s�(�
{z���D"�3!�!�D���	���vu�6�C�7�!��!{�R-y1ǅ|o����T-Zx!�DQ�m�T�JU�Z�*���� /�53�!�d�X��C�'����1匈�Py�[��Q����:R�4h�'����y2#՚ɲ(B4�ɕ�^e��.�y2�٢IWp�,Y3����ȭf��,�ȓ}ƚ��D�@�|��uAͳ2H��z�2��w`OX0}�d�+IPhp���x��',
Ӣ��*� iæ9�ȓUR���eO0���"Pmˣ�B��ȓ;`RĠa܂h��0�G�ߜ]=0���~C��0P�� X"'��N����69��X�R3��"5MK26�,|��*b��ǭ���B�b�C�h�L]�ȓ"�<C�bE�zEBtbpl��.vQ��
�ʗ��&"}%���4�N��ȓT�L���	�����I�'����ȓ8�, �bÚ-%��|��P�-����ȓ�p��bj �;�����X�$���Kr��̇F"EB׫�YX��ȓe�P�r�:�H��g�N�L$`��H����E���x	�NQ��@�ȓ�BQ���v�*]��%l����@m�m�� H(!����U�н�ȓ`�]��lĉ�������d���3`ȼ�N �7� ��r@ƒ�P��S�? ���6	�9��`$#W��e� �'\�`�AK�By�fEB�f��q*!Mp��S�L��E:�)WH�<9c�/O5��T�L�09܅Q�l�<� ��E�n$XWD�Sۖ����p�<���AS�X�P.�[��C�,So�<Ѵ�B�"�D���_�t�h`���q�<9��L?/Τ[wGT+�!s�
p�<1�ƚ1>�	�(�2,ܝ��$�n�<QSGP��sp�ZV7^��)lܓ+���'7q�Q� �΂a��e�����L�c7O��?9��^�*<"<�0HT<t�� �~M?��F�Y�kb�]1ɈJ -�I�:j ���f6O�����#-���'�(����'"�"��D#.tc��WG�>�u����x�;#Ǉ���	6�'�p R�Ǭg����P�I��a� at��7Ɵ.;չ,O?=��+E��:B蒂=:���%�ɂ.Xp�rd X�!�&9�'Ja��T,�"��$n��n��0�t%��@Ւ@�B+K���)-L��}�K|҂ǰ6�:}��i@�@�I���/LxK���(t�:�=��5Y䨈�m:(+�'�$]Ho�����C�Bg!�Գ$!�ú���Vq��&��2a����cc�`�0Pg@lF�83�ʉ)�M37L>����C$ �
:�_:l��-���+��%�޴v2����);�>����$P�'��9���d
�#s��Y�O'{�'C�T�'*��b$l�t�������wj}��R�G��Q��}������L0u�TXxB I1T�ޕ�'��������,o&�Z�'��&��a�G����3<�l�<�{�'�h�b&`+��@�P��"��'����������DL�Pa[
�'��<h�����l��bD�D"��
�'�x�@�OĬ,�Q��K�8>d��	�'[���LM3�#�AN�-z��9	�'>V�"m�0-�mjd(�����'Ů��4�B�a�:M��͖L�<�'���� ���*1���E遶;|غ
�'���§�#��J��`�F�	�'\ ْ�LM.Gj� E��(WT*�'-h0r���.�Z1��B�`� �'�^��Ć�b�X�
���w��0
�'�L1�J'z�$@�r��x)�	�'�a ��@*u:"'�+�1��'(d)�T��1C�
�A�Y5l"	�'��Q�oU!e�V�),̭1b��'6D"�l�_r��K5DZ;T5(
�'����J̹R�z�+d�G�^���	�'2��񤅾}����Ȳ�p�R�'8�),��I�i0�W}Ih�"�'6 �!���i���A��?{l���'�D݉g��$Qi�}��N��5�
�'��(zEG͗SM��aLI�6)��S�'3�̊�`F55�pۥ��*��
�'�%��80��j�&��
n�!
�'t�ÔGNu��p���2S�x��'6�Te"�t1���ꃄ$�J���'Z<I�j�
i��|�4N�04Y��!�'��� � �/��H��#^v�+"O��v`ף=��]j�σ;	G�9�"O�mI��4�,K DE?`<X�A�"OԡS�L&2 �Yq�̄^A� Af"Ov�Y`��r�n-�a��&Zx�"OtU��a�xM� ���I�U#��1"O<�`E,3����\6"��"O�<!�"N�T�T�e <���0"O�I��)ΎO-:h��d�NX��"Oh��d�Z�qej$�Q��/*
�W"O>`���C6r���bU1����"Oظق'N�DV�zU��wm4 pd"ON�k�������܂0��L�G"O� t�:eɖ%a�a�f�(s��|rq"O��9#ŀ\���$N�+�����"O<�b��O�aVʬ#�$�	��d��"O.�q��ͫ%g����ޘ{j��8�"O��Hf��^��q�R�|R�"ODM��GH�8��g�ޚb5
T9E"O
݉�JS$j��	g�ْ��X��y�
�]lLkp��(G��E�`� �y�b÷�̽i�̎-9S����̱�y��:i�0�T�E�gv\�DO��y��Y�����Q�\�+��L��y�HňVO��d�Li��C*�4�yb�ހ)��4	���Es`ī�h��y���Z$�3�ʬ8 X���T/�y�* 19FH��m�h&����y�IM�F@X �QP����&�yr���XQYE��)^��ና��y2�F#K:d�叜%����^��y�e��7zP[������ ����yrF�t;�xm�B5�a�Mȳ�y�U!9D��V��%g��!��$�yB��'V\D�A���`�Bx[����y��N�wo��E�6S@VP�R�	1�yB�@
z찰&T;S�8�Ô��;�yRiԻ)�xU"��I� ͒U��:�yR�ʥp����DL�Ji|���d'�y��y1�qY�DW̌Y�o0�yR"ۭ=��͘���)L�Nh�t,��y�a��ULСo�F#�X�s���y��__�$� �^C��R��-�y�F��h�h��G��N�B$(��S��yB(Q�p��<A�l%F�Rl���Ә�ybII#}.���6��@P�5S`$ۂ�y⃗}L\I�+V5����
��y"���j��b���
��ĸ�yҊ���hH�3m�K����6�ٰ�y��JS�D2�H�*>:PCFGA��yrG0�;�
�
t����V�yR$ș���wD5�<��*͉�yb��$�Bѹ�ȳN{��5��!�yb�?]��I;���'K�2`�5B�y�(X�!1r�k�NDJ�V��)$"Ot�!�(r��qe��4Y���J"O^E���K8&4#S�M9.�b�"O$;k�}0՛5d٦h�p�("O���d�^yN\�ʞ8,�*m�6"Or-Ӳa�7���[U�
��uA"OƬ	��ТNδ����f���F"O�pb���T�T��)�a~�1{D"O�xxt�́p}nqdH�"pt"O�H�t.�I�h�cBƼo�>)z�"O��a��P5%b�	`��P�W��A"O��#c �G�|E2$��(�a[�"O�T{�Ŭ`F8��GZR~��$"O��s�ַa|2
S�f~�Xt"O,����H�R�~�2V8/�Z<��"O�Ң�D�Jq��Lu�
�g"O�(��U��6E���(�b��5"O~@`+Ӹb!��b�)��|�$"O���g�Wau�X���)�����"O���`Ș<[�$����(-��%f"O2����/S��QrWM�8�Hs�"O �P���K���G�FՌ�;�"OX	�Q���l�n�-
g+F�	2"O� ���t��8`� �k4aX�i%4�&"O�ZW*��72�q�͖+FAr�zq"O4����!_,�욤��l�`�0"O�Y�5LB-AƊUI6�<ui�"O����D�'(��F�ۖZ��cG"OT�Bcb�.,Z��s��6���2�"O2����#/�� { F�AԦ��"Op�:rیT��tłJ��T)ID"O�9���!?�0%�@�-o�~]� "Oh�ړ�\�L�LA�ףR���e"O$�a�ҥY:���@�V\�s�"OI���F7Dr�H"�6,P�X"O�Q	Ul�R��1�
=:=
�2"On9YĪ�,TX��b��F�
�xH�"O4��T!6�u95C�5�f�C7"O���6�� \�u1�D�	���!�"O^�Xs���2�*��KXW|�a�"O�a;��
��L`����u�� "OȬ᫝|d)�)��%���b�"Ota)c烉^7��b��˴S.d,K�"O��`K֞*=)a �̠N@8�"O�Mz����F��T��"O��ϔ=|�$��.�VAv8R"O�@�ت/A��KVϋ3bΤ��F"O����*ʾ@v�3�#?��@�q"O�u:!�#R�t�"�dS*T��͡ "O
��&�3E�p4�B%[u��Hb"O,r&A��Uޔc�Ԕe��d�"O����]#j���7��U��"O��b�K�;^f@���3R�t�Aq"O<T"�cҕ&p�㱈��]�^50�"OXt���*U���U*\	��}HA"O��;�H��h1J���q�5p`"Oj�p�J�����AW�sb�7"O\�5�%Q��sW
^y�d��"O*����'b�D�p��Jq
1S"O"LY�.p�D�i��^�dd��X1"O8�p��; \��ON4BU�=��"O��Ӡ��kp��A��G�u�u"O��
�FK�i����RD(�S"O�(0��O*���Z�z]���e"Oh�b� �"q�!�E��DBC"O��� NE�q���[D)%���X3"O��j�V�ҥ�.1�f���"O,d��B� '�*��-i��QF"O\x1�˞0�XdJ�Ҹ>60!�77
8�q��.Qrh9[����\!�<L8�����.y<�"�� !�E(�0�3!K�B����$B��PyR$ݎ7h^m����=Z;��b�&Y�yR	B�LjE�_5[}j󦉄�y'�&6 Ieㅇ$��9RanÒ�y�R�
vf��ՠ��H���� �y2�%3ZZ�҄
[/|)�]�&�;�y�SmB��@O�r8R�녀��yr�Z�|��1��D�T��сr��yŎ}���9a���Ωs�,���y���%A����0,�q��;�yr���!r��C�$?,�84c��y�hS%����ʏ�(��I�� �yB�)s�f�aRn�6$Q�=��솴�y"kA(+�^e�tk�"�rL�Ph���y�b�;H"�q+D�n��7��1�y⇂D�lI{�$�354<飶��8�y
� ��k������3υ�\�0sv"O�)��;)�,�R�K(@mМ@�"Oh[��C�gzM���_�Lk:�J�"O�(��܇X|�qKǽuk�ɻ�"Of��랴&R6�H	���"�=D� � iG	H�N�����G�����>D������mN�6Z�Т��<D���bF)}���a�-ĊC���4:D�|�_h��(��j���O8D� vh
y�4�3��]A�d��8D�Xb�  f_��Í�\�0�O:D�x�c��p��9e)��F�"���M+D���!��?���D��Lw�P�A+D���U�ʚ�j� ��ĚE$��jFL3D�l:1�'<@�f���C�C3D�Ls�@�%���pGaA�#üA��-/D�(i�*F �0<���_�7��}��+D�4���v�9fm��bF��3�(D�(
7�%u$PP�0$[�d/4yv&D�ة��_ ���W$���H@#D��h�$A��N<S1N����t?D����˫=�����+�h�����.0D��R@��M�M��璞
�|URF�"D�D��aM�"���1�$]�B9��`%D�(���?C�Q:�J�"^(y`m(D�Xyf-Ҹ>�8�7
B2`��ȩ�.'D�X�м0��ַg�4az����h�HB��505J�m@�hL��b�i��p�n��ɌDS :��B�5�ȓc�j�˗�"SS��+�&���Iɟ��BFW�f���ia ]�SM���<�EDk��&�O��)�4�����l�>��O���q��,)��V�Q�\!S�'Ƕi[0��	d��+�;)�4s4c��j6
�Bv/�"�����uA����	����Ox���i'J"�	z���}X�!p�H�`�T���<�����>ҧcRz���F�4Ed1��fɇQN���MS'�4$��"`�Q���x2����yoZ��M��Q��7��O ����O.?ǔɸve6F`b�_�.��d�O2�$ѫ>�X�O0�1�i�H��*�ǀ8j�Yu ��I��Oڹ��c� MR�~B�@��$|��"G� (�I ��o�s�u����0%?)�Om���b��*�r�#Ǫ*���զ:�$�O��<�`��/k2pA��<.MAZo����4�?��O*�����;�p�"��iRVe�E���D�<�Ok��'�r�i���� ��+�Μ� �W�����������,k��|ҏ_.l�@K�.)0��a����$K�DD,�(XR��U���@I�w�')~��m�P��&�iY��r�X�0��	ʟX�޴�?�;�g}�iJ�P�)�6I�4,�|豥�	,5�����<�	ۓ������Z� ��צ�>�P]�O
�	ͦ��I��P�޴��I�O7� �n���C�V���x���l<��6�ܐn�ϟ��	��<&��S�a�#d^�W�ze�!$W�J��0q�9$�Q��o�*�rU*[|y8Qc�70e�$l��n�@ :�ka�Z��0ƦZ+&��z�'M?cOȄ�%J`��\k��'%��|��')b�x�c4h-�Ǩ	�'u��#ɋ+��	SX�`8�BN�$�A�30�Ag��?�L>�@�if�Z��2�gD�M۴>�TujvB%R�,���,O�E@p�3�'G2�|�O&"��"d��'�6l�`�	�ǊH�P:���n^؞@T�F� ����0NO�`!�`�ÒG�Jv-��[��h6�'��];��?��B�K������q(���cW9\0�'�ҡǦr��O�n3`(IV��Is�MB��@�2a�<�e���3�����.�M'�ݩ1��X�l6mCߦe�'c�D���g�8��=��# M
�Q��ʟG� �ѧ��S&���ڟ���$L'����K�S�?E��ӓԗOH����M?�b��h��������i�n�O�$jQi�#>�H��1�O�^����}b�׮�?!��_��Ol�S�	H����U�$��!�5p�v�����'ў�n�7w�4٪6��vLX:0Gə"(�z��a�llZY}
� ��!jH�_Eԍ�fG,@��9��O>�D�O�OZ"=yeK   �