MPQ�   `�   p� �                   `�     ��     U�     �       p               9       �        @  ��)�N}�_�h�d����)�z�:b=����Dss                �tIS\�4����Y�"1�0�����8�?�H����:~����|�}B   1   �{���Xq����ʫ
���.O�X�.CW �< ����V�R����2�@     $@  Nh  �  �  �  �  ��  � V �3 AO Xj !� �� h���w8�ÀqdE�޲22�!{��M6){edf���d&DF����G�L({d�~��{���p��9γ�GTw�lѺ�z�W-��	��%ze;�����Ō^l�������~��?� e@\]�]u���g&Z�,�b�|�B�xgk)�!}��haa�>2Y�*"�y��:)w�n�2e���V~�Ö�)�s��TQxL᭛\�l+^A���ݺC��k~��9x2[h?�vZ�����5���N�,��PgL'����;1g�탅�d�*�U�2�_���'�k���Z�X&l�&0`9J[j{�4�nܫj�aa-"�p�00E`M�ll����Y;�+u&� �A�[�P�^�Ao����/��MsF���uh���D�����C��R���_�@1�i���H�����1՚x�3�܇��Pp�]y����2����}�6��@�����$s��ڿ���Q0ۥe�_�if��� ��l��1`M�����t���^��ﶃ�_�JTu�Nx+��D����"�T�?+��D �)E�u�}n-O�%@�Gvǯ��p�
C��N�yÍ��q�<�\mqZZ��;j�~�EY_�dѫ�Xڞ]U�c*����:�.�?-ǉj�)����ց%����	H0y	��=�$��q�����<l�����=��6B;}�&� 8���(3i��8MJ�~你�KQ� :8F{`L2�����F��	 {°W��xͧ��:�i��avү����c`e�]p�žY����i�>���N	v~&٭�7N���I������-���N�Eji6��K�,������9`x��MO��_�^D�Hק�cK�C �R`��h�ر�LB�R���H������qٟ�b>+�;��ϒP��Q�c�n�tn�xX��UD:�̓.�<"���W�6��4�����g�#�Ѐɞ�D0�#izG��P<t9�r�[���BO������/	�>���2�`Ś��-ND'����E���ܷ�j���=N�D7$��$$Xd����oY�3�����#��	^E5�nX&(,��I-���!���wh�b�5Z�ː"�Qqv�s�̦nN��(v�)�W��E�c㳘a�IB(Vc�ͤ�m�L�w[�Y'e�7zP�mO���u����0�_{�P�-P������(Æ��Ǥ�́�~:n�:�f�S,�>��n�~�,df�?���g;��u��_�Oz�s.���ծ]�858UŪ�J(�m����n�rO=	ջ<CŚG^������*M�b�픫�|�)��}bN��F���R��k��}���W���˧sN([��H��r� cg��m^&k?�&"ꁭӝ�%yb/���6yv*3����%`E�X,�4Q���Tw�������ތ����ϩжr�) �I���_ʲgpy1KR��;��\ҥϼ�5�u�Ut�����%���
����:*`���fI ]����#*�ծ�-NK������+~`��P�ر.������n�rKm��l'0Q`��V��VV9��!V#I��=g"�fݢ��lj��[j`N�la�}sf3���ƺaa�������5f�N��)��Ѯ��eG;+�K��P�.�Q*G�����p��9�`k��o�f�����K�L-�f,�5C/U��§�m3iM$0$`�a�A�N�4¬�}�,�Ks�Y�j��<� ��/{0��N��Cl!J_軁��<�?�r6�nPk�3&�b�E�b�
�nKӀ�^ˊ�0F`����_@':*`^��7���eV��b�Y��h�S��/��������k{��6���y.��?`�k7�;��-��Y�	^�F�ͰFzhւ�-��`;`_��E��+�������o�6��&[j�X�y�\��:�8�5#�Sq�+����q��F�%�#��I[�"�y;Ͳ�7r�_C�B4�7I`-����؟N�{1(��A�^4qc��q�i)���܊>稲C¥b"ʂڏ�Ft	{��'���݊�3R�|��Mgr��00 �fXفv��Zr��d;�OF�����-o�b(�vn�o��	zpE)�[G8F�6��$�u��u`Ek�M��w��|�D�6�Q%��i���z�ɚ��<���w�8��G�%M=�_�#��]O�[��K������|�!�O�Ԉ�E��r}�!4��<N0^X#��c�cNS�V:k�;�e����mt�9ʓ."RNV����zBs�&x���z��ُIL��XǏ_&\`��xH�Q;윁�̻�&��ߋ�{�EnƋ�Ls��d	�����;�]g������Q�����w����%��0\]�����?����j�n�m�\/3V�1�J�d���0+���X��%,ꇘRk�#�[�>al!lW�a�����7u�76��%t�^��D���c�����r�|0�V�&�4�mI��j2)d�{�c�P���#�#z_�9��@� LاC-�}������^��v�RZ#7X�.6��/�w��d|KC��~/�)�3�uXNY��_&�z����Fy����\ĲQ��XmJh�0G�X&0g`��,<���L"%������>���bN7�9�TDx
�R����+X��q�I�lgu��-���r9w�WN�6-�<��4m(�MeJC\���;0`��4����:+�ߖ-����0I�\p�?�!
���'�Zۚ�oM#�!:�Mh�"��)-�=�%)3���F-�Gl�:��ft�6՚��p���y��G4R��%�;���vx&�[߳��`��O�')�ྨ�����A̔���2�����q.�Sx�f<	0G��v��ckY��d"h}������'�nB�;\Y}b=U��}�M�7�zM͠X1V�~>a��G���[ږo-T�X����Qw�J�Y�x��D���|'�/`��e3n͸ګ�_tx��18�"±]\Ex]�>�,>7�E�_�)ѵ���Ѭ:������<�����N�>O�����@Ҫ�����۵���q���K7C���Lfc�m���Y�įB�>Q3�b�9tZig9�sB�)e:���f��?�h�.��~��S��� ��	,�k��wr�h�}:�u�F�7.�a�F���MHB��ÿ�#��nU_��xO$|�!����Ћ�a��3�,�,��b��|�e�9O�+�O�ٛne≍A� Y�I��W��#�������*��q;�q�y�W��s�W�t���6�����)Pk
X0F��iR@gt��a!�b6�h���b����;<7�+p[���p$#��X�MAVO�0��r���o�)A���V���ia�WNE����e"ˁb���o����r�DF�CL�	���ck�-����o-˲� �ָg��C�~���%�
,�H���#3�>�5xa���=��'D�ͅbv�S��ܕ����8�Ɗ%��=�bs��zf9����/8i{��݃b�BQń�R�E^�਍�rB����GvR�гٗ8Id�X,Zp�M�<�.�M�%����-�m�,��5�>N`D��Nb�}q�d��+!۲T��s�[�XK�^S���Zd�����B�o��K(�^P���,Iho����D���AW5�����H��t��*9
Z#񷭌�m>8�8#-ִ��@�fEC�a��ZK"��%ⴣ�������*PP�*�p��7M�}��G�x��N�%f�+�/�ф� :`A�{���t�,�όm������bB1��!���I�(��<�7�P�q�ů��(�%EIぷ�7z���V�����T�Ń����,ٻl�Ƹ}�;0� �a`����_]�Q?���:����?G_����M�b�\��84ÕV�<;�[f;�P̨`��(��ӧ��c9�
�Va@��f}J���M�;����U��Ϡ�����겧�o�p�b��h�����;~[��M��e�h�q�w/dU4�'�co�y��7a���B��J��c&�oPHhB1ɧ�R�W�h8lh�6���������D`�c5#���I����|PL�GV��b-W��J�.�:�>�	���и��Rg��.���KL¤�c�n���n��k����#-�M�1�*3Ҳ��c>�i�㬮���h��1D���6k�� �^�j�����Uk�s����A�̌��Q|N�WЧ?�աQT��brx4RX�%b߹]ȲsE��i�O���^��!GU�5)���W"}�y�D����(��w��L���Ŭ�b\�+"�2��d���b��ws��>[��9���Z$�[����b9krɺ����ғ�(V�{���Ղg7C#p�Y,u�ؠ���\�����ӯ�X)5th�<s`z���X�!�I�Kv�1A{���Zu�`��Ͱ�� ��cu������ZO��	��z���	�1�<���eLw1�1r_������&(V7M���8�����rn�Z��{(vc�8�W���؃H�!��P�2d(ˬRբ��f�OCGʽ��Fh�[�����ku���}S�;8��ϫt����0�#�[�&���a�7�筤�&W�z(�&�~%��u�?J�*�R��rdSUPM��Ɍ�I����� �(F�V�%E}�1�����5��	����O`WZ#n�q�U�kV�´7���c�U�N�:ߏyW������������s�Yk��$f@��u:V�!ʜ�R�'4~��r(���&mY��a�>�oNs��[32C&�\�B���*���jT|m�Qd�}�dz#_���C�v'Jv7���&�
N�$��[$t[�B���Ȣg�^0&�z����	 3 fsh�H\�n���%�l�8��>�b2�;gج-S��$,�	��v�k��:id��*J�	�D򏠘(y�r ����[���@k� (���뮼.�s�0���1��Á���c�ԏ�z�ճA���BFp�_(|<0O�p�`�����_]����'�ǩ�B{�!�єu��b���)�8���L�ٔ�{�i��`$�Jt�ǻ�zVd�[���X�QdS�P;���S(���.�Pl���ŭ�Ft�
��5a͔H0V��\��Q[IN��L+����o\f�c����t,l�A�AV���4̾l����b�y��vI��ŧ�d���(�B1N�ƅ�Word5��]y^�WŐc��7ыn��_tX���{2pB���.�z��T� �P��`�/7��[p,���^���<M�c�]�,OUM�7a �X�Il��rR��*�˻����v)�P��D�I!G2�`���]�e�.l(&N�wV���� X�	U���9ko{�:Wj���6�4��Ї�6��1	�nD}����|�m既g��1�PL�qb����9�P`���%�x~�ʪĠ�5y��/5�ɋP��iw��,YJ�0K��</n��r(��)���RX2��^P33V<à^:�����a"�� ��5���d��������t�y����FW�`��;����v�{?D�g��.D��*wU�iO�������cp+cuWT�SO�l���`��M��۴�b�51�4d��7b(5v��xoA��^o;�=q�������-G�B���.-oIċ�{�4~��zn��@1
-w��ML���3�?پ�1`
c�z���*�o�	�`������>�5l����`�����z3n)��(^:2W�!���h�N
J�G�M3�����Ţ��2��v	1�����v�j{C1���9�߷�xC�u���jPǜNh���p7k����V�=Ps��Kv�V�cEF�(��Rt�S��]�]s�޻�}��v�$�m�7dL�������M�+3(Ve�c�΀r��
�O���{g�C1I'bC/�^1�k<N�Fw�ʮA1�Â�&�,
���n�I������j��.��~��ݽe����شS�K	���Q�����<���w��L[+�jeý򠘝0>�>�>]���>�e�O�b��m-��b1ؓ�L&i���
���M�ۯ�5���H�u�<�B�<��-��&td3~���rZ���Y;nǺ�@���\tA�l�M��'4؝��ӯ��X�B���^{���]7��m���F� ?'Cz�*|&�삃���վP���Ui{gC��g��u6ߌT�z2[cת���&w��<�j{��Q�5T�TXT��O�&"G�U�#��_��m}�@�]�!cLze(�?�#4�ZxV�}�}��c;������$7\m��'ei���P�2r\�PP�\�Ϯ����s�?wf�G��-V��L�jjGk(F��K����d<z�XY��9j'�?��
4Jor��2J�YaEs���Ǫ�?^��ɔa�2�5k:>��Mb>�Lȑ�	L��I���aצ��J0�H'�5ze���ߣ��"��#�Rf�;����Y}�@�����$������v"��K������,!띶|�*�����9y��c�m�_�倫y�U8X�kO�Q��z�=Vzh�RolCh�>�
�d�X�=I.��0������B�U�����t��P}L�}�ԫ�΁?����jB1���޺I�S*��7]�+Jܗ�bb����H�]2��\��H�m�0��q;����'���.�Β�$ݏ�-���d����Y#���:4���V����s�o>J��D�o�b+͏f4[�k�5e��Tio%C�����2bcn2���n[��#5C�	�7؂�D�h>R���T�_
���ߚ8�`;�EGFsF����e�X_|S����mD��Z���O߬���A�Ū��"�����Һ��^a5]�M�1K���֧X��Pn�^�����E��;��}���y�O�&?/�ɘ�n9��E6B�F��&t�;���w��nf���.C�b��3�{�x�d8�F3�^_�׽5�
�!�j�!ķ��"��h��`���Ob����9�?r^}���AE�x+��v�߈�(�����Za�������lh���w<֍���J%!#d�̆=�3��eD���=�%IV����a�d�"22��L��}v~�:/�����|��?ˋ��:�r8��Wh���܆��E}����������2�����-���Kk�y�����|�۫��g���fCuq`�`��h�����D%ð�76T�S�8�v��,�ˤ������U������Ƕc8������g�3X����܎��DI�[M�a��w�O!�G���9Y�6}�$u�`�k� ��5�H��m��4#�Lb��h��9wS�ıֽ��a���=`
`O���q�]��cY]�WnQ<��z��o;����5�ݏ�έ/��9s�Q&oj;��=�s�L�D���{��S���}m�1��a���I�'/�ߎ�}{�f;��9zCQ������w$�i�Bo�̄{k3?���v|^�S�o!�r�sV���\�4X(��1n����Y�a?��eBN�IS.\ڻ�����?��OWm$<#N�n����m����V�)�E��ݮ(�O7�c��ɛ�3ks��DJ&�v��G�4�������.q2a9���d�ao�0~�������s�?��i�wtw��/ĉ�{F�_�"&����5ʳΏ����A���_�õ9)�i>����L[���۱�IR_3s��.���~���4َ=gPp�W����ٸ��%��c91��a����i^��:�K����L�U�ś`�2��7�� ��1���,�{p��|�˾!Ϥ}�q;F���q�Fe��Oab��ۏʿڶc��vֶ���b�M�*�����:���ȭw���=��a4���cRvo��R�B�է�V�ס��,b]�m���1>��R7��ȭ�)��G������c���i	Eۙ?vW��p��.�h��:7�ܩ�;G]Ųs``�����=�$4����CJk0T�z��ji>y�q^�\jy
Q�t��V�u��!1��?Y��/�#]�2�D�����+>���J�ʮ.Q����������	4�\�\}2���S님��S�?�S�������wY\v�F��C�[P�~�!��TfD�J�S�{�Hye�`�6u(�|M*����k�<�YH_λ!�OL+�B]&�+�FÛ�*k�TXl�N���{��o6�P9�;���E��U���t�~g�Q�I�����%�G���&�v�*�<l���!�2>/^0k0m�au���e.N�Iv*Oa�ޡ���K�v�z�פ$y�>�Ӧ5�t�ElaNn[w��IwKYL���'��L2�5g���	��w��0�5W�	�����c06���x:��;W-㻓W��}y�*)Jڂ���>��lN�X�˟)4�|�L:�A��
W��9���?_�^�%UR��t�m��R��r7*�7vws��R
�Pc�vmg%�ve���
���YbO�CCv-�7dݎ��]k����>�XC5����]H���y�!�N���i����e����YE���*W|MY���	L,1q�`̨���r�E����V����OT���O�U���HeT�����?�&e�x��N��������+VT����I���f��%g���K�kV9�y�ü���O=�8حE���eneUS�����Ӄ.���tq�.�Ͼ���6ͤ�>J��rrZW���1�+=U`2�)�_�w@w���Q�9Z��>���&vђEV��N�X�S�i��x����Թ�<��,-M����Y
;i,��]�"L�cN'�t��ȋ1Kf+��Z{A��M�C������r��\L���S0rt�T�[,����j�m��le$L��`t`��]r���'��/���e�J�r�~m@���������n��o:+W\������ybۗAy�3�~�;���eV��b��	�B�;������ꪡ{
F��z���169���b�Tv�M�jjq95P]2�T�nz��t�؝l�z�RSbF�Q���S�)�w��:k�͈������ �O�,����J�%�����穳s�\���/#f&�1��,e�U{xk�������C���?���S��u�\Ĝg\�A��oT�~rna��[w��+�^���忶���d�.R|y�M�>�9��V��-/�6K�,����5���b;6b������芣��f�*�*۱���~�4x&^�ڢu�b*O��w;F�5��Y�30�@JTS�"K������y���z�>��a����\� K��o۪3��JN�����bt*�t���30W�K��`x`�X��.D��(��@.�wV���K�c���F;,�O|���V�W��5��ߎI���ҟ��SI��|�W�ނ�۱�1q���tDE6����F䭷c��$���=�yǽ�ht!*k�G��>�4M��@��ޣ"�әS�_wd>eK��s��7&�e,��6*�,v��h��󏡺בM��q54?��Q�9��~�a+�yP�E��r�e�?:�;����e�}; �y������N���`n`OP]�JRM�D����f+�?�U���1l���$������⼂>م3§:~�?u3b��٣o����M�~�PXS~h�	b�`�`/�����`ӎ���	bYx}�їtz�.�%��F��Y��Mֻw����P�y���ׂ#�5�6Y��9�<�
��(�j�)�+dR��Mr���������v7{uS��_\e��4)Z�|~�%'��� �7b��Ӄ�T�?��PJ�L��]����wF�(U�[v��Y�����`��?����:��P�&�_�#� A�c�+��K*_�Z������S���c��;�:���9N#����MWǮ����^���c�Q���G��`�!�'FFs��E��2�ȷz��4�?6���)���c�J˭�)���{X��v��WF얟�|�������P����nj�Z����w����;�wj��m�籠�1�C������M��7�w��(��f�1�R417a�X�N�%Ƃ�O���
����+��yL�}�8J���(����&��B�1L�� Q����j����i�Z�U6� ����w`����͘���I��֗�
��v^̶�ߎ��ҚhV=y�P�,��da��/�m.�c05�"?��l���t�&�o�ws]NX�����?�ƶGH��X��
���M������1xK;���f��4�`�kr[�?�����\��+��H�?�ey�uڎ�I�(��U�v��I3)�m�\,�$�O��.r���ȋ[f��q;��ǣ��h��g�M��/��۱���ࣶD#O��S�o]��t;f��)�Eh�xG���ܸ�{�v|	۱ �������>��S菊�$
܎��9�E�rx�U���+:m��$5�M�2���(�Å/j�;eu�1��� �?M�r�ٰ��FF�fF��NF�ݍ��'ߚ7U�&���=t2��(�������q����{�^!m��t P�Ad��pBk���
�T0�P�`V`U`,`�`��l��?d���O������9HTu��D�L%0%0b0e� 0-0��`�`-`����V48lc�|)7&�<�t~m���L, L���X����ɾiט.q]��>���1^�5�f�&
���L���ܱ�8V�k�F��	!��� rG30<�,�09��`_����I��X��\ʽC���i!�e�b}��8�:X#XX7�� �J�NH�,��yh}�1�I�n#9/0Y��``�`?���e����������g���*�.�'�Y�+)B�V
&�v��l�6���Ϙ�'HߎM	L���`��L��(�X ��3��`
`�*p�����p�T6U�e���KZ�[�;+��8�a0&�K�ir��i��Y��B�G/>�� S3��	�L �X���\�<~5s�"O�j��F7~��q��"�m�n�<.���Ia�O�_��+A��H�&�c��%K_fA�Z��tC������W>�8r��,��>�m�[�e}4|��o�h���ص��4�޸�`��0+�F�����0T7�2����&=�7ԟ��Rn�#�� ���8�I����3j�dv;���=o��Rxށ8y>��&+L@����(KD��y�'���[�Y�\R�����Y0�V�2�I�`u�-�`$M(����Ϣ�j>�B��}R3~j@b�{V�E��4+��3��,M����`ŏ�mD� b�ڃ��:��Q��˃�K/��'����Oe��]��Ի��Lk-
cƨn�5t�FkK���j0���$s�]�ۅw	�~[�/�i�L���˧f����)�Ԛ�'�G̤mf����ԍY���T���7��?�n���#�P�m��F�\Pv�ߝZD�'�=�*�__��˝��fC��t�I|�+�n��9��M�b�3bv�A�|?c��؛�u�g_����h$��Pv�j��B�5{ړ���l'W�Ȍ�x�n����M2�0��yޠ���e�F��)|5�&�Lt�����P�l-�C�^�x�����	j��'��ɜ���UcV��x�>�.�X1!�!���;��BϪ�/��s;$��>{D�l��mg�|��z��b��:Oߴqn��_1Ƣ��>�H�ƲA�s`2`�ȋn����cҦ1<����Y�_^,2I�fm���}[�q���Yab��mv�|����o�4�z,)pS�q�19��,�LӉW3>��Ow
�URfL�&�I��(���ecٟ.����ʹ�Crvі�(ѥ�����H֕���N &][�oòw1�j7J���w��I7vW+�C�����������]S���D�Ӛփ��{G�&{�6��=w/����r���S��U~͏]������j�Y�Y�=�8fy���P���b?���'� b��%�<���|�_�K[�� V&&��,���5������u}dk������;�L;����]�QRAa�Nd�M�@�Y�C�=��-�`�`�X&��,2�랷��Q�U����k��ެ���zy�󃭎�\���m^Xƍ�'	������i<���,��')��[��Fl"m4`V`o�6��uOJ�O��<j�_�tDI-�X�49ѦFƆe�_�����$��}��M��P�
�%��!���(�kSx;4��7t,��mes8n��2�����z:~�8�_�FVf6�m���bEu쏇~�mi�â���dO���66���Eu7��%mOI%YS%RU^��Q[���#�d��DUTL1LB�/i#������3��]6<�����x�maޥS�Α�f<�,1w�&�6�p�t0Y����1B��m����	;���B�8b�`��:0�z+��s����=�R�OR��Fۨ\��������2;��#jS����e;�:�s_S��.W�������
�s���!fc{g�Y.�� S�EuJk�Z�� �I0F�*�W`5`��^@[%�zr���ŧC#�	�f?I󕁭7S/m2���+�G�{E��k�-�[ě(�~g	8I�CK�\�0���MPG������ w ��Ѻ���su{�t��U�Y��5�)��m�Cާ�).�Ly����|
&��������!��mZ�,U�X�Y(��u�0�K�>�}������
%��K�ik���Ƴ7��k$�����I7��;҂x�e"�Ꞃ���G��P������y��;�������%*�c s��t��U��M�| l���%ru����q��q%�7a�ss�X�6�jw<�~��X��]7N	�V��8�a�]���8��a:,�٨}�a�{�L�]�4��k��f� �0.�G`�`^X���_����S',Xg<90�Tx��ԋ�`�`�`��M�76�� �v���M�wX��1���v{���$��<F&8�8W�/c��\�q�R��0]�3w�{5e�t�����\4�B��?�%�8X�~Lw��2�*�!���we+�v����6�fV�ա�5���e�?��g>i�X_v!�)o��	0�Ic�A7�%t��:�\�[�l�ATi�<ÒSMeڳ��{'���,�����hb�$bg����<=���&S%��_!C���װ;>l?��0Ĉ9�Vv,���mfè۱���;
�c��ޛ�4!�BG݈��4'��k���9�O���:T!��=�k%b4{FI*�|��~7�	�c�� K��B��>v��ϗlJ��Kj��Ȼ�����X���3�1eTO�]d�v���?u��!�0�l�q!&��Q�ɒ���Vuf�;F�E�}/�*����{^a8��A�{�17��f���h|h!t��i��(�Rs�O(]:H����~�ˌ+c������$��{�JFsM8�NZ��)����_E�#�60v��X];X�~�۪]�_�߻5Q?�M�l�i�h+�2�Σ���~�}�oG�[k�0A�I������T4ܻt�cY:boeI���Q5���{�$C�v�,LL1�8�)���22��ѐC�0w̰�͉�^�AHF�&�ڏ�|0s0~�]�	���=f��X��\���O���G�X]���J�h��Cm;?��uSG� �X�Jص6:���Y0z�```j`\`����8q���z�T�R��2�候�}�D[�)��M��"l�lKe�>��۫�L��(b����k ���i��W�ci�멼���^=6�T����z���R���m�X���+�{ v�X�b�Dai�1sH��S�]���>�w���f�V��䒌4��<Z>��{��%
�7C��	m�	��䓌��ڟοt�F���=�i�Rͫ.M��s�Lݎ��Ø;tkӓ`iyW��Wq?o�ê��\���߉W�b����= +�k�����ve�����������(փ����16kT�d���&�ze�#W�F����9I+�?��xI[��
]��]�%��{���̅��9��s��=ґ�<5��R�֢�E��^���1]�T�Q��0+�5L��`���nX�a��J��<k^
�������ʱ:��t�(���}U�A����Ȫ���r�?��6�Ubw�T�gd�G��I�s'�?�0K��$h̺�U�I�z���a���c�/�P]Ѻ[!-g�|{����!��ع200W�}`b�)ˣL�L�ښ��C{ܾ��!���P�A��M&}m�`�`���޲�^�NN�����׫�k���n4�-e������qT���yB������/y��8�����>�U�-���ml����<���d�Ԫ����=w��Ʌ��		G�y��&�N��حtfx��Ā�W���_l��(��r�]ޭ.�\GQML�1�Z��3��Q���ϲdV5/�Z���}�G�r��K K;&V6(x�ℬ�2�B�R�w#C��m�``"`$X]$X���%&Zi�+
���U�E��/�]C[�)�e�ʢ{���"�ɧ46�͂���R*��7�>I��cRJ�	g�(/b�ČGN&�4]r-�^5��j���b;�	�6F&��{V�Q�I�ř�n�q���ĩYY����(q ,�y��a�h@[QU����10��
5A%��Kwt��k�Y�:��1��Pc�%�c��
t���U���f���^��">�8�,F�H���
,�
L�ssWX^Q,��`hSi� "�РM��Vv��m�`�`k��Aئj���{)�시�FƷ�
b�j-,	�tWw�?$�1>��w��w��%�gTW�_��ϳ�\
Q>�3DXF��[��s�e~�X�LOg�\p.���ӪR��5b���6 F����PS-��)3�Ҵ`�G,�4bg��IE�c��̠/OKVq��k哢'���2���L�8Ƀ1E�-�����2�>_1y���W��+XT?�i��;vL�{��Q"X�]�ꈵ����Ǣ��+<�|Y$�~�����rd��u�m#�.N�����c�?3uO�p��>f�����d��	Y��x7>��}:���	����5s]���~�u��FL��"%�S0:�Lw@Ý���¢w�W�,�l�`��h[;�6�ա��3��+�$$��Uո\j�v��d�ғ�-�1`�{00b0����#c�n(�7������3w�sN�53ٌh@+X�RZ�ޜ��F�e���D�W�4����Oԝ-�IA�C�Sf��+;bΖhc{vq�np��l�0�"�]J�c�jѓM�Ì�܊���\����m�Nŏ������|̨�~l Lz\2E`*�����2b����+s��2��T���k���?��$���i-��Հ�Q��m�M�L�^>!Ř��9��,tj;n��L�<��tĤ���l�!�H�-jz�\�p�_h���6($h+΃U�)�=S�7Ө���F�9Xjϡ�;�莭��)��u���i]��.��d�n,3B�l�LlLr5p�S*�uk���S�J�:����
V	�F�ա�m�����F�Ɍ�͍�ܭ�fehk�c�2Tg�&>���:LR}�܂L�M��������Gcf0&�����)��F�eˈ���58�i:
���X���m�~
v��l,L1Y6���0q�1�|C@,�2��㋓��l`j7D7�t3����xP&g��ޯޘ=I.�,*b������~a����?q��_j���c��[�~���j�)��sk ;FV����s�8"zD{@�}v�A.-o�Z1X �8��0ڞ"&#�>��mb�������h͙�S�N���b�(�������4�%X&3�/F��<�)C�?|�׽�N�!���qaY8b��1��:�L�(��j�9�=y/�(�vͽC����'!��ɂe�5c��G�F��pԞ���:�����bӏ�6
&6�e������&2oپN�����)b�]SS���0v:�T��f�e{��$�k�^��e,d!4/og��&��Y"f1�� ���h�m�w8����q"+{F2#�RJB��I)#�LF�dKd4U��ddd*�gɖ��=�������}__����8���|�}���V.1�<x��W�V4mޫ@���*1��s�o���e=ĺ�"���j�G��r�Q��i��L���Sn73��	�K~��A寄�
:�}�OM���F�,5�J�J�\0S�s`������L�Z����Z�ћo��h#�
�����p����YgVu�ǘ��	�tv�T�?��/F��@L���k�#>�-�2n��a����9�#�@0���!�t�MA���-#�j��X����Q9��w?r���o{��<�/X$X?Xj}�����%��Q7/��󫾄��C���:����
b{�ހqa�Π�����C���-7.Z�e��8�혭|:p�"%�V��)�2}�51L�w;h�p��gR�÷~4��&X	XX��t8���T����D�i����~k���p�6�4.w<��fc���
)�V����6��>�����z�`�``�`�w���Ҍ��9Wu�N�������离�\�.ؐɜ�9j�`�`-`�`�`�`�]���[�����b�*�|jn{3�	�f��p��/RfGe'W������v_5L_quy#�vLc������S�EI�֐o���/g*4��yu��k��̼Ԑ' �~}cJ�I�}��=���Ն�dů��?�H�������郅����X���@�n��Cq�G�ҥu������v�o3�Ģ�\�fq��1��9ke�{*��n]���DC�ix;)�3���i�K�t=��H���m�K���->�����k�v,��
����&�+��f'A�ܵ�,���/`�`\`3�}C�Q�Z'֊6K_u��0�mKvN��Jp�+c�`����v����-�(��ż
eG��r�� )y�N�V�W���Ub� j``�`t`��$DZ=֛��R��(??�^7��5aO�x�R���$�������7�~d	jj�|m6����)bi`�`"��[�&ʻ:������eq'��}y&}�*�NQ����@��A�X�e��e}8��w���RfI#a���Jgu�?X)X�!�uL��Z� a�_3�;���2L$YO2cH��Q�#���fG��#J�	�x���+9�)�/EM� ��`GW���0����?�Ǹ3��c�z��r@�H㙭����]��(0&�\������3�w6������f(䚗-��6�D1/0O0g0L�����A{pE뛐rǄ#�GD�a���M}U*	�(������iaP��O�Y߸o<CZ�1����>j�8��D��6��-����p]XΜ��ǩ̽���m����3�`U`3``��uM"�����/�v��Y0W_�)b}�zMj�6�]F�|��y,__�3�_��m��Unٙ����d/]jy!��͗��]�0�ѝ`���8{���b���ݼJ��899�)�i�I���邱�GG�3y�
�?�/&)�$6�]���~�"f�	��C޻c�1C��?-ҸoaI~���Yc'�I�'�d`�b���$���V�Vƛ����������T^eԮP������ʛ�%�1��?X#����|�:�J����������F�E�0v0B03L�,#��ќҾu�.@�7�h!�9�aV.b?��l� Zl�װ�F��N�3�eTo.�s��+lL��N��J�2���T&���+�� je��Y_�=��M��C,�!:L\6V���l��9���6fo�҇�Or:s��L+I�)�+�7�f!�Q���=��M�#�%��VkTy��w}�>f_���w���������ډ:n�5C��M�S�P�LN~�Bۘ�I��Y�X�2�_�e�`��w�R�%�e���y��n�K�|�V
��.�XX9X�v�e
ֈ;������g���_O�Vq�	�΂�V���ųUN��}x;F��EVl~3C[�؟��%da\kn�w�H���}�I��뾂}�{�ss���F��wv��s��^͆*f��X�ʨ{���'�+Wy��,��ȫB]�����v���)��
X����D�B͈�D�<������|�ތ�k(�:�N/!K�f��˿e-��V91�u���E���E���`�`V`����va:{Ԙ���ꩣ��{��"�팾����0�
��R����mfe��5{~�qÅ�>v�t_k�6�j������	��ux�����н�ۑ��,��4�ڹ�Y��d�W�x���%X(��4��`S�n��jq�vi��t޽�V:�f"��+�+ ����_aHęܮ�K$/�'��^f
����-��X��k����mݲ ���/�kj]r4eqM����N�yI@����`L5\W��<�-�U������]��^|��}�	�L�5������6��xus;F^��h�x8s�a��6;�����-<2�Z��9&w��r|�Ҽ��SϛQS�c�fԞuW�\n�tԚ�`S�-8�}7�Ol*��4F� �*�D�7 ��&�,�?�6�US�3�$:=Q��8��{2���{0r2��Qc+�d��f���H��V-h�\�{#�Gfo�X3��h��������=Tb{E^E$7�llb]����
��O3��婔C��d-�\�5���;�Z	�,��)�90�O��k�����?,F~�%S�6Ԏj"�Z���F�,��>��k�B�T�.��g6W���qKt����ptU�i�<���������y�[T11��U���<���ZQ{���u�5�ݶn����SrW��l��d�iswg���j�Y������	&��Ob`b7�6:�=�A<��`�2���zXW�޳��̵�Q"e���4`�b���n�t凍�J���N#�JWt��Q�� tw��`�����T���)����{���w�ȁ� ���#�#����V��r��(�a��,@6v,� 1j�a�`A��p���?�������W�9�\C1���	��)y�^/�7�7�����1N�6��9Hӹ�y|��x��ⶌc��1�Ƀ1�كe�a��/�a�,��I;�DA�] 66���b}``�`���� "�{~'ͤ��֩�ډ�jb`~`������-U�aO���������O��sɦ����D����[���̣'oZ��c��C�c�Zs�K��D;��0�9X(�kLw 5g�G�/si6��*IRM�e�wk�!0cԒ�I�L�E5b�NU޻�������GÚ�_v��)����ԉ�d��j����F*��
��5����:?���������8J���2�5�XX��+?�����8u�5��A��&!�^���	���Qc:��0���̯aq��c�󩹒���̢l|;�?�M�k��5@���(�'8[�;Ya��a�tN���!�ɸ"`WRY2��I:c���h�C�ܸC}c�Y�[>~�W}!���g��d�Z�VP��D�lL
�Q��޳�9�/5|<Wj�n�M`�դ��	f�\T]��Q��6��x��?_��*�����W|�P�4��t��A�m �ć�ļH�3ELu��m�3K3�����g��G%�Z��=\0����'�%G�N�F�|[��6ˁ��u����� 2>n։�#s�`�`����Y��]���#0��#��!�کiW�3v��Df�c������=# ��	�����ܭ���k'�_ΖmwUw�v�	b�Q� ��t`-Ǜĩ#ӄ���C+gH/�et͟@��N�Ѕ��K��s�!Y����D�{������?1���w
o�sKLC���b�� j����Bk8�V]��~��gLK��[��^�`��B�G�=�D�����ׂ�;����*��F��*B�ٕ ��X��v^WM9�xޚ&���~r�L�;�7�P2��O��-�tX��~����p��rZ��So;޽P~5��D[Ƴ00s�A0^�60�sۻ��bV����) }7��A7XXX�5b=`�`����Xc��"?����w- �G%�����q�d��=�ݹ�x!�kC8�+b��%��@���]��5�Zޛ�~e1F`�E0�5\�f�F�m��0��#*�9M���x��5w��Q���woW�~�z���ر��ӁpQ�\kK{�1\w,/8�l�5�ݹ����umx�x�����8����:0����x�*��v�3z�24����]�X$�?�.�_L��Z�W�� �~��f���$7E�)z�fP�|Pq�o���@�5Xfy���~QJK�ڀ�i�>j��N�!�����V�6�/Gi��n�#�w�9�K��[���l�*�
Ɔ�
�2�2��_�$���.��dj0���w������ZW��B�
��X=�Ù�ºR�����\w�?zic�r���0�`C`�k�K�d�!��F�3?v� �{��^�Ҷ�Wr"Jk�}��Хf�ew1փ�'X��ӎٛzA{7t�?�b1�I�v�7�3jE��CW�#�q�;)ƪi�CsgO�Y�m�1�X	� �:���&;����ʞ�%;��w��y8��/C�f��t�L�;���u�"\��c�����eG���$3k:�Հ��������gU%�D6;i=�Ub�6�9Ԃ�^FL�$�YYI1�6+��e�Lܭ�4[:y�S�U�<t`�`_��
�Q�A��7y"�)�걭��'A�L��پ���g
���1����yԨ���d�����hO;�H���"��B�+=]ݙ�WӃP~��X(�	�C��%X�y9q%�gL�IJ�'�<��mCl�0�4ư�I��R�Iᄊޝ�y�����N�vZM�%G�vu����`l5B�1
!�?J$>��z���l�LL�	5�(�4�赊����o��XS�>|�����6�G�LLg���"߮3^���$^��e���.���8�[�:�#nP��Y���nK�:`@�����L�K��j`�`�`6`�`{�~��n��{�wf�Y�K����28ƺ"
F�)11��2�|?b-�a��Ԙ�F��p��X}���c����A�୴F{Ζ��N'��j��/8H�[�9��On��ϙp:�h0F��k�S;��#h)_���s�9�$����,#�>�:�:��C�����(>wt~�Y�V|��4��A��RG�+X5X$����c|zZ�ڝF��.�+M'6�xO�W�4�q��>��	��wo��f�ӆ�,�r�~�5��M�yS�K�0i0;��`͘�j��`4tr�{ߑ�K%0s/�Oް~H��ڣ��I�m&��3X�3��|�~���Y�<:n1��d&����=�yWǭg�`"��B�����p&����3��mS?�ו�[|�l�]��v��FvL����#��S�)���\��Ĉn�a�be�RP;����
�ř�|�^a7פ���4	G-���nal��`�=.�@pi��f��̜��;Z~�~s�K��	l�H����-�Ƙ(j���<m�����+�>�I\��S|ZW����>��M�ˎX.����Ҫ�'�r3���w�xb�͚��<�h5Z?�!_�_;H��HW���ܨ��@ˀ;QKEԾ�N��V�	Q�a��:0Q*��{��4��J�Ǆ]PJ�wuA����G0�����_�k�T������S��IϦ$�f��@-bH�k~��n�q)c��򵦵�T�%�uB�f�������~�,��s�b��R5���*u_�n.�s���阹?E5�EWb�=\�81v5��A0=0~�}`�*o�p�Ҍ��2�<�[6n�g�Ama10i�G`Әg܃c���|��dWx����-w�!V&�c�n�P�qU�$K��t�3��K��zkVe_�D������˽-c��$j,ϣm�]xv���W�ڍwi�F���F�����Cm��`)������4�66�_e�7_��/Fqާ�o�%� & V &��}��Qd%�ז�Q���|��p�[�$+ُ��~�����1�E�zF>�����({�fJ���������[y�u�n�#�*����㉏��u�}K8�X�}Yhk֜��ɣ_4|"-�hz���p��=c���_����ޮ8�n'�<��m��Y���L�ʻ����ԅ�lc����͂��9��Xl���5�F�e˳���ْ#����by`�``��N��@���+����Q?�%Ɯ��Q &vLc��̉�=*Ё�ϕ�3/$qޫ8����)/���q��3�<�QCGp��	alg��?�I2��vɀ�����۩���]��f���Ps�Y�t�}��#r<�Ռ�����!��`g�$�lշY�b\`'g���L��?U"|� ���|p��X;�ºw�d*U޺L*�����:[|gF����i�����_'ט��-Zj��6 �
f�f�����i�f]Q.�Q�(S?n��ZT�8b�`�`W�Nc�I��6kQ5�]q�T��8�`�M��@E�� �0�������C�y8p����(���O��6)k���2X��s����z�'cĨ�:7�6#Z�K�Y姤��?x/��f
vl,5�W�m�E�у�fi4�~vB���f�XW��@�m���u010Í����������"���T%fQ�:�y�Red��1�YL'oT&)7��XS��Q�ծ��ΰ{�μ�C���2��t8S0��ܙ��/e�D������90�H�d�b��N�J+l����5��XnH$��{��WP�&��G����ؐ<��}x��x���uM�o��-/���N�>[�|���`>������	&��X�eUsl�۽�=��t��ѱb�ިE�C,
�,���@H4�b����;N�~���iARK1��R8�Lݒ��'�5l���b�!��:���U�6_��v��<JYדғA�wWKH�,�Y�	��Dm�I�N�������h��g]־��1�ف��;���1bZ8Tbr��y�w��~�w�,`E�Onl3�qĢ�R�8q�3}�j��!�&��3���7r��X-��,k>Ý����9��/���&XG��Y	�u��"v��&&
�,k{�`&�!N���bZ>��¶��<��'�O2bK`n`-�e�XS,�<s���7�TV����6�#�c=t��e��#/��]����:O����6ܟN�(�^���2!�]C� �X���2�D�+��'�~�����m������*�]�`��<��%�ɖ�=���oVQkA�X3���|�Ʈ'��Ee���b���.���)����Y4�Z1t;���l cJ�A�����:JN�zu��k�Ł�������`�{�Q�{��������ˣΥ�k���F�g��@�6�,EL�t�������m��,�׉}t;�[�%��k�r���n��������[�c|�O�ԓ[��g��kq��c�"X(j�`��������у��;B�o��-7�H�Z��	���!��ւ����z
̵�,!^F�t�$�d�ds�`rX�c9�j0J���ك)�]��[�K��3�P��Fo�>���2[�Ȩ��
���[���-K�X6j�`��*��|k�J��2L�@������`U`G���^��e�-j�`��*��
)�dD�Ї*_��@K��b;�XH�mB��߿���k����c���G8��Z���D���W���ŢE]�n�tL��gV����4?Q���0�_)�[2X�C�O`�`c�ѽ�Yr����yJ3�_cxM.��v䀽�A���i��Y1t�C���c�DΒk�O�f������L,씬�ygh[/޲&<���Ơ��/<�Xq����}5���C�C��Mʊ1��Z�Q�V�u�"�?`�]>Ԭ�Ϲi�˯�J���&.5+j�4����nb�L��"����7���qߎv�[�R|�	�	�^�~�a��]/���.����\͡:�S��ѹ��ڱ�/������۩a��0֋��#u�l�l�������<�����V������P|���\ѵ�Ճ��\h�>|�_�le�"�����}��"�F������`�=ֲ,���4˗֛�������t��q�R�W9����m�Ԛ��w���{���~Uc�,���n��; &vm{g�L�Gߩ�����m���ؼ�$�"��3ĦQ�TK�����������Qf[�k.އg�1�F�f[��(����v���0x�*���_W�mE��Q���u���=英��:J� 060j5��[{&=�^�>u���R� &��Z�*b'�6��u��]�	پ����!a�Vn� j� ��c�t~��C��bV�IW�c8����yr4�Wc�Mi�7V訿�#�^��^p�}Sܹ�:�K�{���R5 ��� ����F�&��B�mN(�)ΓL3�m�1AF��yn�m����`$U7N��ks�y4��ݻ� 6�d����#�ɭ��_6b���ߎ��������7�5��v�����L���LL���5����%q��I`]����@��K`�`�g��/p6�ʩ��ʮ��ݰQ� �1���/�!�z�)b�;��M�h���lqzR�o�f�Jr{V��[���������Y��y�r��/�p�0m���Խ�bv�	_$���V	���/4���=; ֛Qq`��Ѭ�����r��o�l�f��b�͍fK�<�\��ژ��[��B��,9��&��vq��6i�[M�1/�g[|.�c���_�3���Y���M]��<����jC0M0q0Y�0���p�5��:EQ�(k�{���`v�FM�6��6����*9eh��|Ҍ��t�I���
�^`mO��GgU�&�M
?�
|_�Jn������R��QRv���H?5���t���!���9F����� �	�
�<����5����C�&�7��;���Q�G�!��
�ÙA>�*y�yR�iq;�B?O�j�Ĉ��O�\�*���a���������
	��#X6�6e2�_p�2tn�ư��ɗ��ܹ�1���=������H��st��]M1#�z�Y0z010b��ј#��͟!貌V⮗t�S�xMG��l�pL+�b�]�ALLLgOZ~Z.�^ۖ�w�z���	W>�˥�xs1�wU���:k��GM���a̒���p}�5�]��`�`��<�������	l�O��=p꽰���#���0��Qk�Q�=�^kOX�&W��R�2����Hw�L�����6�p��nnBb��p�g6`IO|��xr�H[id2%
�~�:�D��+�ݐ��Q��Ks�#}��ǎe�;fV��n��{dpb����:��������;sj�����\<#�]�vnVN��]
1b�t0m��90�V���bE�T�Uo(M3����H��Ե.�%ݜ����1����
c��٪��#&vw��x0��f�r��	l�
�ӭ��� �0�-)�0͓WxG�������;vL��L=e���G���}�x�_�;�-��.��w�,��Q�M�q�k�]���$رʐ_�D
�t8����U�=��.�����AK:0y����T����$����d�f��_LH���Ry�{�M���"V66��p��:x~	g�FWN���U�}����}e�a01�Ub:�k�n�3nYYo�>�����}j2z�`�9��+�,l��JP� ��n���(|��)"$�D�{�P�[�"�F�T0^��K�K�P!��ck��r�dX�F|�g���m���X0�H��$�>��]o��Ӄ1�C\�lP��I��7����U���ϟ�2[�}�rK*Y^뺗�b�}-跢���<�)X+�t�qfxSe����>M�T!S��۞d�l�b�P{p���mv ��V������/�GS\:$�{̨f/�I�0r�Ò���KX���%#���K[�䎐�������S�h��L��iԨ����5�̓����.���h����?֏��qB![T�VB�deB%;+�d�2K�(e�M��2BI��"3$�ޟ�r��=�s�_���xj�t7yk4n�vT՞V����!�Y���
����C�㙄��x+Gދ����/���)�Qv	�,�0;5�ʇf��b�5����t��xO�:�͎�c~Y_���c�0,mbXk�V7#��h�0Mp�%�D�b���]��cSD:ʘ�.ʋ���rH7a?���F��A
F\B�{r�e��������z��d��3��o�$�ZiHE���1����R���V��m%zUqR3�Ϟ�/p��z�ܞ�
��� ����S�>���M^P\��k��i�
L��	e�h��dŴI�9��N�(���XJ���f������57�|����NR�a��O�3���	+}�]��`���Lôцt`�`&`-��-Z�W��BY�?��L�$�P&���v�k�x+9����|�Zh�V׭�:���5�4���d0�O� $�*#�4�� +~;���8�m�r<�<7���Fk�?��a�q=��a���d��m�)�u2�0��=�[ �{���-�<ؓ1�pW%��(U��3���Ɠ�@�c�=�F!���E��#=U����$��h�p����DD�4H�$kv���w#���������������/0��_��6�^�!�B�h06���N�ȉ��Gż8�����O���U��L�l �C��}u��N|V����T�
�O�Ɲ��0���a�F�����׫�XA�)�k���s����Z�n��s�{Fj�cM�6��#�{JG8�q�#�������.���`R`�`�`=h�M@YXX�4�d���d�nG��>3A+�}D޻��e�`|`a&�H��3-�r�a�Xx��S�+�zh[h�t,,�Kg��L��I���"f�O9�����t����KI�.Vl����[�Y�X�:��j0��"O�����T`��QvL�|�fa�.��.[�Zk��ޠ�pk�����5�y�0��gX���UO�p�KQu�:堡8�J�@�v�H�SJ��1Ɗ�X��`&`�`l`�`
,G�^��M�f��l��@۲ʶ�����M����+�(�����_F	��2Y�����`"`#���jV>��(�gRd-ƾ��w,����H�s���m߀X�8�@�D�������̩J]/ş/��ł�#C:5�9��L�m��>[�,�4�|ɷ�C�s�D�`���Y����e`3`��P7qr�|z�,����������aX���;�v���K�:+�����M��6�ӣu����L��MGE�R�|�s���H�g-���l��i�&���.��+��b����c'�7p��%�V�����A�dR�WR���5�W>&�m�*��{R���N�w癧���T|L���~��t�G9�� ٩}������Z�,�*s���L�<��^?�2$��ʥr�aސ��\��мΥ|-�n�7�7_�s�L�#��2[��)��J�[�O�٠�>GĠє�^�b��,�ajPIx�l�tJyQ�GZ���&�Ǿ����x�'�b۪�P~xP��{���G�?���4�L0ſ+���$h���.�׃APh���b���>�j
=~`Σ���cѼE���_�>6�U��G�f)[0��(���f�eo��ΰѩ�x�i|�2�:�:��Ϊ]��6I�@!.���GK�48E�f6z<w����y��N>~�ˊ�P��D o۹�q�3�X�
K��e���h�ɓ�ν?v�93m� ϕ滝jO��<WhЗZ�H$�����'铊m��xy"�*�v
�h'��S/�M[}S�J�u^+m��L���#
�&&��Io�=�y��3O��@P���+�\?�tжf�a����x6R���?��2����"4M}FU	V�%���'`g1:�4��g݈��5n��X`���fF�65� �S���=q��<5/n|9��� #��A���ݬ�kʈ-�Q�y��bt��N,����ҷ1�ɱ-�D3�T��3�`n`"�
���;�
,aǴ,α��mΥP�I�ӚL3J|�llS�bv`ܨn,	ll_�@	��'��Ή���C��=�1L,�j�J�.�C�T�K�yq��+�w]�n,_����QFl�	,� ,�&��r��&kn��8��lĺ�I�`N``�����l�+6�;�Ab��
��}�`�k��&]�s`I`gr������X�6�Q&��d���s���z�<)��^������mK���e�����~Ċ�V���p���gC��p*��µ�Y�c+����BY��9 vF�!F���n��M"=���[��d��"bF��� ���5=r;�g�M���1�b1c��b�`�`-`R%(�E��Sm��B�h������+�o�t�2hk�g�v�o�1
�U0l���έ��r<�%���WN����r0�I��D��̓����> 7�L'����ʣ��1�m@�فK`�I8��	�&�������R�ɀEk�s7eB�>��^��D[X;�ـ} ө|�܍��h��X�9�����1��S������[���8��!0�p��u7I��;jkŚ��5��qb�;0=�v�H�-L[�7`.�N����!��9g_5�Nv ����CU��՗���`v`J��]^�rV�A�\����,+�w���m`�`�b����V��绿�1:�����v�s�8b�`�]ml�``]`�`��h�~�p�3��M��G���U3����Vv	�*FW��r��[���i��✦��h�O��:gAV��pI)L�����{MWz��4�s���K�}G�����T�.c�=��Ʋc�M�'�&�#|%X�4�4���������|�]���t�3]�.����a�i��^B����[�D�A��>�~���0ë���Ri-����R������w��IK��,_��	�Jy��&'�]0L����1��u���H���1�bG7;��	�՗�\_~���q�-�	�i�1�9"�R�:(��r�VzbB2.�M�m,0�Bל��Z�;v��ц�tk$�ߖH>��M�[��L%?�	F	&6��.���m��H�v�����[�	�W�+��Ҵ�3�[��X:Q�M9��`�݉v-6�Hi��~0e��6�6�����&Du�J�H���n��������7��h�AwK`g��"[��f#�	����O����n_�\°&�sh�yt�q��[������g��Y��� �����.�D�f������A��i�����qr���O�z��������݆t.��qyϴ%�=���P�?��������,��|U��0υ?�O��^y�<�H��4�� ������K`�`1`��t�.(n �F$z�R��ǚ��fVe0���Wyl��lV��t�K��ܼ8�B̺����
�SX'�+ ���\s��֑-��k��*l����R��g��,y�I�����-ݹ�2�A�ST��O�f���}�>��0C��J{ga/�N���������C�5|_�jέz�,�mq0ۆ?v�̺��1[�5<2�؁L����GU�;F�6v10.�`�0�EY�>�����Ѩ��K�[/J<@�6m�$�5�B�I���S��i_�<=�o������7[��#����Q9X��'�_��B�T&�����I9�&XX��Fҵ���tE�3Ԗe<׌Kb��>}=_&&&k���o��;��2X/X�~�ׂ��Q|ƽ���9�r�:*�6_��`k`��mz;f�6I�Kx�g��d^��F��C�x�Ю%��;Q�Y�	�u-I�y��#�EY������Y!��}�ͯgM�r�Y�́Y]]�E�8�]���6:�R�W$1Ӽ.m���~磺o�:v�,�}cc���{� ��O��T�����<�~�P�^�bJ�;�M�gl�C��=A�tG���t�`}�C�F��}r$��/�虩E�2T� vl�l�erh�[D���>��a�O��u�٥"�$�v��d�}J�	BL�?�>�=�F�{O	>m'��ܜ#�w��8L�� ���[ʪ�vlm�-�'�FV^��۹�2¼MǬ�h�䗋��U�*�s`�`�`��!��+���4�d�ET�:»��.�f�2�����"X1XL�h� �ѷ��
Q�Z.�s���&��KT#V6f��S��N�5":~��N��k���^m�q��M�m����D���Z�#d_����5���Y�󑕧��}���	�v
�;F�A����lx��Y.=mj<���Ǒ��^�s`#h[����1�Srђfh�z�h��[��q�3`�``t�6���9렺C`s`y`.ʑ�O�ۙ>�_�/w�Aˍ��ك��9�}��0��m�������꒻w�$5/KO�v��b��⥦?T�]���%���T����쨖�>�A��ЖV���L�|�Ew�6_/cg��0U;:yy��6]�-�.�l<l��'0)�x�i0�P�)���$�[4i�u�n �6ѐ��L`�Wg;�6!t7+�]�t4`�آ�~�Du�7�
�m';����,� ������:�M�M"6�E�_�\�)��
��.�LP�.x|�1��R��5�Ձm�Pq�0����ŉ�Rx�J�~�=#�ر�Q��Lm��헇�u�E�-	=�_�z2�D���5�%ڶ� &^]6�X�$�X���]���8џ�Ѫ:���[V�
&��Ǌ���x1��'�)�������?��-�?�l�R���b�x��k��3��x�B��B��>M��n������lC��o��
f	V�am``�)����x�%�X���.�v����s�q��ú>b�`&`��1��dT� �/�a�閐p�TY��g��61`1`�1,,�/-�/�&� �
^v�"�n�~��8+0�)�:� Y�b~`㞨��	�4��@�q�9�o4���R�8~�{`�q0e0�ߒ���`�'����T��eI�'�#��[=�{,Zb�1|�/�p������L��U��I�����H���{0�1��(ع��w��H1�;�[��x�+C(�il6�E�A�I1��fml�F�f�c��a�(�LU8��sE���Hz�E��`e�yD�ecX*�S��{�*�<�2G�{tv鴷7�+��3���Z�9�كm�������u0��^��}�k��|;�U�tC�KfX�-��փ�dx��X;�
X��)��T�ʖ�sdY�g�M���F�;���,��։l�;?����>��>�oouq���Q�/"�Qُ�"X4���NW�'�{����R��*���GmO� c��c�`�`�1���/AG��K���e8_w���{#�2>؛�PĂ��Q�)bt���7�-�|��Y"`=dVa��qä�`����P�~T��y0��/P���K����.���!�C`z`}]�wT���d[nJ�s��A?cg���u`>`�V�f]���Ŏ�v|m a���2lR M^���� �!J������
������ZW+Bwq�
��H����7�0,���b��tѼ�lW����V��c`���_
�U̦F�
�]���@�>�`|`~<h;/��r��M���m�Yjŧ��S`�``��`�օ�K��Y}-'C�'�ٰ;���ni�,L_��
L�
l,��C��d��j������C�\CmU��6���ӝGf��{Ϯ����[�a"#�q�#���&q(��
� vL�"�C��;���:�$���!��x��0�]&6=z�1i�d0'�C�3X����#^������'��(#�+��F�a��-�E*Zվ�z�~霩"ٌճ�0���s��n$!�V �F��u*�1f2�&K[�vO���gA�,X&�%؍]6C��ݓ�:&���jr'��12�>�!����L���X9X7�M�ѝ;ҭ��Z�3<�s�R-�s�G ��s��Z�E�-��9��0���W/���`5
^��4�p�F,LL,�pt���R������mm�V�o|L�9�FY[�:��6�e���m�_����@����������0��W���`�`F`�!���Au�`������eH8��l��|�.6�iΚ�T��eL����L�F���6���������z�O�׷�ƅ�&���I�����[`�i�̉�<O�q?B��K��3
0��h;����nC��>B�`
y:�j�AI9u�iֶ�̬���Z�䝴j�
�,+g?z�/����oHZV�Sh�DoTB"�{��ȩ(�E<�J��2�u\pX)�{��:�/��u��+�N�K�sz��Y�a����5˟������f˨�K��W9�vx�v�'�,$�P�Pn?�V9��;}��l�
.��6�ѵ0jB��jnv��_Ι*�[�[sL����g��1�\}�Y�Y��c�S[�Wq�8y5�V;���)���[0�OQ�0c��49lܒY4��{��#s����68�5�!M�}gjG7��D�����4h�S#6����������J:�\,_��=ng�y�m�et�[��,��0�$�/�W�I�7�f���V��`
���~������3mMۄx�M����P�*�`u�#A���86k�7�Cm����(m��Ӛ([��&}dm��R��{*[W��ʥP]�c�墅�`���t�ʦ��K1ԗL�3~�TܽN�'.r턡MvTv���P�k0����P��%�����!��9"��$�����i`�`v�f�;��-_N5��{�8�Ц�񧛱�W��b��!�A����;=�����+������v��Q.�L�IbV�çkI�r���0\�� kԼ����*�l�m�`u`���er���|U�}N�B�2�~_k����س��)P���i�Ǐ,�-w���V�[���ʴ�[s]����S��ax��o��yi�����G��&�N�����ց�%���Ƕ����ȩ��9S0�N�ۋ�~!����2l�Oz���߅.�?�}ehS�����k�Ōˮa!p��ӝ�����4���`T`w�� v�ړi>���_q�|����q�<M/�A��u��3iq8�����������Ƹ'A�2����R�Bܟ:��|Ո7����L��/6������|���Xh��U���4<1��i���ߍ�hH�+���<����q�(�E<���/��mX)Ůi��_�G<1�TB�Ȋ���6;�&e�~[����Ƒ����h˻&|�헐�W%���|0�G�H��1L݁�~�]Y]�y��Tvqm�X�r������r5*><%������Nv��MS�Y��{}��Γ[w|�;�Ɂ?]�3<N� f�!n�c��ݔr�*��ې������&�P��7���.zL��^��8�k���<�e�S��A�Pi�`(9�܇Q�R������<�D9Wv ��N�L�ث́�⊅����#X�G���?�i=48��}��W��4�~�G%3��:;�N0�1� ����p7m�~�2uH˔Ȩ\]u�����O,����跣�����ޱ����v:Jad{�.���ޯ"�U�9��	�H�$z�	&���89��[�.��w�y���t�b�+�����N�<v��g�EYՄ�$���xfT�.���5�1��ʟv���Cu[��)G	��U���5OeI�?Y�sMa��I�>�<�
�������`;@ѤPQl�𳴴�@����߬�~���T㷞��c6���3>�9�;��R=�xw�[��g|�k��v��w?t槭��=_�ֽ�D`$���e�K�xk��И��P٭���{1�����o���_�ɕ�3������*�e�Y��^/8_FR���µ>ׇ_�9._������M�5�%��!]̭�h�O(k!�YYo*��^�΢n���J�e�U���-7��T��Z���jݒzK���\�/0��"�Q���%;t�z�gI|���^�"v������uI����R_?���Yc�r;���5�.gp���$�}������jzg���,����΃��=��lW�G�Tb9�ӥ�z��-�%��2��lt�K��G��qn�/F�
;�ͮܖ�?��7�W�j1[�yr��4=�$�os����\$7M4g�6�T�:u1HnU{�ҍm�wc}Q.�1����:����i
I�՝��j3[��y�����8Cf�ϯ4TKq�!��W�<�,XX��l���|-7�#{�-)]��9������󯤒=�0����c�����Y��eX�nO��Y;�?-.�����
~Wۋu����Z0-!c4;=2�2Vq.��XUK����7�d&b󳙳ͧ��s.��<�����#��xv���e/�F�9��Dy�@��!is��^�w��u,{^�mZ�"��fֽ���Z;c�*����\�È��Ũr=�;�ټ.r�b��oC������̒閚��>�fn�cy���Vp8���uU�����U��ɕ{1�4��\��/��}`j�`��hf/�]a�P��*u$`t�L�-^a~/Fy0[��]��*���{2�S2I�y{1ƨ��J��S�����G�{�wϙ�|�N5�E��3�8�}m@f/�L�a2���gM,�w�V���"��^�?�Df���|T�L���m������H��iN���.SD����DƵk5�����m?����#ў�ҽ�t���B!EG��wW�&��
j����Z($���K�6�D�ڋ-q�<$������8tK�uj/6L�@r*�kK^�5����J)ީ����~-�G�	����{�?�r��l/�i���-�Ž���"����L���ؾ�����"D�F���ł�R5����	U�᢯Ѧs��v/��Xk~�]����Ǖ������ۋ���;L�DpeX��:k]Ć���X�#����ߺ����z���%����"Ne]��t.C7���F����C{����m�mN�ԩn�K�Ck����b+�]��)�"�Mw
_��������4�L\�+�����~��z/�BK$�t(i~������7��p�b���J�)ƕԸ�i�[��L$�{��@nV�t�dل��T=3�Gj���b!1��X��+�;𜷝���-����K�O3-X,׶ZYڤ�bx3�]yz����a��mr.+����L����k.�	^;ʶ�T���(r������k�<1�_���+�!�F�;���Ig��hEq�'ؐԐ(�!A�#!ޑ��������*}毚d���s-<ڋa�g��ţ;=����[`�"��o/F��V3V�w�����5��b�F�h���u<ދÀa{t�����crL35Ƙn�����fbr���k�g?;g{�����o��v�7�w��e��D��$���Bβv��� ͭ��[�"@�ՒV� �;��!�8��3�ۉ{^bݒCU96���_b�v�/��>�����x"���y��}ƻl���A������Ҁ�e�k��լ����\���=[i@l�cl��܆�޶��d~uֻ�@l?��Zǆ~t�q)ް&�>{�K'[_�ӥWa�]���x�}���$�P�dV"ȴ�X���"@�Κi<%"���)V�v:}�Xx2rW�sC������be���k��	����[yY� ��>�f�H�An�g~;�`�-��S@̋v�<6"
�H��>I���N�@�t%%d��l�ɨ�����ٝv �Oi�E?���)݇���v���%������o��\r�2/�N�_�0Dy�U�F�ⱈ@�����b����5�ʱ�:3EK��"8�AZj�}Sk��cuQ��.�R��Ԑ��ũ���A�*�^V��Ϻ�uZڸr�n�@ ����E���M�u��`���1z�5Kވ�m��:Zt�͋�4�of��_�]�K�?�:����v��g�$� Y��7�\�X��dONza�������lG���+Wʆd�Ux̓8�jJ�?�O.��s�[���{�:4mo y�`aKv~��u߬͠U�l�ũuS��ؒ���G$ F�t�t6HNf���i�B�I���1�F��P>J�����+we���N����}h{b8�ڝ�1��������us��X�՟�*�w�p�z���2�ĈN�*�R������ka{F�o�.��^v͋���aJZ�賐�1�iFh�fľ~2�[&s�'���s?�9?��{>��+jM�_�"�n�ʞ"V`8N���^���~������t"��g����ߪ@�	Dz��hF�s����i���L���ES�-E�x����p����4�̡��Ґ:�_�*Z�-� ,ZR$%S���:=���u���Ԡ�F����2M�n��0���K%����Y�ez#��2:F\�9Bk}6?�G����9o��|�9L�.�D��uM�$�4gr��;*�C$�i��-��c�o�y#<�~/d��&����;�T�[��9�N�KF�K�|4̳�ATq�r�gB��AJ�Ks�E+<�O��Ԙ���p�/H����A��h��Y"�,Bp�.)P�z
%6�������&e6��k�"
qe
u��d5\l�$:�|�l}<��X?��w|�%�=���:^"���:"[�Y�1S�S��RB0�W�&��:z������p �di�?� �\.�?�1��G��%n���,Q��_Y�v?�׎,@@��P�y��ѫ�Q4~b'i��7 ����W�r�sX���-Rz#�7��)�2�Dt���i2	+��5S�͐x���-;i����ثj�Ǚ�A��Z�;)�߻گV���m	���{��@��uU#���cu[Ӽf��t�R��ZI��0�ZC����m����N��SJ񅸦Z�t;������X��T�s������h�����0�։��$K��I��2r%_7���VO��H2�L.KD���"��k7�e�A����~���@����� f�$]^T�P��|`u+!�j�B3D[�&'���$�]�BHU��s��T�V�)����m5�&E�M~PϫQڣ�G3��@��/��Q������pm]m۞e�P�)���Hmd�czھ�7��,ve�wޅ�ٽ��ZY��U�{�B�kc��PTn&I��V���V��P�z�W�Z�1U?:��he�������;�98{�*&N�ս�۵Tyæ�4s0���d�ۇ�1����v���[�/6t i�>s���<���|���U-p���n9�Ou��O���;���WM���7i�n�zi����5�f�JTN%OyK�tH�QU?F�h�y7��B�b�8����񆱄6�Q�_�o]L"	��Fȗ��w
���.���,��e���*X"ėٿ�z�M(�kU��c���<8�|٢7>�x���&����*�?:�xq͚~�}7�w��X�	/�Q��sr|/��Ye2NH\���tZj�q�d_�㿺�o�E��2�N����؁�=��oF���l�_-.NEl�EML�FW�ed�%2Ʈ,!
�ɄX�� k���ډ���Z7������< ybV/�7cW'�6m�y9{d�K!��M�|�N������	:3Ae�~���~���K��OЄ�i&1�(���|	E��"�O.{�� ^No���M;�F�,�k�ԁ���s�y���t��#n�ʕ7H�����Y������F������j�˙�
Q2#C���:~��C���&iHxZp��t��K��y������
�S�D�e�fw^'��޹y�Kƪ���<���M�+����7 �����g0r���,J�[w/N��p�pp'���֕=�c����.���QW#؛o�&��?�B攟�i�G�[1l@6K�dlm� �c�_�}>���pxy'҈���"�d0_�<԰��eX��4Ӽy�j�P�;s�W&x�U����\A�������B���-�Zv�l|C�8��3?U�&S,���+˸yH�Aft��n4G��|�L�Nv�2ÜT��R��0�,�����4+#�o6����;���Ջ�&���w�[�F��Sh��w��P7X޼7���4R6Z��dt��D.ˈ����ט��d���ˇω���~�,y��(rߪSkD-J\�~���9��(��T��A��;��f�`\m�T�[5h�qH� EH��6�����&���)ιQ����4�P)����_��!�/]��a#X�$T[C4���o���ͨ�C��6��qi���{g��7u���$i��I��#}��,���x��K��]7��]���O����Q�A�_�l��|�Β$L�?��+�7]0�a�}�	��q��R���ܟ���e1�g�Z��'�u��~�w��lE=�����oSr=�K��r�i[�</�'�~t^.��9�6)~Z�ʹ�������Z����E�5�8�s��B��3\�&��8���苂6�6����0b݉�Y��f��nNV�d��
Z���}�����E��nh��+z4��
.�J8�dB����m.S�L=uWG�k]��8�;�$���Qa/����@�:�G��;��?!�I����O?�3��'4�*��O�o�!(��S{�d��Hn/�3U�f����7�lY7{G�6�U2�~��ƛ	��Y�T�?�p	K,_Sjl*זs�֬��l�z��/�r*M�3�V�Qk#7��ݗ�{���^7���bbi�yݾ���2����7�jw����^/�kݧ�Z���e�2580P�?���S ���b2��D�L]>�æ5�)�.�*����>r�����{��ϕ�&s+5�ؽ���a��ec&\�}E*ݢ��L�g�;_��8˟�d���������D��9�����Ŋ i�w��-ME�5����'%U!276S�^��;��&X�3�Տ��^6�[�\3�!�;_��g�&���DS|�3c�SSԡ��76H3���8-�|�~�
�Gթ�^��'?pϽ{k{6���,�wZ�	�+�X����}FTy��5@Pʼ��M��$؂���z�c���1���~�'�Z��QA�b�j��Q�sJ�|�V����ݭNv�-���Y�U��;�Q��@<|�M�r;��x������%r�|kޕ1�
�Q�]ﮛբtY��^� '��w���V���75˹�5e��+��/��C����,�!2��l]WK1<}5o`5S<r%��5VB�$�\FZ��+�dekEe2^l��̄�v6Rs�	-�C������Řk��~�@�b����)�1�����xl��IU��B��΂#�E�Z:6ɼ�k)�.k����C�I' ��#o[�T~��	��\Ym���2�����Tq���8�nJJ��yQ�)yc�f�:\ox.:�v\����K��׸{۵�1��]71{�Q��(8�{�d�iO��w�?<a��D��g?m�6�}��H�ӧ��rwE��`���(U[d���@�u:k歚�c �P��VN�Z�o-+��
�p����Ht%w���k��UHDI'��^�-Ә�=�%i,��\ �n��(��-V}Q�='� �a3�4�fHM�0�)ۅz�	��>�m��M�ᄚ���kf�W ��G��[̤��y��	�>�}�	�}4%�]��G�.��16������<��@�h1�H��'���b��4Soj,��U��d��`,!�������e�Ϊft��Q���"�s~V�f�6�!⸩��FJ�	�m61ϭ`('Mj���a��y�X���}��mn���J�*P�Ĩ@LG�cūO�]7��z܁L�i�-�1��/b36eTj�u����PP����֪{v�
M`ј�
��'��� �\��-Z�10zpĹ��&�PUn�!]���J%�L�&46���܌�̒�*k3`y�z�E��ь��	����=�0y�?�&�S�%<J�{�9esk��h[���.���u����'sX��;Y)�ب���R�J�C��~���@��SF�~��j�:o�wP{2��|�~�e��.�([�[�5u�x 3�WE@U��\,Uy����f�[��=)]D��� �)�^SaZ��B�<��B�<��^^8��9MW��6K�	a6È������Zȗ�瑁Y����$,춚?��<rU��?NC+��b��b%Yhy8Z���P�aZ��L^f�i&�	4Z�:UAzё<�h ��ּ_�{/�{|? jj0�m��=���&���c�D��;�
R���E&nJ9��7L�-��� �b��!P`qR.8:�"��S]�@l��c� `�>i�% 9�}(&�9LzDN��÷)=�l�+KߢZb���Sj��f���v���7�!Y�y���|�>V݉"�8�)++���y�Z׻9{�	�� �ه�����a'GM�H�
��1�8��;��v�|���{���@�����fk,��K:����b 6.�T���&r�UQ����hrb�ú&���GP��m��>��G bvF\��3�r������8�bҥ���6m�6o��_��n�91�.a���91_1�)#	Y9n�h fQz�%7��XܻK�)s�w�8�E��l8 ��?�;1b�}g��k�rp��5��;v-�@I�rwD,��4��q��ߠ��S��1ι�f���wx��> �F�G��������-�e
����CO����YoR]�{����*��^ �Y\�Wʇ�3��S��D@���g�:����<o�@Q-��AUL��`�tX$�����9d�bv���i���7���;��1Hf�HY�j�!�DF����t��A����qP�*]u �OS�Fl��}�N	X����ǃ���EɁ@�{���Q�{׭a�V49&w �?�DZ��ѥb��9��≞$��?�uv[�����|�1�t�b�[�	 ]ؔ��ŁY�O�[@�]SB!�@�q]D����*�����
P�q»�d#(LU�Y�;���ǆ	""r�T��׶��KuV�bc�yj�Y�O�b߸�,�|��F!b�x��:a}���M�pL.�h6@LUT�t�^R��#����a.,�@�q�]��V��8���o������\�Xw8�+-��T�VJ|��)x�{�S�;f�8WtrF�~T��Rf��1vM^�l*�	����$���t����	0����f��2��=c=Y#g�m����N�iݜx 6�6�����Hq�Q�bT]p�Y�n�	���=A���7�	Ģ�<�$�1?е3b3?a��, bڨrRw�Tw����&�ٽUq$��~��u��b��Ð�ϵrC9(��h>�,�..7���-�uQ�Z�G^rZ�f~�5�����~e� |�S�B�5v��C����/u��wk�-�ѽ�#����\����ʽ	�A�5Wb.�H@���K�%�ۄ�y�,o��Ì�tI��6��=Ns)�bhKLr)�5h���q�*ҏ/4p?QI�(�j��Z]� k��2�9�n+��$q9*cA/jG�����ҭ���
S �L4{���jގ�&ѱ���v519�6'�r�lj�M[�h�= �H?�J�?� �SMt���z��
�}�.ֽ�K�*�؋$�H����s2q�lg�H$��l$���Ĭ�)�.s7?U��&=�p�.p� b�
g�#�r�$H��۱F��.�@�@�i;k�B.��~�N->������4t׶��|�V�9͗[�bo�$Bډ?�d�bv��s�����*+�d�%#�ɍ)��3U�N�l�xD�<bvAF�3�`Nእ��ƞ�<j?-N����_��N'�����E7�=q�����y	 ƫ�6(��Ĕo�N�o�����0��*�_L�7����K�7�ɫ�巖��=��|�a#f\��������L�+4��>#& ��N5Z����Eb��iwn�����5��<,�q����Mlt�?6��	C��Ι1c�Y���~(,�m�vRDns��L��I>�L8��j?:vV��ˋη�G�m>��V�`�@�Ec!O��n�F���zc� �#~�G��܌��W�����V#|�X���%|�؎!5��!�`��建�2~�@D�F$�GA�ճN��0��bJ)4��C�dm��Otw��M=A��fJ&�"�gmJ��>��z;�ΖꤌW3���5�by�m
_��+X"hԢՈ�ݲ�"���,Ӻ����*Q���ź��0�#Nd����
�0��Q]��������VܜO��K�����	�}{8̳ۏyi�|���+�!x_��*|�p�6���p��KG��ꕲ�^�U���p����ZgcQ�{�3D���]�����ɠ�M��X�\f��"�αbv���X{C�hu�n�yPz���E}�y�rỗf��Hn�I��"߭��c}�8X��a�0J�`��J�o�{?S���E}ep����"�q��y���#E��p���ʠ�?�*[~�<�P��t%Z�<?2鶷I9����M찐_��6�}c�p�(T%1@ׁ�$����� ��ooB��{���]��-��+�U.�q�պ����T����q�����;yJ����T|��0��E�WK�;%�w>Kǌ��-<�Ԕ�a�<h����#��������-�K!�W�
�j=�|]uT:��{e��H�'Ea�:�S�D�ZI�t��#�Q;q��ԉA����g�`���zeP2l`	7r�`�e#t�ـ�ȳ
�>\Z��֍��?���̣����N��I��Zה�`�v�44w�,Gc�=��[HU�<�R��-��jؕ�ȡ�r��sWvt/{}8b���X?����8vQ�)�+�{(�92�m���n5��o3a~:���mXG1��-mb�;A���e>c��M`��ޮ�STI#�m�5�~L�Ʌ��X~M��G�/��BE��� �T�h���u\���q���$i)�II9� ���!��T@B�A���HwJ���v��mw�����pM���v��h��=�W�2�e��D�z�\��%��8��.?�����Fg�'�6}R��{J5l��<�ǥPauE��������J6{�4�x�:�|pCQ���=�0J:EBan���h�o7z�l!K7�Y-�h{&�����s���D�d��M����D1��F5�;p�C/�����j=m^qX�5L���ZV��kG
_]a������=��۴oq���~{g�Tcc�tX�"�)�3������i:�T6I���/,�$���D:��EPA`������ғRձJ��5}�o��ТA�N޻�bf2I|	�~M2�ޫiI���-�f���
B���EϼC���{Zm�~���Vm�>#<�p���@��Z��6��z��ih��4�M�l#]htd�i�1��#ўBw�@���*J�y��k�LY���t���[Es,�x��[���=w�u��k飯�n��>�.�.I��D9��K��P�|0S Lz��Sa[��� �c�Ǽ �o]�Y>&wɦ���V��P�`-OЯZ���c�(	��t��c��h=���xN�C�j�֥�B�,�3'�4�?2�x;5��Jl
��?'���C��1��U�2GfdZ��Ok	����N�;]ѥ�1��Up)�n��j�AQ�s�Z�/�������(��&! @�����N8���4Wq[W���WL5���[(�Ls-��)[1�E�_�wc�v��DH#D�����+{����b�i�n��}�N�*ڡ����j��Q$<����޳�MQ�i@-5C#����c/E�M��W!QJ�������?1�I�鷔��$��މ��?��:9�V�M��I�&��\#�ѽ�c{f=�űh��]}<�_�߭trizj�������-EW�)����S�	�"�R�F*��lm�K��q9 P������O�j�݀n�Ӊa�}w�ov��±_�w���ð�/K9�c�u��gbyT�LQ��Fs�>to�2xA��������[Sw����!�)*�s������4�5+�� 1��!R���X�(�*6� fx���$�C44/B��hQ�j��nz�e��j��O�ټmS?@�Y��$-����^S��\z���A�d��&���(�O!؈&����p���	�C�NNTz�co��fA�oqz���j��v��x7�����K$(�UFEQ��-�:�o�i�����ͨe��F��&r1+a����tՀ�L-��"���*v'�}��������ȑ
�?�Ҕ�o5C͇�i���ɭ���'���&²��O�9�T�M3���r	cKr���ϺM�d�x<=���-H�H&��4���� f;�g��[7K(�^�e{��oZ;�����r��KU�Г&؞�ĆDx�ڡ��w���b裨��P�"�����U�����ьmwn��Jha,k��!HĐ��yx+E�&�Ǔ�'#�jT f9��q��5�`�3jG{�Z�o�k�ɏf��g�=�j����O��� �Vk�7z�B��"[ f��p��J�O�UM�[pB���u���F���<+�,Jp	Cz�Z��̇�c�����A��]τȈW�����98ĸ���S�#Q�������ܐ��q��;�_ft��=tO#>1��2�ɜh��dd�%*��V�8��0l�M��t&oPx!���ą�s�3=�2�x�|U�>�*�8�E��]Zƽ(�oxjP�'P�'p����3�f��?w��^�SS�'�2�,�nr/������5�1?d&���@�"�똢i�p.����G"V�_0��|�͐��Xip�N���[�I����7�oD��:,�/QzA�Ǎ�gɁ��D(C8���Īv��{�q)���<M'��������Ú���T��W��b� �Z�z��Ȼ��)_��9�;��,x��|6		��Ҁ���X��yU�F��R�k���LZ�� ��9��F��޴l�G��Bpb^L�N+xf#{mʲ_1w\��/A� ��ޖV� �@����:���x V�N�h>K��)Q<��n\`*�Q�X���!&��0|���*�� F.���� ↫����(;3R+b��Z��a=	g�)0�&�v<[�!�C!i@[zN�f��T�j�b>���E�ʗT�K}2��@�J0N�f��Гu����$"� 6n����i�P�S͙6�}Zdlb�3�i�)uhFD�{�/O�n�ÀS�Ui{Q[��s���8�uO�gF�-�K=��W�i��} 1�z�#���eTq��z��t��o>��P�e���O�R�����5��q�Owa�Y�WDm<SŎ-�K��U
��w@1�m�;����p���,\���#A,�b���jlS�Κ�~g)���2~���8���-{���{b�F-���ئ�ݰ)����G��A�8.�F��u��Y�s:�(}�Θ��D�j)%7X��b�B���E��Ky/�A�ms&;5����ý7��n$�/�x�5�e�2L��HE�+jթ�"�#���6R�v�JC�&��/���f�cyw~�)���b�{����5-3^���݀裏�h�z?E��8����=L$ޕvN� D�_�R�a�1e���Fݧ�\��\�	C�6 �xv����L�0{7�ֻ>c��>|��s܊H�����5��dW'6{�m��k��s�41."��bso�^I�Ym�5#C�\Q��+v�J	�t9�}���A��J���ē�6ߋy@��3�Z��$�d�<������S{"B˭o?m($c&��W�j95�5O|FH���O,�g3��+8��XM?ۂ��s��g
U;��}d�>H~:O=S��K�5���a��� �Eby�xRl���
�����i�U �w>��/w;ʯ+��rY�0L�@, �Mk���e�nEu�b)�8s�<��a#��`�K�� .���b}��7�r�[���?�9�܀ؘ1t���\������ ��M�!��qrK22�92#orTb��&Pb5�|�=�Њ5���	y���hs�G���z�,�
��xa���:~����-D裩��TI��8�埡�F�Y)Er���ʈ0�{��n����Uۀ�]������W����H��#y�_�B��U#��3��� ��|�n7����m�K���b�����h��W��6����0�@�%�:Kz�x�dr^bͼ��@�K 1ۜ���7��&Ih���'��߃�yL�Ϻ�4�.
�:��1���:6�}�k�	4&7u�3�p�d�ti����ؽE6�Ng�@�y��9*�5��訓�M������
��7��?f��b{��ҽ�b���m�u��ep�~��1�bd�J�a�g��8n���m��A(��:�Β�4ؼ�z�`�${�m��X�.��j����7�c��*�������/���Xƅ��%�ʩ�|Ϋ���n�h=��U*z��_�A'ȵ�֬ڔcb��E�ǜ\��3���.�4�X'Q�Lz���׵rÅ7b��A ���C߱��+��_aĀV�
��՚N���P�W�~�C4��� &��������&��7�D��R ���| ���̆� zM��F�4	d�����")qD�*�����@,#[�^R�;��]K��~}�+�]3��E���_+��D�$��n��7{����uF"ه�_J�A�ݖCh������.*19��r��^]�_9c�gS�X��D����?�1�"1���O��Z7ᾶ�� ���z�NMn�외�V&�'�A�A�� y���4Q͋��n�~�)�}c�����M#�"�Lat�<�:)XQ�omץ�6*�\��l@����҇+z�h8\Vͱ@fF�boXT���^
���s�\��0�i�2wL�g�κo-���bq}�{ �>��~��c-��좎�dʆ�f{[�^��)��}�q*:�G���	�(SIf�ul,�厶��`�<��	b>������͟2��GZ�s_���XD̍ߘ�+F�P��~!��4�̱�4��^�d�Z��CI
A,9�����a.��,�En�z�0�m�<p��ޛ�hql�~��=�b/R�?Y�1?��}�?��f;b�˔چgm�����)I��,$m �a�2-���G#Z��/��~�v�(C�϶��=�v�%.�LOU�X�n��A5a�_����Ӫ#?H��E�WX��Ҏ1�{N����q�C�"�b+I���1�3q�\9�v�s~+^��!�Y1��}/	�L�*�WrE��6S fZƕF=�T�>�6�ӭ���!����ݹ�ۛ!�@���i�Z�; 1���s�G�B�U��y�&��"s.G?���/���M}cZp�1�m��~�p[��Tܼj�c��8��eu_��i��Tf�{�Ξ���b���K]�f��r���z ����灍k{�_ o͕�)�I�!��|��r����af7&�RM�6bbbP��Mf��H�x���f�@���C�Mb��H�����	q`>�e��C��A��M�C�R��u���b���.N>{�^bv�\qk���%ru.ֻ�س��������fk�ٌ�sh׉�4�#̈́�u|Hy\b�+_4��vxlχ�����m�b3P=��BV�*|��LiYͣ�z�������ސE�IW��� 1g��DSz�Y���ލf�C��ӹ:�0���me�n�"����,�1��v����Z�f�na�s;�}C>_�Flܩ�a:�4�:�8Q�Q܎.:
l��B4�6m{I��%�ܙ`���L;:mV��!��*���/��;j��"p�:9�1��������Mi����5@��9i�~�P$;�R{�wgՏ��ޒ��\�EU�G+��i:d!�g��G���yd��~��N���M4dd.S���zN D�[M����g��E����|��Wm}AP75n-D<S.��:���ͺ7��$c����$�/���}�dM�;�=r'1�3��pLW"ںp}=�gX��@�WX���R�2�e~$��� b�]*�q�ȉ�Y���픲�}�@��%t�	ޞ����D���rbl �N큺{l�`����vz�/�C
b�#/V���ҿ�sE�ۖ���1|�z����|{l{գ�P3�?���1�o��4�h��A�R
nȕ�/|�/�����k+r@l�14�c5o�K����̲��Ca��t���HOjVkbd�z,r1���o�GjjM@L�&O-!J��3��)^�q� F������`5�����K�:� ���T4��¸�b')5v�1�7�GA�,&mw&�E��a��.��6�O�~�j����R	~"��-�g�m�>���8�_w���g��;�JhǗ�da>B�S1by�ay��$�"�47�::�� vـ䓺��rɫHV
�U��1$M�3+��L�'$����;� V�AO� ��d׋hOGo�{b����ÑP l[�Tih�w �$ �#"x\o�Ȁ͊��x�Ż�b���;�Y�tp~ʏM���� 9� �_��N��j�����H�Ѥ:�r�ݔzd�G���`P=���|�=�� ��3�N�z��Z�.1�jx��}���r��������Z�q:�x��Ӻ������}��i�����Qb����;�X�@�S��pڥ���6������e��$k_�	 1�`}�=HV9�OX��2�4����B`y7��q_:����롚 ��=r9�(�J�:-��T4�pB�BW"ŗ#�1&x��핰֭**���W��W�k��I�+�<�#׃ f{�0�f�"J������F�]��W�7�H�*�Ɛ�I��X�Q�nrQ��nY��PM�x�.��F�S�-�L(á�*Jbo�[�Z�����"8��4���~AtD�̪0��.}�K�}sR��k+�$�媺y6p3���<��h���g8���qd��-{EDdoQ!+{������l�[��{f��-;2�d���s_����s��{�y�����,�e��'����_��wI�[�ْ�-O�����ݡjV�3��~�����J	�6�j�����,��I�]�$n�2q�$C�y�}c�b��������	QG����X���O~�;e������;�6���b])�֣x�1�,��L��bAdM�_8��~٦���L����ʅ�b��l��d��x?Y�(�*>��T���!F��o�
��!ϡlU���5e��3�sOկ����v���~�kH�&�o���*�x�Х�"b��j��^�%�s�""W5� �_y��N��-o��-[��Z]bZ�ǝ�L���>\�����C�J�a鰕���SF�|�@�(�b�/Q�\H�����|�.^U�Gy�B�ux�j]�=����=%&�������V�nfH�o�w츼N�!�����>�)x�h��Xg� 1���g�A��B��3!L�9$�����O��>&��g�k)H�����۩.ZOX��qn�z�A����H�r���	J�"���pF���g�}�8��7y@bH(0()1��՚\��.�y۪�Ą��mU-�e��Wc�5p�P*Klbd�2��sά�pT�dH�����L/Ě�7Qۃ�BXC3)�;��;zo�C�܉�ml�)g�"Wu���af1����8>z1���8��V����GCM�251	ٸ�C��k\w0Z!6��u��� �B��,�5�*WO�!�:�0�g��!:�^U�=v���
b)ah:(B]uf�8l�g��)h*�.���h���ao���1�z�&<CFD�{d��JZ�|����n�4ֱ�G������b=(�������~ӈS��ʷn�����IE��ߟ�..��_}mqV �a��J)�++j�,���o�Db��w�=�0R�8���E���!6ܘ��ף۹]z�>�۝/TZ����͟e783���"�˹|��c �ʘ��\W}�9vw3]T�ęb�yM�fV�Ԙ��L�
k$�tՐ"�V{9�AfB�>&~ݑ�1t��~�q�,����
�q.��!&T�}$��f���mP`Z��{�h��e�?e\8�o�eo5H��O��3��-��	��L�o�IlKsdbE@la�b����nD��gd$h�o� ���Q��t��N�.�JƔ�:�&R(uof�j�+��O�̯ �iyy��X�G(j���a�~��A�$-0������M9G�=�|�'��^a�"+V Ц����=�1wn<��j�U�
�ƺ_x�w!Ǝ�u/a�鄘<E�\��ػn�K�->�[y�Ąa\��<��$ƣ&b�"՘\��ic�����|��!v�:��TP�#�x[����O��.<��/c�E��p&S�텘�՚��R����Tm	�/7�l�d
��v?�D/����x1�1F)�	�N ��u���+���1��?E�H#bx2�}S9�T�%<���ը�^�0I�ڀ�*
sv���o�YG@n�-v�w�bc�w�u��F����B�[ҍ��� V���Ŭ7���~�6��a�Iט;{(��sĤ�ƿ�͑� ��y�rbT�����^�n��S��o�Î=��ǯ������N��k�7�Y�}ܹ���̓�Ħ�:��]��R��ߙ���-C9v�ʂ��IY/��ҺC��	�Yǆ��;{�q��Q�Ĺ4߽�J�y����<ڲ�� '�NW��X5�A+��`���{sa����?cV��Sb&�}R^n��hh;��G�(1��C,n���1YWٰ {��4� ��g�6�Ln'*E��i�N�C�īs�S@�#uл��'�}k�1i���r��:� ��ƤeZ����*�)M�G�1�*��܇!&�6�옂��,u״A��@��R���O�u��gD���^��u�^�o��C,��5���r����r�J:�Ɋĸ�zUfDQ�%�)�D��&@�u������wC
�b�����!b�M��U�p�U�e��I�5π�C����t��<�Ґv�O� ����+�c���I�
�x|̚6X�؍ޭ�mq}1�X򗧺F�Nߗ ���$����O\�e]wQg����x��U�R�AU�}�j��c�U�e�$ܫ2�BX56U9�<�����b"V�C��T%Sc�qn����!1����:K��
)�X	�kb���]S�7u��
O\IUs&@l�O��~;%��|?�3�g��C�a�u0]oҺ�<g���dǆX�Ѫ/w�j9�PfN�����XT������q�Ǫ?ͪ�p>���>"{Jo*�����\�Rw�1���P,f^��`"'��AL������b5+�C"��?SA�@y��a�ʩ����w�O�!���SK(7�Y�w�ԝ��_͇ �0��Ћ���l��]7�P�[(�R�ϒ8m����O�8�
(�3 f�^�>���)G�Bc�FE���?y VM��B{�P�15z��4�b�Z>颔��r�Ig���u^g�B�Y�_�g� �o
��h��6͞%�ln���_rz� .�ت��wICL�?+�G�O�!�� -7��i(Ė\Ņ�����nw\�� ��8AlcV��!��ڦ��7�+��!�G�SAw�J���Ϝ�w\��� L�c[�]q����S:
$��.B�Z��������tW�
�- s`��9O#�VO@�*��1Ł���E�فή�s
I��0�Mസ�0Kg��4�_u2{|�Xϧ{��C��	�Ȋר���!v���ǹ��n�&H�	�-�e����NFfON,�����y�qK &s��û0&p���o�!��oq�A�1�\>�1���L}Ds�,I��_&��d��O���B�R`�9��@n����\p�올���������C&SrT	\��̫�&��_����L:&�Tks�.o^�oZ�?L`��k)�oC��K
}G�!����o>�c�X���+c��o�t�2�e����F����ҝk�4>x��ȍ����ےŤ�Xs\����6(�6f����dt`��gh��"�#��IUAI��J���}4f��"�p�i�z�k�S�� C�Z�O�Sz��`�Ӭ&�C�1��o��+�:!c��e���� |J�@6��7��m��cS&��N��*y�&�㋴egZ�剹NK�x���NKU�c~��Qs4c����/�O�eǥE�;��6;�ќ!�w'�Y���UơZ����Ķ���X��H��^Ceׇ�26r���lhֆ���3�G�!����D�h��1O�-�����K"b.-ʷ{��z��8��h��SR\!���\2��U�mS�x"_�Q����\#�!�Tz���(����l�1�iKқ�ζ25���-�ZG��r���������;�7��_H 6~2N˥,Av�&!?E���b5b���4���ɕ+��b1{Q����eV"�mʕ����i��=�p���Jmw}y,#R"��FG�!��m�!I<=�j�j���S�ͣ3�U�5XĶ��x�X��7!|�[�Cl��w��M���1��$mb.cb	��n�}�#/�ְ�ClAli�˾~y��:a����	ľrc�+qc5_ۮ6&����XDe���yr'~��oB���n�QeR�~eE%ۓy;� r!F͈���?w�/z�T��QL�A̷Q��;�n��3~:�z���N��rUs_m4�%�\P��mEA�{}����yYT�C����%«����Ks()V�l���������_ʷ�!�f$�v*<NV\��j�V^l��������$|6n�c��uLmȻ�����ۺ�E''����D�f8�-o��m�/��
9rz+�0�~<����]V�19�UoMe�J�1�O��sX�C�����TmIyM��}g�.�	b3�[s݂��v���'�7
� VOO��dH\�;���@ˣ�W�*�z��<�/����ʓvj'�3r<��˳:�H��tK!�$b{�K�ٌ?ĝ{1��,
�U�.\)���JL���Kf��Bb퉬_�	�.��[�|�t ̀X�}5����%,�*:��x� 3��|��D��JB$�{�~1̾1�Ტ�L�JT1��"�ٚi��-����1�/&ea�	��@�NJMj�\$�G��;������w�qu�q�`p��#e�g��_�a�\J���m���N�"O��JW�[�8�q$�l��)>�Y6zNc�����כ�N�K��ly��!�I��fH�%�dF���vxO�� �Y�tm��^���v�!B,U;C�̊�'[��ay'��ُ�^���:s*����H�ϑ���q�)�N$����"��[y}{��Fb(��{����v����!f�C���ᱩ�N(;�wQE�������G�")B:q�y��ˡCL\2���a���G\����߱N ��zNS����Y��M�}�����[@b���$vԿ\B�A$d�C�K)_?���Ъ�a٩�H�f:;���#�;=����������D?���q�Gj�օZR�l�y�|&�m�=3�5�2B�'R?�Z�路��;{sH�WQl�W�M[���{�?�&fәYג�?jc˯5⁘�g'��g~��+�Qʌ��DK�����j�t@'?0�Cԑ*B�Dc��g��,�>S8"0����	��*�zӦ��DA��/��
��#��3}�(�7wb:;3�a;��W����bt�yb�JQkBL�\�tNT?@��kA���y� Ą���{5�e������Zk�
��X�kAJ���rԃ����z4i�=+���=_����3��E!�[R�QL���šb����������L��
�4,v�дɝ
�w��)F�(ۨ��}(�&Fl��l�q�����̭;�q&?#P�#N�zU�!V�M�a�W��ԧ�p�5��1�]����o��ɳ�����A�6Z�m5#u7E��|�t	QiČ�
�wLd�����LT�~x�ZA1���k�d5�,����jg��<��>����2���*Omׇ�W>-Ų��o��_�&��i�b��#�?�;f�{��ڍ��"��!Vk|;h�O�%��K����Yrq�MF�&��)6� �e{f
c�b���B���;&��J]��6J�uALۺ��S�WKؑθK�N�G1��ҫ{���Urn�yx�3=����X\7��*�c���ء�4E6g���]͔c7n�3L��ÒV7D��Vy��]�%ܭ�A�H�U:�iN��K���(���x���]}�1�4㛯����\?c�ҏ�����=e��t�������a��T�����[v��x״1K'5V�b��3z�ਫ[Ӗ�w�RA�M:��^��_�[U����,;�U�ad>.)?""����W�*��Q�ub�q[���wn�x4�%�?����+�z'F'J�Zs���s�z}Q�&�J�@L��-J�_�S�`~��d�������q�K�&W0u7H?��t�c rE�Ȅ!6@��n�ˊ��Eޞ�_��a�O�� ��4mh���ePj� `Z@�.��N�nAB�E�A锔��.E:�X��K�AVJ��3�;������g�4�W�l���Ji=f��7��Ј �� �#ev�ObB��QI���� 懑5�k̲1����h���o=b���	�xm��q�^��cE{����tx��~�,�b���bS�4o�%P��;�9��0T���������Qv���M�ԯ@ץ�v4��������g��Q ��ٳ2�q��	�-�bN� ��O�N�ōXco�ޑ��U��)���=*ޯ���o=~+݈Ɠ{����Id|eA;���&�Md��&�c�؍��Ed�^j@9�IW���87ֹ���o��G-�7�K�Mw_r4JGzw�����9s�;߸7+3���Pw\��b59���S��ֿ��oRd �n���wԤ�ahLi�$c�q�:��uos�Z\��w����e��3�X���u��������Q���A�;_[�N��f���H��F0+���HZڲ��Ǌ#���9
bJ"�6���o�`�K^�'��F�X3�/�v�]�SĜ]������[�R��>1/�<�tW���%�1��΂a�RT�������w�<׼���*��g���:^���F�@,k{��yN���6Lk�Jlz���,LC�ٚ;�yk�Lݹ-��A�����+˶%z$.pgb�Ķ�\�S�*Ϫq���k
l� &���p�ͤ�H�\#R��b����޵u��xQ�&�ʁ��놻ꆜ��	�7�1>w���qI�s�A��x�V�y]���@�?�o >�?d�Bq�x,��kbbL乚1��A��!R��' ��y��X����H�S�p�7�3�[���cm⎘�YOe�$�� 1�7^!�-�i��1;�U]���C@,��f��,{w�l+szBy����r�V_�=b6*�8��c6���1�eDw��-C��yEmu�LwK2�lQ��}���2T��r1��-$mm�)��� z���' F �RF�A��*�s.�殱���q�4H���"��6��3[@�cN}���౪[����Z�|���rӋ�`���1^�!A��P�/�1Ta��zN]�I�N4:�,Q��Gbێ7���"��%��D��xb�v�ۯf�L�����3�0Rc�X]�KX�e�97R��
�eZ�v�g�t~�D�a�Y�eh�1��˫-b��.V��Ū7�u@��k]}������������qL� f����/fݡLB���h-��2��&��k��[3�X����
�
�-���xz����)�B���fCN�#�/'�T�o���;�H�������V#�커n}x��<�����dwM�������lTɁXj%�A����ā���s�A,�nkI�⦯ȨgFh+~��b���goÓ	Rt�q�T��@@�)s��H��ҿ��ډGȍ�E���2���_XU��t�O�7&�ʂ��|fl�!'�ϟ'K��u�㳀���3���BI>K���'��3r�k���-0���R+�	b�J������ ��j�&%���K �&L�T��L:��Q��g���!�c�L6j�,x\@�7�,�t@,̐�,�E\[�y�b*iQX�D�$T�b�S˻�z&9��OoL2������V�6�<���kG�j ۀĮ��=���>�TW�N1��U'Eے�g���2uj#I���(�|-~�s �4�"�6����A�+s�wո���m�׳�AL�m��ɉ1�ט�%g� :���NGy�ȴ�j�q�?b�O�A*r�i�C�rA���)]��;������5#��4�Al�A�@ˣ�u�q�z
�W��x�eS�8�b�H�~�&�T��25m�1qd�K���͵�[��wŃӼ@ls��/�^Fۡi7!OP��{�|�T� |<�Pۗ�_��pZ��]������|�J�T)�@L��.f@�`T� ���dG�&Mm%�Q���z� �.a՛b��'ݧ|�b�P�p�2a!䧍��'��+�C@l����>�e��p M��a���?�����~Y�����:r��H��쵨�lY=3v{��mR�R�9v*K�����G��Y�%*�����4"�b�XUb��j:�{�����_e��X�ظ�6��#��V%$��[R9壚8���"g�[\�z����Sw�0Ye�qqX�f,���L<2���LC�b�N���o������C��>���®z?�T���=��r�^�j�.)/��T��ҿ�|Kt�k>*ZEMN�ĄE����{�s�e����B'�A,xi�������Ԛ~ g�&[���P�~,?���˶��������;�O�i��0p�a�I��sӁ���]C��՛U�E����6<x�{��z��p����_��ʃf-�0$cU�?��؜�l���؛!�ktC:�ް��#������>��v�]6NC3O:��D|�"���Z�-z�^�w�Fh����<`I�+�a+��Ĉ��׆u���џ\3U?�nPb����Z_!�w�J�<���&~د����n_����b�W�{�F�R���������(V��ov�]��RBgQy���i �E��t��^E@������q�5�dJ�8�t
f�oE�q��4��ρ��;�f}͌�;��1޵���4O�DϬS�#��DC���u����Ö���	$���d�i׮��^�N��L+�B�[��^�s�'1b�����J��×��+�����r:����@O��Ar��s�F�D>=�
b�7��H)��^ &����G�Z@l�KvI�\�l f�;`	-^W���]a����u���E�B�Pqz�f�r���H\?4�#V��I��b/�G��ˤC50�O��q/�D��$��A���H���^�ؾ_��:�|�������3\C2� Fև��Q'��Ѡ%Z�}�M̅�BSm�))��1�Xf���>2�6Ăd�I��M�R|w&���?�bB%��;�lA��O��9�7B_�XB���fX̾�M�d�@`9Eş�x���s�pt�P�'���$(IZ/�b�hj���Fđx��P�&8��;!ɢ��E�
eSN0��)�X�p�AeNژ�Z�t{�x��J�?-���Ӎe4k��x�{�g��p�`.;,9(�4�":�n6�� 4?� �݂��ߟ�\����)n:F T�+�a�Oc�a��6���������;���̻  ��ε�K,��Htc�����i�?3����A
�615$��lS��ܧ�@����~�� \9�L�$}Qb�9"���Nn��e�v]՛��3��\��7��*���!!�n�Yg��e�W؟��|�g�kZ�۔F�L��Fv_�^e���=��y}Q\��TC7��.�ޕ��q�
FZ|*��\�t���5�0�zJ#��u��41M	i�a[�\����!�z������ɫ�����g� f7i����`u�vKImm�`Ě�N�Tux΢w/�,x�4�V��]��o�
uYN�v��Ӎ�L�2A�A�Ft�z��,�C[B=[.� ��k��,��*5�T_N�����d���ߡ���'�b�v����G��M��&�i������	�����z S�M*Ϭ�ٝ���uf{*�ibqֵ)�l3��yh��wm^7��{��E����ޙ�Mǘ|���c��\���"g�{VZv-1L�4Ąz?�<�{�+���J��L���ļ���m��=��z�$��J�����b����(9��p�04[h���_a�?l��m�H��No��x�t�����w����l��,��X��詻�ҙ �[T��kO�5�n9f�|����n�M9aN<o$�-���Ĭr*�OO�N��鴈o`8���إ�^n\��Px�_|1T�`���Hnyv�-~-����p��%ipw�ea���o��Өnߠ�Se��`D�<	f����b~�Ŀ�-s�i��C�'�D�
%ig�@l�!�>�]�U�L̞�Ţb�-�ף6���=^D��d�1��
b�e���7v��9���ۓ#�p��}�n���Rޮ���K�Bݳ�	0x�����AOK�3�b'V��:�)�T8��B<�����t���P%%f۹�i�~����4��թ�}a�����]�!�	_Ϡ��ler`=�c��n��[Ġ�������)^�l�?U�Ǫ	�ؙ�fp�s�	��ģ��?K�JE}�nВ'|�u�U�$�!>�1�1�v_�2}��i�:�P{v��-S}Q�{#U6˯O�Q���<\s�i׸8�7��E���iF�Zz������H����� �ӌ��^�Mׯ(�)`�8����u���0JR;�����J.e�`.b��x�T�)j�l1���k��Al�Rf3�tS!�a�*A����𯰫�"II=�G��C}X]�c.򛂑�Y�_�zy&����[o�ub�y��23;��~��Ǉ��~�s��A�_b51��9"z�7<����!'����A���0�4�RQ�2��s�X���7ņ�4�ivS�P���.���m�,��&l����чs�+���vv\bh�3_mj+B�V�[��� f�^\��\�~�/��6�;�ĮG�)>��#��=3-�^l���lΡ-_�o���r����<1�b��	�'�+fh��^��s�� E��Bx$+�q�4R�	���L���O����=���yb4ϡ
b�^�w����S�(�}@���RP�*%�Ir��4W�^ʄ���s.eRS���X��d�����������g����_]��R��otzr8�/�+˼��5B���u��GN/�#�I"҆K�Ŕ[Q�f-�ض1&���0��@�?�b���[��� �&�����Y�W*�l���� �@$���~�a�^f�,�I��5�ߚ����VP4��D�pGǋ��M*��i�i�Ի�zo�Y�|Ž�y�i���}e������I�HR����b�iyߚ�P�'��E�ؤ��v������pO
(��rb�z�9�{�A��A̠=���O�]4k���Sw�>���cۻ?���!�t,fq� 1��V�4u�m1�h�fFK���3�-E� s�>v_}�S��ݗ�B���z�L�/hzE����z����0�������dc��(�����V3дGZ�.r�N��E�F��N ������\���3��tp�c@,e��<q.�U/��i��St���Ĭ���Rnc�
��	tڂ��o9�����F�j�4>� &�65qG#�9�6��c]�����kh?L�wpL�>��x4-DZ��և�e�aW��&־�=���K%�ޭ��@�<��Ĉ��'���J���n���h�"��`N��B��`a��-!�c��+��Ӻ�bW��?>�ډ���*L+��@ b�<�'��d�qR\���э�@l�!u�0}��#�?�[�$����2���D_W�V�{��w��Y6��
G��?��
��i��=YAб-)�1ù�Q�ъ 1g��t�����X�(n{4��fy ���H��*���6� q�pW��M�?,�w�qw��
��c�,��j� �hB�$B���~c���<ְ;�[��ȺN1��ˎ��c>I�XT��Ha�^mڙn����'��pWWX��`v�<��|?� ��b&w��n�P���ȴ���fR	����g�h���ePh� `��EJD�4��4H�4H�%�%(݇n����!
� pwg��q�ξ�y�`5���ro�=�g
|�ԡ�F�?���1o����e��	s��^旋�� fOW�B��+}A,��p	/Jy	b�OɹiZ�~�1`byA?u�_o����A����Uƞ�ީ$���R�i3���m�@k�*Y�O�� \����'�q.QY;�B��{1��Q �f�6��T��}�k���Q�~�����$tE.����@X�;b^6ہ��k�%Co.a�w���:�� v"��_:1��"�d@�";?1�[~z�K�Zܺt��
��(�	��y��v�	G3޼*���R�C��>{A�%��－�|-)���d�	�N\���w�`E$��k(�� v��#켴�ȁY�*��k3-C�l��o�,��'�,Q�d܋"=��b���(̝ڸC��Re��C
}@�9z��h!D+�3)4��ޣ�e�)���-���m�����N([���A�ɦ��
���.��[e�r�>�Ԓ=���_E2�X�:��1��p�������k����#r���P�yWS�n�� �S�2Sc�;�V�;Zou��Σ?��CB�Ak1���B6Y�-4<Br2T�� �(�ܥ��74��R���Ё��\"�!V�������<��>�Xg0���R�%>�v�I�^_{t�I�;UQ���:ݴ��;
��w#�+G�4����M�R*�A,�Ĵ��d>��մ~%�aV"�9�9�S��r��+G�Fp�m���a�D����	�j����"��s�@�����-�C�ʳĔ���e2��y�aM��h��լt�uNl�����~�+����J3���Mq���C(�����Q<��[�Og��'
�ľ���3d&Qf�p'���t@�M��	���1�Go�s�eﲾy�qU�eʢ�2T��8�`=l� V����������R	���#�9c{
��Bx_쨯��[�gP�9�c�w؟��#�\��n�uS�Yb&�`��D���i���߂&�y|�bX�x�����q���>�:�)��m�aFa~�n��F��u,"s�A���Ŕ����A.tu�P
�.ľ�Vyv9ʝ(,U��l����b�"[�׿(��K�-��WG:c���;����%,˒��F<�qm��x�b~�k냙�"�3;[�3�{�� �"���)|J<F�sf��U%{��.����/�=���{B ��Kb�t ��
�xj�.�{���lv�I|�ngq�$� IQ���WtsW����K�@,>�p���UuE���MȲ$���6�mSb{�nf�f��S�4�����VI�_���75��fn@�@�*\MAZ	��O� ����߬�sE�k
��{�nW��v�)";u� �Tp�c��&{�"8�x�tTo�X}Gt�'/'�����n��>���^���QI��{ ��p41;��
�|��\�Һ� mC�iTGh:;X}Y�0`D�ggPfb�'�)��V�����_Pv!�J v��P��~Л�AB76���f�$�5f��{���LWH�psrh���A�՛�Hrړ�a�[�k�G 6�H�%>:�Z2�ǋc�����*���?O���A�M����ʠ �X>IM]�ﵰ#/����*�y�1a�6c����x���*�T-��ݢ��u�)oi?��8���5� �O��ҙ,��wm���� ��bBmZ[��>h��}�Nf&�:y�S�^Cb3r$������z �u
�X���\��$�pm��K	��rAl�9��d��&ƥ���)�C�W�UH�̼�%�D�L���^s� �J�����*�!4�G��i{bNT�_)sn����󦬒F�߃�����_����'��t���h �Kp�&��̍���
B��V������v��We��n�(˂�n�MEg���n��r:����$�e���xYKl���h�`��H�b��=�N��T���4��Za\�a�zW��0S��A*c鏢�� ��z�G������������b}q�%���ơ�(a�Q(� &�ՄK�I�\�� 9�2��9ľ^D���!`�Fm�f֏�؀ؑߜ�7��<�g��+�e/���yJL7l�ʺ����d<�tC�߂�����qYl����j��c��� �ɭ|/2�����a�|Ӻ�<�%E�����g���]��K��-�a?5�Iqu�ʯ��>�����`� 	b�qޮ�^����¿��x��S
�>
R�T%�N�O*1}+Xh�1����TeK�$��FD�>q��_=�	�'�,����!�M��bie��֗��HH*����<�c �m��Ŭ�'�����9��t�����g���[��P��b�~�Ѵ�����-,WY�;�U�:P�A�2�ϥ��X�R���9m�8c��Y��e5;c׏5~}cJv2��\&f�V�i͜���-�(��0���@�`��aj�% ����u8s:�4��W�adx7[�]�����UU[h�����+���X*a�u�ڬ�}���=�ЋY[۶t,z�C�9�l���l+���*�D��s�sJ�p�#���A�QP�f��<���(�������u�e����D���&��S���Ĳ��.f!M�C�D�'�'O�^����+��tyI�}�>���<P�V�=s�Z���DC"A�L��Į :�5T�!v2�1R%D3 V�C��~���N��v�)bi"��0z��1���0�n�87�%ʿ�c~�d�0� �sñ� bS��]�G�!Vp�"�77�| ��Q�_�4z{Ӣ���HMM��	�
s=�Ѭ�&L�9	i�(��`8 �2��ć�����<�ME��N ����?����@�?�T%Eѕ�Y���S�hr�}ǎ^4��!�.T�X�8��hނ#�tf>*���]y:�=��*�8}]7ػ�4�M<g�1kB����h�k���G�ű �i)�ă�^퓣���i����6�څ
�Ri��Y[h��É�X�Cv�Mi�t��]�{�L�f� ��~�F�(eb�yC�R �fbX�����:�g�`y���� V����g�ǐ�b�H��t㏯ V$L�a���c�`^OΫC�Lbp�d��#����f4���$�_�1ۺ�e��P�+{���v+d�L�b�N���
�&6��1#��ؽǳ�����o��j��^Z_���� ��%!�oi��c��-4
?κ��O0T�q�G8���Y���q�}�:->�3��tr�����Sg�GE�ӣA��P��5���� �0��rQڱ�ѵO���<�QGb�2n�I���𖅓�/�A��S��	c��ɕ�Sر������U���� _L���'��-�;��8�'�����jWg�~�ӕq�������^L�"�	dc�j��\7�is,�����9��+�,��>�e���H���X��
:���a0p����.+��*��Q֡��rl�,�	q(��=��q� ��*溭��moA�$��ek_��,��rw�sV���꣐�"��~S��مG� �o���@�kHx���ڈdwu5c b6_�.={^6��-��=yԢbQN����N�	�m8)U�P�@�VHt�kK|$5n�Z[Ԃ���P-S�Xz�����m�|��d�@��`����Y���eB����F�1�q�;��ٰy��sR��+4V�o������K�Ǩ�k�}��H�1K:c�Zt��[2x��X� g��f��(R,�|b�+�6Y]�F�#����#� &�&�$�IM�k�RKh��12~b�Dv�0���:}�38Z2)�����gOq(>��jdyɆƀ{��ӥiĬ*�ŭ�QʾmIԱ����G���1�H�P��v:̥Z-���b�ѩҚ�������̸K�X ƷtKѠd����(��K)�bifcqV�o�_P/<H��#տ�	#[7��'����J���{�� f�FFn���A.,y.3�7��8�=r�n�Q��很��P�īɮ��=:?u�zVN���`IH��اk�i�����]���/(���@�	�ٹ�v�Avw�P)j�����^�O�4�_G��FD��Z���b�b_�Ui�r�הPp�}�3k ��0�*�Tt3Wx8��}�,#xv��P��1���J|H��y�C;��ٞ
�v��#�p=�嗠p��ɾ�[������������X�����	�=�q��γnȲ�g &,'�nlI{]��_R�c��8b��[��=hI�z�?�{5:@��������M3���z�R�!�M���,p�Q�>:��?�T1�CD�U4E��}�ȩ�G�a� V}�h%�Q|nQw��\%��<��w���X+4���jH�_����"�@gUt�Z#���o+�jB��t;!���o�e�4��zi��
b�I)�%��jۉЛ�o<E�} 6 �Y0t6��3'��øTG�	b��պ�NIQ��<fVCD�5� V2���&u~m>l�e)q���4�����m�'jk��{��we0�����Xc��	�d�0`����,���ï����m�/�	ܵ]�g�:�9���#��)YG����|s�t�m��^Ek�t�Y�gߡ{�<ӽup�\�R�VH��٩^:������&��è��Եy%n�h�[��O0ﰻ��G���Ѩ]�w���H4����	�e���ZB69S�\b{�h���6����G#�j/���5�sGI��i�L�������:	������!�O[����boX)�z��&��B �Ϯ��@�<Q���I�F:���{��i��F�u�Q	�^$cTG��+���1�v��ށz�K�Jd�L^1���ϣX`���L8�8��ru�H��D��]�a���q1��kb��B�� ru��Gʅ� ��1:�����	<�-����NA,��&�77��+
�`ёg�Q���I�̩�h�����.�X#�}ϖxR;�9���ۑ' �F��6��}8��pt�vz�bϲ�mE� ]$JN�Lo�d^X�m�w��o6��1�e��-~����x��*[��A����\n�t[ˉq�-K�Y��)�_2ęB��4�iO�d��@L'�[�Â����@ ��:�����<��ߣa˴ʪ��*CrP�b��\)�IP�Ӣ�ń~"��؅���8��W^��	&N�_����m�eԋ����P�hXI��f��g>�)Z�	��M}�u������@��b{�J~�|h$" ~�B��9��� ��I~#�.`5�m��h��A���6=N!�Ƨ2$�'aɃuZ��� �m�@�>ŷj{���V��z{�J��q��N9#o ъ1����L����BI���$x�%͌�c��*�3������|�F���Z�a�'��Wq2;X�~؃X�N�#u!��"�H�L���]����g��Ub�f
ru1=1���7k�ؠ�7Auػ\9�A�t���HƦ&�̢�i kD�� ��5f�u��7�@&R�_�.���f#X@K>E0�������j�wM�Ba �(������t����y�a��3��'O��G�����Bػ�@L	���\;�+�����FԹ�O�?4k��h���ePh� P�C@B��n�ኀt��tww�tz	%���twwJIǕ��x�3�3��{o��g��;�VF��в�w�)wz5��� �ǹŗm�� ���y������?Y���f��n�q��i��դ'���c�`z�t�<��}動��숤x�)��ϒ~1[a�y]WoV�h'����4
�� �I�PK���c�d���l�O�b(�g7�m�s�xy�;y$ ����u^M��M8�ׅ2"�vz bH�ȍ�j�r������&ƍ�@r\���I�8��u�hA��+3���x���6��ڑ�v�ed�b�P͋ �r��3����?w���[=@L�nZ�:4�1ͦ#��wc����r"6l=�ãs9Ve&%��ע�`����|��+��PN����ևAL`+�k��f\&�
�75~��5�I�G��d��MM|�v��#���/��m	F�Fk��;����o�����$��X�23�o��Y�X�S��"s^l��315_�wq: &H�q�;��^.��o�����w������^�i}�=&��@�s,�\����i���v��q�b/���@l�����smE{�Kl��i�f;�Ъ�u߼4:�ʙzO^�qS����c�����>�vK;��}'-o_<����.�=0����u�@GJ�v9'�y���:�{S�b̷�Y)�?<$1��� �o���o�$v�TP��m�q�-9���ǖ�!����ԍ�^c��Ǥ-A��sw'u�@��%y��rdg3���I'~Y>��&�����U�Kn����{���Qv�r���h�SY���Q�H�*{t�_��[,�m���2/�5�Ĕ+�޵ ����`�4Øb!yl�b$�~��d����V(oS�q�~������'�;�
¶�����EE7c���?����]kIɯ�EZ�ա��Gfv�����,$@0z��U�R5���j��y��z$͕�YmE됼�D��꘩�b�CZg�k$�yaBݍ��- �`�'7�c��wK"%������uw���c+����q�=E��#/��������0����_y�L�O-ն��b��ˋ@�)���/]��l�0 �_�AW@�Q�0��Σ��/6X�Sf��@�I��$3�V�y��¡ț����6SQa�5��op3ybn��D�>�'�o��5��\c��J_+��bw-���7H/I���g�5y�k��`�?�y$��ä(u���>�rx�`����l�/�*��x�c�#�6�x��k�?V�����~3�������Ӝ4��
��G �4U��2:ri�yG�Ӌ�bޢ�c�l|D�]�p��"V�������.j�e�dx�P�A�[���6�b�f�>,ݻ\7h�lk��J��OwkۇOx�,+6��@L���s�'�ې�S}���ق�����7K������yn;	NT�W3[�l�9!I���u%!��~���'��D���,9*���>����܆ {E]�(��%V��d+��e�!'�9���RN=33�p�@��s�g�W��_V�X����x*�Ԯ��V�S���L^bJ5�њ-1�)mte�Ge�KJA�1�RyJ��P&r��}~*� b4_���C�"�ܝ�XQ�F5��AldF����@q��C;~(C�	�FF�E�/�\��[���?�9��W��'���3evsf�m.��F �H��UkM6�bU'�E�k���� �./	2BXpa�2�9����&�@�/�9eA�1>c����%��@/��)�1�ık\�_��5�5cd��I��ηt���
W���Y��$�����Dl�n���SKФ�}��cl��++���$ 1Q��̨��ȵ����a&�㥒���#	�u#9?��4U��ƃL�v:2�P���!�O��V�A�e��Z_c����ԅKE)-�u3�y��tS��ҥg3`VB�|)d���H��}s]qL��״m˭ζ�y<LAL�� U�T�L_φ�S4o��_m�/�3���׹_7ٮ|�_Av=b��Y��~�9h��]b:�?�g,Z��hALitV���I���Nw	#�Ġ�.��I���!Mּkui��~� �;��su����&�E�*��F��Sڴ {_!+��r��{|� �&�S�Qn���H��l��YbEb�#�EoLY(㔇�>C�x`���m�Q��?�,�B0xB�A��; ��{���L��0��9�+�;?Ų"�Y�Y��P�K��$���
!I�x�	$�y�܊� ��@V����蒰�d���u��-j{z�@lK�*�Di���*A�esK!XVOkUحJ2�S�'���o�ˬ3�?�+�������V4�T۟{�R��\{"}�U !K|V���՘ދ������2J�戙B�����
?�z��Qk�%ɭ����qj-P�uw��b��,9��"�f3!�(�2�H�
�3�:��K�K�N��'S���A�ؘ����$4t%�B^�9 ՟b1����h߇㤰�z�R�q+���x�Õ�s#5}��z���mۛӽv���#|�����bXOV�ӱ����/F��h;B317�[�����~��O	H/N�<A����u}Z���M��m��r��5�)��cdPD�ۮ��C�X���+�؎V'A�8M+�"�e��`�=���(�ۼ��ᐹ�yR�eӚZY*24x7Q����K��t�'�ӽ{�C�7#%T^��;��2gJ�n3�9��pe�6}l�A[*WFJA8�O�ş���y��Tb�[��utP�ι�1���-��Ƃ�,������\�6+V�sL֚(���B�^��7�[Q���96�؆�g�mUm�����nhO�O�=ʥ�����iǪ�ʵ�؊޿�b&[����6?���D,~�E�
bS�*\qD���F�4�|O|�`cpI!�1tB~�M�0tc"Ϩb�	ȶ�5�C���Q��� F�H�U��:@�j�aA�#��ŀ$��Y�j�����0hh��G�c	����ǰ���|�q.4�o�A�j�PG5�:yxa��4�~�gL��Ԝ�VH��*��=��f���A,���s���=!u*�Wu8q�e�زX�	gݕr9�����T��ف��A1*���M[�s]f F����|NG���0ć����D�;�-w�d��Y�EP[��T�G'?���h��q{F/�����@Le(k���5��I�߄���]�m�դ1!2��Bq���I<����A�Q���g��{�-Eߣ�A��Q�]��f.r;W�孕�1�����P�M[�����oA,�f�z�����K?	}(&���u��PV#"
r�d�He�i�G��X�L���<~
aF��s����6�݃�O����g��ٻ�y����u�bB�"F�E�\��b�h��F�;(O��W��C�NM�� ��M�P?�Аa�+s5$����")�M#�ލR�$�r�����a0�s�Uj�l�4�4���X�Q &w�/s1���M
�9 �_穈 �!F�&�����m�t6M�&�BM#���*�}���⎊NxT�bbi�<�Ut��5�����N@��sn�87��U�'��E�X1�o1寇�@Zܴ��S��'@�/�Bi�ZrP�B�[v���yu%�����y���UMZE^����1��8�k�5wcy�8�r���Al��V��;�zǱ���k䯸 ���pPO��Y�m�DPIA���+�i�����!z6ta��fM�XUv�!R�M|NBqCU��"LdB�}��<a�C��M,�Z �a밿��Ni؞����>`"Y�X��D��F�/-�hVr!J�\ f�x���!e$��(��%�2w��Kia�ǜ�7U:��5=慚�ظUn��S����s�u�P��:�I�-�t���̃)e~��l�9���U�F{�2���u�L
��lQ́�k��B�(�f��"F��Ҡ����׵�ݏ%<�թ���b�b;ٓ����F�f��Rm8'@l���^�a9���&]�Ҟ�2	�r��',�`I��i�o��!Y���h�������|��Y���<C�ra�O ��1��Q�9B�O�TT�7�Z�'/�͂��5��1cv�U�5-af63GR�ڑ ��� G��M��8?�E��p��:�LD]e��?�yB&��Q�c �,B�ѹ8�>��Dm8?�_/ ��j�o�/�[Y1g˵��A�Ѿ0L�Q�k��sxb��|�.��� 9���њ���7 &?>{X{�SO'2^���tb-�*�𵅪�U{LM虅= �o�4F��wN��I����pA�8-�#�5�S��!i������bv��7)"����]γX7^���@,W.����N����u�� ��ƶ��{lǑ����jPg�O+�?�1�$�$2W}Gg������=a)<j����KI��i9rsF����J2}W��e�H��/b�W@LyNPފZl���1>�5�l�U��k�J�<Ҹ��g��"�@�֝uD`U�DK`'N�9�����72}��:~������Mӛ�*�
N�vP��im�j����~��%������P@��@r6Al��.�0ƒd#�ׁ�e�yb�8q/޳R�pQ~���G:��q#

W|RdE4������ Ɠ^S-����Lh���g�G��lL�{�)���>z�	�Û��XO�nwCj?�7���֥*m�� V��kk��~�Y��.�x:����+ea0�q9�9ߕ�>�Ę<Jū�t�Caޅ:9�� �<"�y���<�Ɋ/��d`b+��
i�.D�p���lq��� &��#*����|��r��I�xm�;Gs/�}$��yY bbA��Rs%-�Q�s!^[�7� �(�<$�c[��x\�H�*Te�
��b%P����=wn��?i�1Ԧ:4ߕ����b�(��
�W�o@�AG�,�1g^�rE�ZY�eir�
�yh<��vDe(�ə���A�bߑN���(�O�	�]���IΥaT�����R*6K�����#���S�1���UŤr�4=O-�i�|B��}k�I��j��Sp �?����z�	���-uI(��G�1b4���7�.f	IU��_��	��d�*�f����4&d1ڧ Fj�#og�[/����Nq�~+b�WH�Y�8Ȱ�.���R�Vu�e@�������$V�*�ڲ5� �eFЋ�^�Z�-����{�^�Ve��L8�t*4��m:5���@,ݣ�e
�E{��ɬ�&**#��~D��x�T�q��u������9��z3��"��P��|1������%HsPL�."Kɭ�b` �~���;�USˍ��ɰ]9���J�n6H_��^��O��۷*���&���j��%�@̎ޏj���;[eҨj�m ���?������::{�M������xP�|���U�퇽`s!{��d��Iױw����Ya蔱�NE����m�?[S�����8#�G�4�-�pŬ5l��g:��cjc��:b���2[�mW-�P��%O���C�M���c,��˴Gg�<��
h�~ɻk"����U��su�	���Pi&Li�ل�-(�|}�Jb򨺛ψ�OHmQ�*1���L��� ����h���w<�� `�+$;do�d�Ξ�++{{�v�앝�P!I� {oYǖ��c����~����u��}�}>��d�ߖ��0)�!�?��V`��P�ܻ��r���=�I�
�����@��,nx���^�c*yb~P�"�Z��T|�.b.�$�-�%��$�ӣD�>\Ư�f�!1��������~��i#Z;,��u~�/R_��iҿ��b�.�X�^�(�ܖ6C���$T ���ܾh�K9�1�n��S^I/ �Z��'U�ߵ>O�7!k���p�1�R/�-��O'�����#�?\��J�Vp����v��wq���<��xC݋��C"_Qi˙n��2'�s�3�c�T>�0D b�r����?���~�G���ɮ(��i�M�������ֱ��^=S����'����S0��F���S����v�-<��pBfы�IbtW���y�8���e��OB>����m�du��+A1_�g�a�#� FY砷)�uI|0�p�)囬 19M/�v�:=�3tKx���T.����'d�c�p{ei��zb"�@l[~y|@�o	[)Xi�L���o�Q��p[��t�Tc��;�Xh����Hz�=����S�O��r�Pb����k�!9S�7��a�\��A���cP�*M%뱿4_6���&(V868�VD�'s��+��
by��k�,ڥϬ���Z�Ζ�@L�!�{�ͫ��/��T��>���5��4�a�0��gh����jJ��$����Y<IdXzڈ��km^b��o#6�S��=��>���_ 6"�Z�l!�T�,'D��;�x�1����wBc��g1�o�=:�HI���Z���7Ia��	�ͤ_>)���_KN_�� �:���$!D�'3}<a�{-n�,�(d@l!���B���*SO�"���[* F���Yfs�.6�-A����b�zr�����ß�Ϩ�HA�:�g���|ͪ�'7\p��9��t>jd��<�#t�����d@�kYz�������~�� =+�o�Qc�/������!d��68�@��z_�?ŋ֦2*: ����˭?p1�	���6�/��aM���&��QY�����e4Q��Ħ�^�-�bI�v�F�;�MڂX��������KDC��9�5���>�%���q�/^7.7[ӫ^�b��/��r|�S�6�gl�gm;Y�XZoZ��:l��e�n������ࡘ�$X� �iq��b1FvQ$k��ԥz���[���@���{���u�x���Z��CG�R;
�'{D��M�s]���L3��
�\�be�n��s�?�I����{=)c�Lp�o�+A�6DL���\?�����{E�0�{G���dE�u<���Sx.��S#�Z����a���Ղ�����퓪�@��[b��b�|��K8ӭ�AŸ f��q����NM)'\�9����|O1YM�Fm��d�҅>_A�����zy���w�!�����WB ��M�60��&n�c+v�K����DG�J�������6��8�D@�s��۾`IU��%���M|&bvP��_��̗B$/�*�#g�VAl��77��u��i�ֆ�8�/ ݫIPwarm�:�v��q�^	b��g%[>~���f�=-�I �.gcb��܊J~���6�/1կj��.����V0K1�}w'K�&���PF���6�����1$Eߢ��j5~hl��� �}�.�k3�oo���g�:���~�
b���U(F����\b=D8<a�@�@Ъs1�P�'s->�m�h��7�����n_acI)��<+�|�F�b-���y>���S�Q��B#3�����TenJq<�#&��S3A�b8��6���^����%L�f�7�MO�rުjy3��=H]�d�vI�FboI�o�J�U��х������ؓ�����'���h��4!������_��������y0mo����]�$�
#3a��xBQ3�=4\��2]A��=���xH�=���@�K�����_�_<�\9cV^�eep&X�9M/��z,������:Y�/q���>{��K���>��_춯�?L�i*=s�3	)����l�b�>"#ss�!���{��;�t�z���X��#���7&���-�_�}��K<��k]@��f0�5Y<n�!�,RS9ol���W���N�V��qwA�Z�ꃶ9��	�I�x_P�$�wR���P��~��W{����C��V�;ʙp��
&r�{̡dL�L�l��rU����W�{ޭ:^����5���0���ؽ�����ڥBB�6�L�,yĭ=��g��6�p��ui��o�����6�o��]�^!�b�������~���x���9ӻxV�f��¶|7a� bL����y�B��^����8^��d��W\.��Pq�w� �����<��$���j����)�u�'E� 5�S7���C��Fd@�\}��X�%��e4+�N$J��,�5�&���+�G���n��'b���(�.~��|#�i{��>t�Aզ��������R��(�	�p��Nc�� ���x��/-�u�@�g>�D̮���˅�{�Ԧ,�y��D�d�����R�-�^1��-�f}S��ϯ����Ÿ�H�e��`^�)��#s+cf����yͅGұ���z&��� �D���Z�f4Hb����ؓ�@LY���߹>���^⮇$Z�A��`�@�̀B�a��C=(�b�v'ŨZ׳����X�"v��@L��X��L��8�|�F���gbȖ�i���+F)h�)zQ������^�����ě���[k���d=�փ�����/�%q��SA��K�@��b�Ԗ��������	�xZ���ܾ�,P�]�gk(mX9��X�w�/Ɔ劦�r&N��� �����p���>��b�A	�b`\�!cn劦��5|�c� ��䒍����>��+Ϭ�
>���R�%�}_n�j�J}��H��}%�|�$l�p�1��Eަ�������G�"�3��S�n�E�/Ȁ�z0���hBbvN��7dy��:�Pw����w�l+v畮f9@�{�/������C�m�'ĉ��I�}JF��ҹ�n��d<k�9��ةd�� A�}q���=���� �!:f�= 0y������[Z�L
d��L\�Z%�"���������(�d��[�����+"�yh>�I�6kFT�M����.��SW=��Oz���_V�U��|;�R��[�Y���htbI��y8C\A�����9h��&(�w���gC�	��_:Vh%��379���z�b6��d������F��j?�@,� R#���~�ե�6�4*�^�q�y��SD\L���UnM�؝"m�
Q[C��٬����i�� vN�Q�-'A��ݐ�ԌO,e�� V���N�Ǉ�W�3:����-bl�q�+���|d��Cx~%>�g �F�Ҏ��#�3��	"�[.-�)��H&	b�Gx�P�DG�v�m��X����8v�T=6�ָ�6K�T���������y31�-�i�6��b�[~�M�ў���G䣔8�YA�-)�����~� ��W�CA,b������y��ި���x�2��H��Ɯ����Ha�?�4��1�x/͘�h�'KQ�D�+��h� ��D�=�+��A*�'��s�{W�NO�v}S��>B�"��,ӄ�b��6�r���̿�m�v5��`����7��+yӻ��%����� Ƣ��W6?����dYGÙ �TJ�2�e�lvBb��;8�}] F�$9*�}�"/���Dq����5�q���U�c��L�CpͶ&"� 65�_Τ��w�16�~�����̘Z7,���S7�R����-}�k���7iC�~�=�� ��:=����i�ImR�܃~�?�e��2n� �Ѽ�R�-���=�t�U{���v��G�灘��S�{lm�l?�^�Z�d�T����sb%��{�#θ`�y��YĂ�%{�f���՛2�8N�@���Q��]�G���s�;)�]6|j<�w�r$r�'�#��Z��$�rZZ���ҁ�����w"���t���w�x��@/�Cs ~n��uU��_�x���B�P�M/��I9�	� f�z���7�L0�g��\N%��b�%ޛ�h[�()�N����ko 1S�Yi0�.�lF���M�!�A���1������O��S,��e��H����n�B,���S���r$�^E�!u����"�r��X���<���tDNܼ/yy|�F֌��+T�D�:Nb�~t��O�X�����X*�C��4���@���(�-�� �J����F[-��u�Ԁ�^���'��2���#6U%맏 ��?fm�#�.}z�Em�+Yb��6e�&vl�wxq�:D���o�XR���U� ���GV�,h�G���$��5Y	e�y����況�D�+7=�4��T���Y�Q:JK(LZXj�*�{���,��Ab��+1�9�b��=R�
E�/@L���LC��W�sY�Q����I�>�Ee~zLm��r�Q]��S��tШ�M���L���%�(�AL��	l�#�J8��O����v v�:1��nԭB�Q2�y��� �}�@��~�o@��3�'t��A��}�+)�����j;�i �c��W��ڤ�\">Zk���ë��'Q�J�����I	�T��s��i	�4�|�`[���HE�Y�K�XA�}t�m2]8|�ž��a�y�П3��Y�]��{65����g��b���$E�o슕�/S����"������Ǒ`�s/�*��O��h��N�P6��$�|���}R�&�}	b�m�_���e���Th�%߱v��|�T%�o��zҜ����h�+�͙�N�%d���';�T�� b]�N��>�_�s�s�\�M�;�i��I�'����9G�C!��
����ӛ�!{��Z$�
��oߒ�?u����@ĄX������t�La�;B�dX�n!7ؿ<D8�,���ySS*x��W����&��/ۤ�"�K�햿����f�L�_[����'�`�;!�Ѱg�Hn�?>��ٰǵ��޲'�TD��C��[��(��次���T����b�
b���Yv�T6W߲�O���̺�۽��)��p�(�`6��Θ�Y��b�{J�BO�j���H8�w��G����o��}��z�!c�������J� ��=̧��V�m��v��4�3���-~y?�8sR�D)�֔��Pb�z�����2[Fz^���T��>����ڵz���56,`�+k���5�5gk�v�}&k�����wͲ�x� �ko�Aߌ�]f�d�����s9r ���WW�`~^���ɷ����Y���'���+=�p�"�� 1��uw,����i�ޅ$��  �}�6�����t�.��m������zh�� "�:�K�|V�J"Z`��s���}F��VS�7>$�)ڭ�bb.��w����bK�[�P8��nO�D�W�0쟬�?�5������Q��n1���oN/@l�ԯOoR?=_V8�!!A(��DT�"6��}}J�~��uC�8��W��V�m��/��q��㴰�|�MǶ��J))>���p���,��� �h���UT�@Q	T@$$E�;D	i����.�$�;�$�i$$�N�~:�O��{�CӦ�R/bl3.���I�exi���](�_tS��zL��5��b4�	Ĥ���r7��\�4����jy�����T��zE����z��Ġ�F�2���{o�^>LF��=�;���� V�ӣh�TO��6�E��!W�
�4�Ζ˦yv���q_��S偘@��@�O���mj:��(�'=� ����c[��F�� �$���$�gv%�W���RK���o�,W�r�c�uu�Ή7�V�� �
�u2�+��H�Ō(��R�����~Mqy�l0f�x0���@��w��=v���?���.����"�tL�Hu_wZ>�q<z�DߦIэ.��&���1���Z��`.�I�j������fF����b�k|Ÿ��R�'3�O:�-x����5��m���g�ۣ's��''c3&��t5ӎT������qJ�����ڹs��d�睜����L��������i8��@l�	�U��ڞ/���� �^�,�7ś(��*>#XA�=��~������k���}��px9(&�iS�����k��<�\��8�ز{i�;�� �/mI��L����/����g��.�h�4z����Q�$�7ID�;��}3�â~5I��\&}���w�W�	����J�5��.�>[=MC��l@�6�>}m��ǃ���M��]�}6��Im��>O���,�ao�`��0<_�!d�c�p�X"�ɷ�� fj�v�� K��e �\��Q,o&�D;���4�ދ͈�;[`1���\N8�:�ɷ�Q��᫡�@�[��`;�� {eM?ii��n���e�{���_w~� bSSϚo�"�Nx�G�Æ�&�X�!2�6[�J"ߘ�-3:��$G�bw��
��3�m�<w��-��f���qoܶ@�E�@��}v�Y������7퉑�(���
l�.��&zGW�C���{Sl�`Z%,����_��>��t�~�ׅ-������z`�{��{l��`l$͚ˆ����X����(�l,�Nt�`�>Q������/���}�bkg}H�^�A��8v�Y�@L,S���3}1�~.��C��}@F�r��rҨ@tEւh����2��8+���"/Z�'ndlã�]9zbۭ{��"[\�5�lW��QU��+�C���ִ�c����w�8����x��b31P),��ocFwcл�Pd����	�{8.|,�_y�>w�Y)���O��E\��7�Rf�nE���u7� �SMkw�h�kͣ�'���^�Y�gW)-U�W���"�ٵ6s�O��rsz�X70k�c���7ͱ�������=].%��h��W���y��w� �V8��7�N�*Lʓd<�!���Y��qh������[�w��wk5���1|o똤�{Ʋ1�H�W�A�,%���ܔs�ܸ��K�Y� ��;h�����XɽϻM��ce�;���}�p�
�1��IZL�$m=r 6�[�o�.��;�k�/����j�w��ޥ�ܕ���e�f%U�
*�����`>������f&��}���U����f,*|�M��WW�}���T�:���7�ƥ�<8��k:���_��"�¬���f��l��օ4��In0�~6����$�&LĒ�ab*.��K�9�p2!Y���.��fw�2�O�J����q.qs4�+�E�f��%��FG˙=�����vQ	�g��[�yNh���P&��g��I��a&{��k�?���ąJ�[5V����� �F@��.���ʇ(�W;�{ &涅�F�n��tK�.?����Y����=�'^�����.$W�+ 1�'T�2Q-(��=���G�o�Ѫ�`:�+��	�8���]R*��� v��.F*�:%ʦ/�mL��b�B��!�П�L���4;&�12䳂[{6�Zg��0��z�p���MI�����ω�-�T
V�c"��ؤMG9V��p��x{��)���k9�l�!٤/��SjWȒ����SW$�rރ7��NL9�YD �fk?8�@�b(z�ċ����#d:S�JFƹo_;�j]k%1���Z��r6�,�]��ʜG fr��N�pxZ����V�&+�`�ďǶ��3]��=���k4I��aG�����2xd8L4q4kr �k�����1��	�s-�VУ��i�'�V�C,�{}6\������
bײ0^<!M��	�`��~ڲ�	b2�����g����g�x�X�1K�{�
�h&K�
(<G�|6�ʅ��UתV[�\�L�}19�X�x�0@$9���>�1��ı$�jؚC�V٪�5��A�r�Ld)J0T�r�V!>GI�����0 WS�f�<ҡ/&�V�W��k޶u��x�Q��w<,�A,3�yUό��V���-���"���J��=��J�t�gqQ�A��D%UH~Ld�0{5���O�@L��o\����(�h�%5ayW�8���;%���=�~w�c�e��}�n\_�#��?|"d�G�v:�!���y;�Yb4�7Fy
� t��a\�����w)G3P2!l�+�D=����,+�1g/�� Zc��c[`���y��%Լ+l��r�n��	�D�[-l��6��bL���͟���kl�h���R����*��]bx5��)����Xp���9�^zo{
bx���ȯ��z��n2��v��XT㱎]�}��C2&�k��	Z� �m����� J�����f[M��a�6BH���1
%�z3�@w��5��ĉ�L�t�7i��Q�F�ȼ/��.ߣv�¢�\�/����@���h�]�Po����
�_4,݂m����ed#�\��Y�[��d�~;n]�nNăfߓ3�M��]!�U���+s��.�ೀ�p�jT7y鲎�c�f�Qó]�&�G���g��M�+�;Z�1�.G�[o��iP~|HGWE�N|�#��"��wvT�I�R��y>
b4�����Ο:i�U����3FA����0�w�j02VW��Jד�_��}�(�Q��Q�'�L���@��,�j ����p��V�js�?����
������}Ү���:' ��F��r#�(�:8L�����:�ݲV'�<�}rկ#��t�Bq�Ġ���Q;$^���~�/�1����橝Y!�;�T��X��V��4�MtF�#��.2S��Z�w��<�kz+��&�?-Ϟ[�bp��.#��(͗:��c5n�WW�؜s�B�\��A��<�Y���Z� >{��0����V�r�E&�e����=P�ŮdxA�}K��x�y��QOBEq���i��(H �(�H�c��9���e����A���^M�S��v ������eK�Li��<j��t��~j�
b�I�!���]���IC��� �m���"s9�r��r��k�J5y�~F}\�#��#�X���aebm�N����#�'��.�d�R�� C'i^%�H;?w�5Ƥ�#So�/kN%w[S��N�T�������t�<�Q;g/���pˠ+��@�/ް-d�c��M�S/2�RRw�e����;�3) ��f��q�~V~3r�����E{R�k�1W�s)Hy�R��~�X%�-�iʾU���c~��Ȟ�b���Mj����&r?i��)J ���PM_���	W���i�:w@���\H�A��>��F&G��4�[L�;���>S�T֝X�F�Vb4SӺ:����gʊ���d� �lIБO/@'_i}��a�Y�1��*�Z���3X��\�Eb�Ԭ@=TE�y�k�7��d*/;�!�u�jJ7�D�o�a�T6���C��L����v���˱�&�G���x���W�JW?}���D��01S��T8[s��L��;}�E� �G���N-�d�S<�ٮ7�b���\y�fKw�C��iY볁X����K���*�]딉A����0C�9p�Y�lw!ҁ�˟?
��2�����QXw�@���Ԁ�R�����ia�
�B� �����r�jX"�'Z��Mcl	�|�y4كQ��H�L5Z-b7������uG��Y�u($AL2V'��
��th���b��M%f��8xhK�����Ą�mƕ�Bۢ��$�e�G�@L��j�e�S�ŷ�ʩ�<�_�رq�ۗ3��BkI `ьsy@����%#'�{��>�ˁ�X�?u��/$T�h7sYJ�r���h*�ߚTs�������@�=z�p$K�s�\�4�{���#>�����l�P�x�F���ͫI];4��A�JJ_�eE���h�.\��4b_�s^��]�1��Kw~8��L*t�j9�Y Ĳ���BB���9O�X23h�Zh���^�!#���R/|3��+���黽��a�(�z�;[S��v���C��=�1�O�?�E��J����\�"֋��W���� �1�V9F��H^�]��wn���g�!Q���~��'}����R1������U���K�7�+!���t��؇e���cYH�JM�Æɍ�����2gF1S^���Ɯ�� �М�B���1�9�٩l^[%[�q�C�{�H}qI����Y��i/��wm��<��/3���ڇ�V%�9��l]~4�H���$s��jF�<�'4�ļp��k���iA=�U�׏���/sC��[N�B��_��h�jea���R�?���	�I�L;Z�`ɰ���@�܍UK��Bv���#�"CZ�?訞�T�Aj��������[�i,[y�(��c֐���;9�o\���%�5O@��H&8����}�G{<�ԫp"���I8M�-����2m_��f�G/�r:��r�����y�Ga��:�)H����ᯕ3�Ō������v��{����!5�=�`������k��Z�\w��������lm?�nQ�pпZ�4,D���ƎW{�]�Y��Qj,��h��%o f���I��"�8�qo�n�7��V�����A͕��I��XJfo����Ƃ�챑�?�	_ƽ��Wz�$��nd�w)l1_:���(㙫�������m�=q*�(�L�]�Ő	_I�8hٳȊ�����4�x�*'���ǲ��;�~yg6�̶�KB���܎c	�>w,22\���6��H?�%�I5�R����v����mv���\�R�_�6�IE�[�R�
d+�<]�A�6�U�<�����o�!_"�0�E��F��'h��Z~-��O��tZ+Lvx)�"ٰDh���H	h��dSa�?���jR�,��Y�gGB�&r
�jaR�	��z�"��!G����^3�*�㚁M�4q���[��A�s��Ĭ�k�)I#^u$�ǡ�r5�hO�"����v�[�ㄽ��[!,�?wE;p*��&�69��=�^�\� ��i��;�,]'0�A�R���~l��9{n����ǮO�tb�߽���a�Y�p���!��Ɨ�A8��aJ�[{#��*oP����vJ�����w��G��76ݯ"nV$�R]j?�=� j�v���2�b��\�㼵m��ڃӑL�5#6�s�+�P>|�f���J����+�P=�H5X6`��qQ<�`}����@C�u�*T���"hK+%9��H�{hV%�l�q嵇�$���Au��e|Mv���eL��g33�ֹM�#�.%��2������<G���G��	OǢ�;�E?3,(D�5��"d���J���R���,)7��ʂv�~�M	mkNڌ�?ؗΊ�)=��{z��FN,͂j��,E�{�+��`:g���I��:�����̐����y.�T��UxY�A۽�W�:J�N��^L�P��������;FO��y/-"ccǧ�2����b|�n�D�aً|�
׻G��Ծ�Hx�Č[*gwsE+^)�Ѥ�1�M��l�?���b�l���ѡ��eS�H�t��-�C����3S/X��;ٟ;�����_�^͎���5J�T��z�ښ'�?�\�tmm����#Wa���vNi�-w�t#��UG���}/�o������f_��N�YE�M���XT��m.*δ�������>nB�xej�Ϊ�������uXV7O73�~4k~�K70S�^[������hI��#>-������]���ђ�TR�F&#Y�0��'&�N���W���2�y\�H����b1fz��F�k0�t�d��D�:��I a$���1y�Z��[5�՘!H� d�s���yۿt��L����Rk���T�v�ȝ~hn���������G�9cQ2��e���Z���?@�n%F0=�c��R״W�,���E��;Z�������[�~�zL����10��:�ԝf�?�]d�fz�1n�9���4�3����4����؇��ԛ�|vb��+�48q�ung��p�*Qv?v?������fEIW���~��m����]���%l��'?��ְ��~���!I\.��!N2	?�M�<=8Y�@n	�� �^�/���zB����H��{���tm#�-~2�j�4Gc�A���/�3>N��.[�˹aL<�I�V�A�jݘt@�/�w�-q}T�"���#y1lQ��x��w�rÉ_!��
=�%UL�PCq���0��n>���[1� d��Zѝ����~���x�M�魌Ծ)B�tc��Z��#c��z�N,�[���8l9���%�u�s��(��q1���ф�$IjZ�]\0�-j&�L��[�����Uݧ3���O.�P�^���F���������{�?t��ˑ��َފz��O�k28(�r��~F��X��L.�����a��VY"������㘜Rh8�)/�n�߾=3G��-�C7<͙��+&`�������Εitw��9��*��Bg�6UJ�l������:�P����[��h���eXh�@a�.	I�����Q�SZJ�D$E:�		���n$�����w����9:�=�ǫi��3?f�Q�*��RQso����i���hG6�5
������<���<������Z�zu��C&ie�AW�j98.�Sbb��W$�,��FT�o^�~Z����Y��y���e��U:<��xS�#Q�*����Ħ��m�*�N+y`{^�1M�2z!^v�cک,���b���	�}�&�S\�)���j��%_N//_K�������s��щ�Ȍf��[uk�F�#��c�C�B�Oͮ�n̥jI�n�4va׺���輪��"@�̲�Xf�g�smE^�:�7%���4%nu�r�����7~�wPٻ{er�~:��ݖ���1�+�V��旛�;h��������.F������MVV+l��-b���Q��Dا���ZUD��X5L4�>W?m��R�p,W\�Hͭm̵Aүm�ゞ��s}���RވK�5k��Bo!���l����ҳx�w�PH�g�qs��66\U���a�t��mǓ�.&�韣��;��<����iY���ta�ɋm�&F6�ɰ�k��^�i�&�k���IJfR�o�]�yԄ2bɴ0 ֽ==�l��G�uD��^��vJ�_��6���"Jʓ03�����-eBR`�x��������B������E���W1:ǆ^/~��L#�i�8=3s�ۙ׻�f�+'8t������T��{�������$�8TD����ԗ!9� ?�� _��2WKM��pcӾ��<DF�T�$�'H6K>�Ⱥ�>�!���2N��<O�i���B���z,o���&�1K�v�LX��K���M��³�����'��n�r�r/���Etvu���!�|q�g�r	���V)�֫�"�)-��Ұ��o�B���|�Ikl=�x��n��V��m��o##F�~�=����v�Zԥ$kO8ȱ�د�ܐ��Mʭ(�P<��66ʻ���J��l>F̋k�d3�s���`5!���eP�A�=�1A�"O(3�W@��aHU�V�onH���{F�.���e.k��P\�(�=��D=��|D!Y�6̒e��/��xW^�} �R}��H���4�O��@r7'�x
�
�y7jW�GG<6��A,�6 � B�F�.$�O���U����J���Y���`�m�f�;�7a1�+��m+�lg�����s��xK���C�D��'����"��p 
�AӐ��了����!\��̋��1����W�GV(��w�=+kBvAl����8\Ϝm,1٦g��2���㯩zPKFl���M+��j��X'O*r� ��l�XC>�ҌEô�U�"�/�~��ҥ�Q)��<g�q���w.uO�R�U,J�j@��3R!�)Ĉ��qg&��y;I7�=�������X��ϊ�1xM�݇�K'�(RW#-<Y&� �8�Lf�^��ײ,���S!�A�����p{5N��)�wF��`�X�R5�N�w��`[uf��3��E�/��]��,�IH���X=}b8I��6���pp��m��
b�Y��y�X!�+�_�E2��A�dΡ��v�D3���n��"�u��|g�@�eo�Iձ�3�E�зҼ�r9�vs�<L��S��]^b�FT��QDM"����I�'~.1���0{>l~���=Ԥ� �<U��#��qY���H(����^C��+͌m2�SV���D#;	�b٢S�h�)�IXN(�8���� ���ɒ�%H������\=�Y�6���mC�' ��Щ���1A�)�Gh"F���KG�q�\�� ��ː�)�V�s�5B�D8��Ĵ���2�"]�)�-.8瞷���`��_F~V�6�C�5�����v�?�̹X�@�K�qFTG[�����׭�
�lr���UO�)��Alw����
��:q&'��5�|@����Z�R�f���d�lDh'#S�|�[����}j�`d�d�bOl�b3��H�`һ�sCÂX����kL�e]������� v~�f�����4"���]vl��� &�f�-*}N���w�a� b۪�B������e�=����� 6?���x?�	�����雘Y+[:e����ZS�&r�(�7f&b�4cUN��y���o_�ӷ��ع_Qt'��hs}�Q���� 
y��fQIf1�"l3X0g b2Ψ}�SAb�]������A��w�Ĳs�y�r�Mw�C��N�>_��	�hؤVbj[<1�7����(����bmu���ؗ��!�Ӗ�;k�[pR�+�P@,����4�-Rgv��t�?��y`�B4��a�����u���m*�;`��)u�
l�a�T�ik�AL�E�*z���E��n���@e ��WE���ޑ��B���rH��� 1�yi�Ƶ�"$�e;mQD:�/{���8�@��<�dNϤ�؋����%5,��AL2��ӽ{C�s��I�ߠ��)����7s=��U��繰�1�N7�'.4��jo��Q0�j;�芖ӝ�)���Le�ͧ�� f�^go��qE�e������tĐ�����*(� ��.U �D��Y����a�qkN8<��ѳ�n�-��h:�u������Y��د��P��f�&_��tT��^|� v���F�!���[Q�)��b!<{���S�1�o�'+��<]����g����,���j��R��|� ��S��O���_l4�A@��`�D�f��/�_ل��#�W! ����&U�{a'�-y���Y(���9��c�rXӞu��!YH�K��31�.�U��js��ܼ^��n�=1����?�#�>��F�[c��1��Z��C�{�r�t�`��ءF�N�7V�׾�,?بq�o� 怂*t�@��,W:�)x��!��	ĤQ��?�@䰟��3�s��b�V
ɟ�$�)�`˗8�ʐ���M�"Ӓ���lcϒ{�y��i��
fqĿ�3��L����|b,$N?��n�d��Nw�¼�g1�ZIq��}m�8إ�W��:.P FPIȦ�e�I;�<v����R�Ҡ�_[�T$�����ʁX-��n����Y��s���-�� V�s��h��=/�g�L6�T?&�4�7���uُ���78��$pmA�ݛW>�,�%RO�&�]J��A,����\���!�����kz띮SH�c�n�@��l-xWIbp�XXZz���U��݃z'��B�a;qp�.�f���n=Q
�6�C#>9���,q� �@��S��b&�y[�N�;��<����2�;_����)�(�V]4�K���*)���3��XFE��=�o�g�x�,&�����T	NU����c��o<�$S�a��(w�omj�#����\�E&�c��Ѡ�0��!V�������w��̠v?�rZ������D�H�>���*��_�kHV����`	�(��z�
>�hS�z���Bb[��EV�o���s�=+�	t%_wY�����w���?����	!�vs]9���T�?�zJ$�J���>�?:ǣHͦ�u�]��? ������?�8�W����} ]�q��N!S�����w�ң:{���յ��Ώ��g�%ݮ�6�/�����P'Kjk������bq�v�-�֓g��q>���~�o����:P�{K�����>�"������y����s6/�U�qË��TV7;e,���y8%PP�mÏ��WW�~��5���50�H�0�#0���[�d2���9ˤ{���W��/�u)%�|}��Ȗ�/1�-Vf�&�"
���=5�{��i��¤�]�ȟ^A`�xX�%T�����k��)�1I��C?#��2e��0�7�NiV��oϽOl�ϛʦ���1k�[J�k� �[ͳ�Z��{Y�C*�Vh�,��4L�\~�\�Ӿ����[�>t�	��L$K+�_�u<2��4�Lv�g��MbV�|���;���(�S�)�n����F%�H�2ÁQ�4[^�fZ.Y��Se�'Z����r<fj)�Tt~�c��a#��}��Q�k�������n�%��ğ�є��L��~=a6��J�jA��0Z��>Z�����J�iF2Y��ø�'���ex��#��F���g#~q��*�:��[@��R�s)��O;���_*������5M�}��oqB�V��؀�|����aqs@�z��~�s�_ލ����X��섢�}��]�����2)XB�mA�\������;R�
ĸ��(�Oך��ϲ���x	��*���.w�u���-�sF���n�X{�T7͛��.̂9ѵ�a~2��Ϻ:�s�%�_��a��Yk4��K���e�~�ߤ`/6Ӿ�Yq�g�-�f�q3t$�."����㴩y�7SŲ��}b����mi��<{wb�[W�Vu#޺�l��y�j1b
=�}(2G�M��d��.�1)�my��2�H�%"Zٮ�k�{����+d}�I<a�QGs�<����V���ɐ�Q�L�2,�C7���_�V��Q)�9���_�����a���M*(vw��S��*{/�����mɃi{e�v�~�������w�~7;U�N����ӾU�<�V�hӊd1D��/�*1�3"^�o�h����H咯@������D�	���h�,�����F$�Y˕쮔e)j�q�6�ؤ�Ƥ�([q�>o/Ѡ=���s�k�G�o�0���?��N.2͋�r��a����(��F+�F�[�仧���;v�c�j��t�z%`��m�9>-~v��/R"�֡]�$'I��&���Mu��5)��ij�㘭��nnHf�2�o�$�@̺��Fr�`�<ꉔq?�"bn�_�^���|�_�Χj�:-���������k<���� IKO|�^�����ġ$���Gh�O[`������]��fs�aQ["���o>LxM�}���5X>�c=��ol
������F|�x%��(�B��pc~���1��<nm��z���/�����ӗ��+����?-��!Q:#c�b�OY����
Y��9�S3+����d����9����e�Ξ)[o�[�d��Ro�Z�&G�1���R��-���>;}~bS�tf�>���܅�&>frK���Ҟ��i��Ԯ1L׻�<X�}H�u'7d��b�c)���6��r�x�2v���k_�`�� O���A?Y��q�KO1���쟝y/V]oo{V۩E��q�`�����֑�rl��°旅�w�&n�:Eޤ�A�B�Je��Uߋ̠�VG�~�Q���>v��b�!seDcn�|;k,d�j;���-"͚*%�g[dD��'�2����*&��5��=C-p�:�B�f�WU.���;���r�z��q�C�R_�`)6M8f����^4���e��g�P�1��C":���iY�L#�n\���/~�w֊��i�	�;�z��j1�x	bs9Tx~R̓�,�}a�2�?Yg~�|���II��]���
�AL����qCKZ5��;���3X��,�<G1�ᦆ`ۗaa��5��>�弸���7�ܠ�Q���R�!�Nmh��eнĤ.5<i�p��@���;�[�%��M����tb(#{��/�5푓¡�LL8� �4WJU��h�-#�_��:�����O��z���^���>E19~*弄-2�	���KOf��]�=^������,!�/'�.H2�l��<oB��m-1#`u�E�W�_Ecz����ti���[�jP��v���׍	~������,�>)���߻�Ɍ�
���^��m�3�S�:��[۴�b�h KK*��>ʄ��l�[�������V�Hk���'�noQt7���B����E�#�j���O�Ь}`� �-��܎��z����N>�}z:�0����5�3���%�������-Y��	�<v�����>K*w�}h����¿ч�H5�C���
�|�N\����io5d�;���w�-L���3j�֠V(�l��9͔�Zޠ���"1�m�O�{�Jc��a3�*�F9�6.��x��
��_aD�B���e=����V#�q�8�9�9��ZA"%�"�����k�e�ǏA�@��;(b�Tpw�y�6����
�/�?8�^,�j4;8! ��[�9@�M$�f��}K�Q�����g�%�0{u��Ll��Ƙ'��U��iϦ6���-c�w׍s�r��U��{���q��[�W��IV"A1n�v.�#c�||���^���o<�nc�r���-�r�s�3t�T��lzWm�2�3�ӿW�����ݐ�������$��7�<������	����5r۽Ĳ����)ލ�1V�6���
�f1��9;{�(��w��}r��wh�@�� �3�)�Ȑ�4!|̼�1��jPT&�#�>�E�hy�M�uĊ뻐M�^ⷐS9���,�S�ۨ��|����.%�ި�'�Օkcr�v�
�n������31[�֡����>O�ych+t�;�"�Zۗ��P��R�W����Z]�2��ߑ+�S!�o�y)2�{�>�\��5A��:O�؇|��S��]�F��
Q��b5-��J�:�<�a_즺�̀G��.vQ�[��%1�^��w5 6�o�Cy�-���2���`��l +���j�ѷ鹐~zoA�*1�g/y)��V�X��[2
�]���NV(DO9�9��֢ƅn��6d���va��w���c�b~�f��o�>���A�}��~\/?b��f�İı��N�\�m��@Ljf��qcN�l	�7���Q@��$/n;�?1���'���b-��?�*��>COJ8�_1�0C/'�M�<�&� ^��N�#�?G�0~h���eX�¨a:%�EB�[��D��[��$EBjQҍ����%)"!%���qf�����y�~;H}Z4!���v˞��-`w�g�&M'ե��e?p6z/��X�u���e�ɛ$���
5m ^�L�\5:�s��ry/o�:<�&��Y�좉���������_۾cA�mI9Q��n5Y��b��-+"��������ɟ�e��Ӛj��̂�[�H���5�sRW���3�W��˧L�؎��/s�]+�^��]��v�� v~��oo��#����ly��k!�5\k&�{�#b���G˨+(bp��؆�v7�R]�� I-� [c�f������ߎ-W5@f!�CV�g'�m]���@�+�r��0L��p2�UOٖD��L�c�_�jϑ04��B�D�3�L��r<��W�Sj�:0�#P��+�Ɩm:�Ӽ�韻҉@���
=�,�7˱jf��WYJnP[�1��UJ�OԴt>�a��A��[伉7�^�Qg̚I�Y�+)�7(��]=�٤��H���3!3��r�W�56[l�����lAb%tz�]��,�y'�e��������TP`�]9��:^d�8����]�YC�ZV��r4]f:;���ߺ�[5���>tM��U,F-1�����R^��7��uz	���裷��yZ�$	�Ӹ%п��[��Z�������~��S��Bh:V�K���s�,�v�b��Y|�����.a?L�-]��:�U��'�-bBO"�I�Tf_�Ø7l��_s$т�d)������W�ғI�3�@L��7�&�~�#�'��m�צ �����FfX�ݕ��0T�z�YĎ����X��`�e�S;����5c�?�=�^I�>6;��v~|k���'�)r���3��QrN|.���;���RE;xԪ�3U�6�	b��[��m|X6];F���)�װ^ Fl�����:��s�J>�G%�b��R�ӎ;>3+��G��j�3� f����G����8z!���Ĕ�_d�x����b�o#��J�Xm�����g�����hLet,;� ��\"�%n�����h,�]���p���Gt���k�}�J�Ĕ�GY?J��^�l ������C@l�Y�(�K���Xu���m�)˽G�vQ�� �s�_AL@��������)���}/c+�@f�u"z��.�6Zz�`(M��fB�����*�d(��!P���F�x*]칷�i�&�����@�6�o5Tf.Z���=v
J�9&ü�ߚX�ۙU���P������	�zbY m]{�){6^��ij�Вy[ї�qJ��~�h�}�;$�ޮ�_�W�I��g���b�wD3E��Ï,�#�)�M�Alc�ݣU�ު������}h �xG��2��&{��r��f�M����ޒ%W`-��,C�����)��W�i��V|�*4\��-P�A�j*J��y5svb� a��b��wkhj
u�Ve?b��&:���*j�AP�M��j����W% fCQ�޶��h+��3�Hb�V�E�H�^
*G�CV^l� ��ş�T"^SȒȻ�AP ��Y/��W�P�C:>mB����Q�qDAW�lJF��M�����'��9"�$�Jw�4FQ,�Fk�4e9�ւ�J3��t�5�����o��M�ҁ���_\����dw�,G%����=�Q��3�SI�Q�b;�:�������'E�2x 3�K�HQK6��+㷝��be���9�LWՁJnn�Cj �uӤ�Җ5֑���IO�����6;�l�����n[$��ʙ�X��S�UsrNl��Fw���Ci-���8�^�8���o13��Dy
b��t��g�h<"��U��n�� v�.��f���z���1V���'- J�uF\X�ô='���f�#)F=����y]N�!�p|���pI_�b�wn��ҵ�s��x0T#�E�A�"i�������(J!�뢭��� ����@)�~���=X{4cab3�w�^Ac���\1�E2��y,mbr�&u�skCg��7�#x��B�
_���c���R-��r�k�U�	��_��������zb�:�
AOb�Fs����??D}	1�m��*zW���������o� �t#V�ǒo/��ES�m5$b�J�����VN>����3<ϸ@�諤��A*��g*�,ؙ!� ��'@����Rϗ��r: b�|�#X֩q�xΤ3����A,ǻ�� ��;�f�d�k� Y��:�6fE�1h쫶x?WvJ�	b
ʹf�|F������N�f� N�5�ɬ�%�~����%bI�r�Q�ƙE�e`�[�y@�拉i��r�'�x�݄��n�T ���0�034WT��Biu�AU
b��Ǫ�$��4KQ�ʈ��`�@L%F�
+~���_;��F"'0ĴJ��˩��Y=Vi��4jEl@,���ê�\S���1� e{(��Ę�2��f�y�C�Qh'��ʂ��7�W{|��0s"W��89���9@l��wQy�k��AñH���^� vϐ�%��e=b�?U�@rC�H ��O:w7\rO:'���=3���2�1��$I��'��Q�.hTA칕�)��}��|V�ɝ���B6CE��[��ѯ4�K�z@Wn���fe���T���n/IH[�HV�X��y!���꒺����S3�,Y���v�:U]��뗞����ͪ��O�Y�#H2����A�;��2��vp���z��c{���0��&�{�h�ܪj���IV^ҭ1���o�	����y���g�������H=,�G����Tˎ��S�����X��+Ա��Y�ݏS�ɜ}d�j�GH�@�bX	��,��UI�_Ǯ�H�͗Љ�c�4Y�רxr��	��ظ��7���l�f�KǉA>�A�m�B*��j��;3��c���yG��j�����F�x�z�$�JR�i��1zK����� �7�Ӹ����q������cAD�����*���'�@��TPu�9�TQ YP �$)�E�H�δL������n�E�b�&��}��|�m���#�� 6���?�-/�������$��Ȓ[�H�N�V߼ۿaRyE1����˺!�/��ӜF��dr��A�2�<ΐ\���ʫ���4�Qz�<�њ��Yi�n����*�z�x��� u�ደ�Ց�"��-ڒ( F�O�ͽ��bT�N܎�1�T�S�t%��(Cn�"�mƆN�fA,�ct]?�c=�\�w��s�� ƍ�N.싕�L�����Hyc��	�wN�^w��%��g���,�����z�Гg$��)�3�	�d�A,w�#:.q�WH����xڦ�x4	�p�QE]��##v������-��dϰ/�	B�86Q���W�S�u۔��W����V�}�J9k���MT��B�Tі�P�|�v�n ��z-f�Ҷ�5���:4�b���صs��]9B��K)_Yܙ=Z9$[�tmNc���I$[Lc��}5 b��o�ŨX%�EF�`^�?�1�L)}��8��ּUX��>�.��ͧC=�*���ƀa��X�R�s��_.��5�UI��Գ�)�l��=��WSڬ+2 ��PC3��r��d`�2�Y�F��Ĳ�.�p�H7�<���K-��A�2�E�z�Os�gUp*P����F���o�.���U����:H�3�@L̐˓�wi@�!=�YHI�������T=4�`�|�c��� �b��k-����k����fC��K 61��䨉kC3+�/��.cb阕s��Dcz�難���c��@��
��Y�����Z��M�'�bGHǌ��;9�䭇f�DpOAlO�v�4O��2�6<���Ȫ9�i�*�v��so��io}r�L��|��F����T��m�7��@L}	�}��'�H��;�~LX�zĄm�sY�	F�=�,25�U�@L�����Ƿ�,I�s�h9���+f�`%�G`�<��~�BS�i�Z�~MyY��i�b��0~�i�Tr��?�XJ�h�|��� a����Z��D�b:�)(CN��|��'�D�?�y;��b�B�8��A�{lU-��Vj� F��l���{2�˅��U=ڣu{�|��I�zeã��Ĥ�I�����-�g���Y�ҹr�WH@l	�eS�f��K���Vz�~-Gk]���0_���N��.&�M��5�.3*�;�y��&.C-U��I6�-7����~#�GKU{ٶ	b�o��U� �fn��I�)�f��9C���'6���6NF��t�!?(�Ԋ�����c���(��1{3B8�P�p�y��jר%*�e�@T��k�Q����Q7E������ݯ|8˧6��1�8^a��}��e���e�s��{����N���/�JuM�L���,�=��_��l-֔�H�L�>�s�.?�u1��x�b���٫r�^� F͔ϠcO�H�if��O���b'VN��al�j��'�����@,����瓽�l�ñ<[�5+l'�{E���P�J7�F��<���}C����Z��,�o�n�A}ּbF��(����d��Q�����j�!b)
63x�Bn�t�keu�� 6v^�ߍ��,��y��\�c���h�񂢆�O�����oi�)?�1L����C:��2��D�#D���5Vǟg:r�O��*��1��I������;�Q\EkY�X��Bn����5w��ؐ�H���� �,\	���X���KF!����-bw���E�^��:py�Ґ���!	bwfP-�ܗ�|����j/@�! b����+Ē3��XF�w��� S�X�}^�����5V%��\�":�U�9�vWJ����:�T�����оy��H�a�N��a�.��sh�F/�ݰ ;"�|�[B�T�WYkA,���Y� �U�a��W��~���5�25�kPL<Mk�%�b˧j14?ְ���Ҙ
�!��꣄� �54�[��Ý���,te�Qb4�8��ȏ�S�U�х;Ƌ���p7�wb�Y ��-�(�F��Ӂ���Ts�Z#v�ޞ�LN6n�5�U���Pg$��ߊ�[��Jo5���nTPk)8ϒsJo5�a��5��<I	��Қ5���Q�y��΄��j�o`�Y:S��������m#/�P+��g8��Ѓ�ݳu��JH���h���;�h}��U��xb����ݨ\c��KlYU�P%�Z ?`��aa�[��5~&�e�y�w'�(�ŉ*&��XVL[̒:��P�YB�!����Jώ��5��$��@�����z�����[^���$L ?:A�����5v��ۦ�$��P{��z6��	]��{P��ӄK�G�x�vh��<S^B��;�����	�8d�߶�Ÿd��Q2���;r9��B�=著͖yb忚Ln�p�K������T6�|GŘd�cF$*.P��Z�/��i���.��.H���Ѝ���<+�b���ä���=�����f�b����5E��c�qAM���C�맩��p|#r�!���XS���E�=�#��9�@����i@mVu�{3�A�b"o]_��F���	Yn����I��Td��P6�����i���}=�6<ȡ�^x�ᣉ�ٌ�%����ƻ�D#�r����0��t����c�/ՙ�k(�P�c<���O������g�-ʭU��Mv�G����<}�01JE%�8;vr2t*\9�07JE���HNF �4����ZyT�8��5��j��"QH%�!�IN�i��/�5�90��n��qC��it�lHj��9b��gq`������M����wAm������bx={W��Jc� ?y���-�p�j�P���{�T��袓і���D��*�o�EԒ�6�7�޵��:r����XP3���k{�reG�O�k0��`L���Ғwj)���b]V�l��b��O�Q@�5�Z�ߺ	�e����ǨPj1}��!��]a��(�5CSn��_�jF렖8JQumVA�G�\�>{@q,�Q�hl*�D̷g27��.;����������N��p�C�Z��,����<~�"�ӹ�S���`?]��o��&W����Z�����b���(��`Se����o��t�PKr[�0K���E�hc��ɕ��l�O�:q~������O���<��{	5��A-�Og'80.@
��>��^�.3)���B��N,M�۸��؛y�[�������l*��r����Z���Jǟ�_���ʙ[�SY羣�Vz�;3C�,�⮯໣2�*6+�j-PlP�(�(�(��}�����rX-�9c��S?>�M��zC�n����	
v�X6�ͲX��3�!Xl�鄝*Vr3��@�X��� �J7�<u"����'��:�����6/�s�8 g~���-�i3Y[s�y��d�^�QԚ����Ix����C;$�8�b��L�y��x�p+��Ϧil��Ļe���o��h��y(��g��Pt��ȯu��u�� z�[��0Pb�e   �  8�{���Xq#��p{���=��ݔ���b?<�[+�*pl~*��=Tݏ�������<��[�����4�}���D�ˋ}-vk�x����k�#��э�_N�E��l����tD�������"�'d�"Ʋg5����j�[�|6[�|��;�fs���c{��b���o�dx������E������Py"&�bQ߂[7_�l�z�RK��u��+WO��v��K���Z�Ŷk�<����͗��bPu��~x�1o��m�s��Q0&�4���+�~�o|��|��`�e_+Tw�$E��ԙ+�4?n�<1�UC����y�!El����`	W�|�.�I��#8;I��z�.��[�o��e�|��^)b���|�k�����r�܍��"ױNy��%��;�,�Tw�ڗ�a�����y�M�2�U7�O>vW��)b�������>��'�GA�w�YR��](-�׭���5��fY	΃��-a]��\�!����3�����&J,2,6}��J��նnz��>�mnA��@���0��ʺ��Ͻ� s�-�~{'P]��Չ/�'m���8���w>y>�����m���t�j.$1û��(,��!���&pr�1����޴�aZ�diC����.֕��X��ǆ��s�2L6��������s�110  �=�Fs��������l�:HP�   �  "%  h���eS��a$�E�n�V��$���A�[��ii	�nA@��A�,3�ewv�������G
�Z�d5W�*�3�(�����b��_~��N���"��Cl;x����d풯t�L�3���孯�n�F���- ư����O��BIO�e^f&�tH+y*t^@uY�"�.,c�b��i�{0��k<!uQKJ���hbu��6�l�'#A���e6����3�3֮�n\���I��'Ą�û���h�ad�m�nS������^���y�]L7\����L�G�k��Pj�K�[��7tdϡG�R�J�q�[��O����q�Z��pL1d���E]&њC~�7���`�qG��J�?x]�V�F����{-� {��I"J*�c��՗4�����<���'�#(�����+�2+� &O�Tj5�t�B��W}�b?J>gS�a{�B0z��] ��N���%����Я��ʄ4��l�igkN��.�׎eO6��᪔���'�R��q
�~�Z3���Bܹ?�9�4�Jr����8�I�9h ���zl��}�5lK�HA+�M:u���KM� N�7}� f�p�-~�Ĵ�!:J��Z���ĸ���zS�_����B�.��k�14mXq��Ʌ�X{o�k����!�쓘QV��D1os��R-�1Q����O��AN��Cm�*e� �=?�4-�22Hs��$�
oG�i�Җm����E��p���ļ�H���?�eܢW\Ah��A��{7̓���|Qi��Tct�b�~��s�Gx��IgO��a�E���� �ޑ���<�>��2��E�$�MLn-%,�/&i�����؆W����MHc��OG�eB��3�AlֱP�Ķ���*ڂ���4�r���A�yc��_�-0j@l)V�����#K9zU佡�n����P���-��R���(=1-V%ʕ�nc�F���C�v�p ��;�b���KGw��L��-���/��%�!�EKM ��$����J��6�����W�u��O��!χ��Vj�Sd،�ۤ-G�/l_��0�CYɤv���ٖ�
b��G��=�X���j�)��Q�9
�E1�%T�V�`Ϸ���?:���<m5���6�ex4qXO�z����WR��g�׽�� �q�c��+y,�<�[����[���#3YL�MH�ir\�^��h�s���9$�E�F���m^���I2��6�յ�PwtOo�MR�l�%�C3G-ԣm2�N��]���
��I
@{�8���s���"� ����䔁�C��1/�+Zv�"b9"�á�ހ��A��h��b;ҵ�2BU5I�Ws�mg�0*�4��	�[�b2x���.zo�Rn���}���mQ�oC�h�p�a���Km�M(�!����a@̷Ĵg�<¾ɸf��D����kb��8�{7Y�*�I+�M�h�z.��!c|=9���ܛ&�R���?ńV���$���t�~-�n6d��A�6<��L�D}�iџ]���_�O|�1ߣ����}e������0]
_��tk�F��&�
�9)���t`g��.yü�����L3�	�Ք�?�㿐�'�<%��s���p��+t�DK!��"��U���������zʆ=��)�*�}����m�BVǇT��fJ%V��J��������������T����G�{�:�_���1����}�r�V~�� �QY�4ĈH�c�'�H��>�4e\�=�y��٠'zN�
�vO,���bm�S'�7��K,��ե���_��C��uw�늯�|F�v)k$OЂ�6���y�gg����|#
9���<�Ŀ�{�!�Ī�u �f[� n����?���k2��\tƯ�Ewg>j?�X�І�&���mR��O�Qc,O�!ec�S,��]��)S��3��VЊ����,�@�������~�j��h�ʌ�u%_yHa�3�ď�1Uc��ؒӥc�!+}��Z��pNȧɭ��l;�m3r��0{����24�/*�/�0Ҙ���kHb�2�E �?��
�ϛ~��Pj!t�3�)�2�H�J3(EO���麧t�λ�j���a�(�T�p��s�΅o�`��s�_��
�~-ox�⒚�h�[���4�3d�qx�#.�6T� �23x���T:��{*�m~��A���PRx�H�?�*%��{>1��������K.��� ���6zՃ�T�S��s�"������Z��f������M�en��Rm���bu�|������~:�7X�������x�yv�m��q$ǍA�k{�}+�*'@��,�R�f�6&�z�������n��dS�S1��أ5r�"���@�y�0�)�۝e�U)�hJO���&��-�D�\�^����9S1X��x?��Z�S�$Vi%W�6�����Է��X���΁�(Qң���W�O&��Χ���7�G<�T+���[��ۂY�����kÕ./cO�[�2<'�%\1��U̪�}b�h�B�w�a.��1��xCn�
 �ը�w�d�bEdJcV��m^����5�X�Ub�)h�yt�u��د���
[<��
��k�dt� �~3��@c�`�)�4j`��E�
b>R�*�J�d�XH>-�V��1����1�A�4TD� 7��! ����ýB���l� �lVbDs����w�k�체�y4�A��+��xm�d^G�&��*��:�Qj}��nK��7b�~|gb�)�v�|�/O\�<kNKd:�Al��H���°,��hR�C
b��U�L��4B)��r��A�!��}5���*���F��L����aC2�$�9$d��h�,A,
�w��-<�e��o]x�YQk������G��\u��c��a �XKu]��U�?�ޢ���������`�0N�q�XɌ�o�9� K�J��ԾX�f�,|g��Q8	b�N\S���,G�&S	w�K��@��&�}��R	~��T�Բֆ9�����2E)R0�8�����耘tNe��&ұ��wM�ω@l9�`��ʵg9޷#�v9‐e��3��\^4�f��H��n�D�1��w	��_U֘���+�m��XL,�׎�\=�K�(<�["SL��q�+5���yx�b�%��oWwc,hloH��z�6axI�[�Q���2�e�$,�%����rKf�x�"�76�vCK�	ľ���,[m��)P/��_ă�{b��{w7H����bhf5�x�� v���?*,�jh]!������� ��7�deHq���F�9��CC31��$�g��ab�ġ��HEK�	��&oj�ָ�}u�;�YdX��*w~��r��cB�\3�'��>�:r�ߝ��Џ9Nk��D��>n��������~�P�Ğ��R���G���:�����Pf�����l[M����9�����H�K�|}!I�j�Z~;#F &1|/��k��{Wm�,r^O	b�����OƦ�x�'�O�@���b�E�i$�~,g:Nrb��,ŷE<{$ƻԶ�y(;� F(ZZ��չ�;1[�"��}� ��)���	���P�r4MB����j�*���Z���M�Hk��PF�5l��Z?��`��}ϵ�b<o��3U�3�����+8��@�ی͕�x��F*z�1���,��2�z)�o�7�.x�L�$">q}����Z!uI#�tg��	��G] V�_*������7�Nx`��3�!RÍ �=�zS�dm"�dӃ��n'u�����,�|����z�_8��c:.6�w3k�*u�1⅟k�)ϴpr��e�����y[�No8Z�cwjLYFv�uz1����X��/=;�������8ĺ��X}6EJ�6�5��������(*�٘q�PR6.iRkXv�"�	e�<Q~7d���Ҹn���%39�qȜ�����:O�O��+|#�0��qx�@+�rڗ��(6�I�5@LC!���/Zene���m��� �밠g���+��۴F.����4<k��e�-\>�	<|�?��	'�t�?�b䰓�N%�
��%Z�Ŀ�㥤r�b�]i�a�.�u%k�����@�@?�=
M�ԛv��73<-l-��B]���t���{
�8�Ӷv��A���$%)�@<�9P[�ӯ���ĸ ���{���0�]R���OA,{Q}�1-J'[�aq�0i�E�v���R�R-�e;%}r�
-��@�����e��kz~�+�N9�i�0���xń�th��*A�HC�&v�^Ԏ�2�'~��� 1��}�%�r,[r\T�)��J�_x)|h}���Y�)�S�xJds�`1�i2
�q�6x�i�<���jN�H��<䟊]r.��leZ��] ��X]��p.s�uLF�Il�7�p�vG�Mbz��`_br1+������V�� �q�u/��@b�]��7ݶ���m�k)\��k�C��`�����m:�WƖ�<�����W�Dl��{_}�;�A����I��Q��.�����A���&�U|Hb�x�a�Q�����y���D�����>~9��`�l����EIv��	(�8���5S���C`�#�f��|�f�q���f����'S]���%ќ�`,y���t�;e���kVNL0<����1�Xr"�<�$��� ������۝J���u13Y�o�L��8@lh8uT;�ޠ��v�X\�9��b�!�vǯ�	)e�M����I���C��t]ւ��Ȓ �\�������V�R[��Ӌ�� ���kL�q?��,�N��O��bG_�=�CWH�.S��{��S;@k�͗I��7������������bb� �aι��Д�m�XU���6e {��m+y�H^[y��o*���BP�r?R0Fq`~��&��󞠹�9�4�l���u� f<�u�$\���������P	�VܙB�1��81C�d��:,@��ӽK�/�i��v��� �Co+�¦LS�$�F���W�b܅)���8�j����E/�E@�Wm�O�w{��b;~���d�P�:Tx��N/��k�����`����]�iC�(k�߆�nU!b'�a������_-������?�����F&9����{i�鎻ch�7
O\�Z�Ē��?�8_�}o��|k<��b�~y_z*�X��Ό'���o?1j{��o��_�OVR�j&A,�kqh��AE�;������p	�h�u]��0��o�D����ALHb�����[�����rkL����Ҵ�ryS$�z�23�,�-�Xc�<���%E�����}�I�� �@�����fHk^��1�&�FĠ��/���������l$|��J���i��-��儕l�`�"v��k;�����nT��`�dC,!l��Ĥ��9R�8��7�,�mkAf�mḕo��n}}xZ�[:���]+�H-mZ��^��Eقb�R8�z�1>�7[����i�NFD�V��>�аӥAMcb�ϯ*~�Ֆ4I:�F\ǡ��q˂X���k��Ye	)Vy*��� f��V�M�:�a�^�&~��Ns^[,�)M'-�cN�Y���BD 1>�=���R'��P����/{E�@�Qy��A>|IE}e6�,]� FV�Gg�b��x�&�kb_gbj����'������{��v��� $m`hh�)O���$���X1#?�@�d�\̄��������N��脎�ڳ�a�Y�+J{��o1�,r%")���i9��7�c� ����w@_w�m��#�7�,Ĉŋ#3����9��]�w#@��p/�v�!�&R�M�1�G-.��$Q"���e��'�}b9����� v���z�+���vj�;,�����dQ�}�P_sۼ���e� bk�pU��*m�aP�.��;Yk vd�����_^�rFg��ݾ��(�7̽�>*b�c�7{Fk�ԁ�%�`b=����׋h�4��Z�E��_�Z�&�@���j�M1X���!��e�$�SO�Tn:㧂��-��d(��-��A
b��8SN��e۞p{i{�5$�z &K�n��ԫ�n9@��:`���jc<�G� ��F���ȩ' 1X=�]�IJa'��c��P^�GH &�M��j�RC0��#�,i*O~bo��I�/Tqn�}�~�m--����@�sQ��KY�ooNl\V]�@,Ϣ>A؁�Xi{��p��~#6�q*��&?��k"-�'�g#�����T�-	r��穉P�9
o�@�S���;��XWc��o�V��D�t �����
�4
�9�>�f���z���h����# `+ٜ-#{$�JVo��Ȋ���u���rdfd+��蔽
9�8{���2���{>>�yEd}h
ߥ��lǆ�Ԉ�����b6�D=�1:��L�PЂ������J�OR�n�U��gU�u�q��ykœz�M��~������p�4W62/&R9��s�c�bd:���N#�Pj�̥���i�f˕9��;�%�6Z�??�ϭ���V�[ōދ�fa��͟�JF�t*�!׎�j��l.��wsE=����0�a3uė�p���M*.��Y��w�d���f���G�T%���a،N`K�0��2���5:rU�_݈�2�n�u�ܻl�Fȕ�6U����u4��6+�L��9�`2/?K�w8��👱/� ��T�8���R���[�T�x��9���g����M�ޫ�G.�R9�[��>��%���T[��rg&����M�tz�=Y.��vU1�Og���r�ȟ�_���aR��ȣ� GԞ�O���XO��#d�Y�jB�/'@�u�t��܇{�����&ȅ]|���(,�8�G�fO'��+ ��4[���EL�������vVT:����<;gC�r#�|�=\���\�!$�(g��Ul$CZtr��b�e���t���b��Z_�C�y�q�}=�j�қ�2�f{ѻm�C
=���fF�۹�h�.o�f�!���N��#�B�#�N��}�]7���g!�=7�����v�O�y(�'�sn�uy���6>�hb�0��B/�'�O��r�\�b��I~&�"����^a�\�`��#Q��sѴjK��9��d���if,�*anǵ�S"�0�-bQ���-Z-��jK>�����ͫ�%�aCV��j��F�����4�J���j3ߺ��qe�7�?5��k'�.B�����>�w��;����2S}, ]?M�2"~b����Nf����r�"6��G���)*K�c��lW6!���GE!KT�Ӵ���V�B�8��*`�bR�s�h����~1�m���DP�Pχ���Z�c�\ C�PK��d����9�q��r�©xo߀U��}��~�2�e�� ���8��(�������^>���NB�3�Q҆QL/�:��J��_Z�[Z?�֓sx(��%����1���.���Ag��9���2�aMݛw#l�
�hH��_��X3�0
�i��x���9�[a-�����o��)��iC΃o��X)�x���ڣ�u%ܣ��>��s�5��!�˙��w�6A��-_j.]��Ѻ���kZ��J!w��a�����άRփ��u��ȡT��ZQ��A;�����"� '$<��i�^�˗ٿ��DQP9�xD���)-��fk�Z
)�bH�M��|y��:���E?��E/��%�96�L&�G(�����#���d��t�51%:�q	Y�(��9� �I	��k�A�����{s)MbӐC����t�n2Z2{s�q=�)���<P��>�h!��[5��v�E;�!�����|�2r�s_�3�`K�ES�R�֢ђv���e��軏�� �g7��7'T��2��զ�Z��]�ܤu��ZKO�G0��{����ѨCN|�կ��i�s�)]Q<}Q3䊔�WY�>��M
�٥e�{�I$sT��
�����Ё͹��r�lm�2	�v�ӌV��y��M!����K�nqS����i�����7�g8�V:��;�xn�o�Bnĵ �l5eȶ�$�>��ziߩ9/��gJm����W�LE{9��
��tڦ�+�����7�~������9ٚ��K�j��F�ޤ1K?�8!n~�acO�A{;�>�?�	��:�^�B�fG���~����(�-�!lߑ៺�#+�0Z��>��\G���eѡ̃�;y�R)�4�BO �^��S���1�[O�q��k-�%�vŜ��ڇޑ��s�R3��!w���`O���ӯ"�>�w7�rX���t"驦M	Ꜵu�*�rO�&'�YurZl�-m5�r��~�1E�l���繘n#���J�9l�i;G�J�A�;�d�5' r-�ϼ���ڐ�-�'f)(
�!�+e~o�yܩ8�rS��b���p��m��]Y;���o?����r���̓�a<�򃔶�ǘ��I{p�4b�,M��Y.s�!.��JB�g{M�+�S�۔�-�_�ŭc�W ���c]+�[��6�Fa��Q� �E8
�3��
������^<����a�8Gq��0�A,�0��C�i,ɪ��j2���(����d9������C��\��S�5��ʻ�ǌ�ά��	n�-�\�=N[µ�X[T��a��_<�t^ab��f�x;ޚ��1�n�[h��jk��Z�w6Y+|�O���>��>�ыy�Tu¿��L~rJv���D$�Nƽ�o׌O=���v	څH�Tg����p�r���+��0���k�g<��G�ۈDk����7�<�mڎU�������d���˧����Y��!wP�t����b_e׏����AN�(mq��W����)!Y��s'�r�"e��v�U�VA�h��\Ƚ�/�$������P'aL��n��� �b�}T������	���$8�O">eo�Z_��2�W���U!�@��S�-E:mž�C.�럷e���*��ڐ�D��O��܀�_&�����:��$�d��Q���܌�����z�8���r�~�����4uR�7_�dM�q�b��*�2&��zsp.����3"�nC�����[��7�O�~0={!�d�Sё��AZ�e<p����&>�Q��E3Қ��!TZ]��)'!W�n����<lv��1
9�z��~Z���Sr�����.�9�[?l`�;���s�^��V����Sw��0O%���&W�& g&�g���۸
FNšD���v��l�>#�:,��u�M�ړ���R���lM�*�&;�'�Y3���c��~�6]n���)g*��r]�d���! ��#��Z��-Ƚ3{�d&���[��|D=��ID�*�Ҩ�>ֲ���nѨ�i�B��~���WIɫ��f�*i+.0�]������mZ�A����J��<�T�E����������*x2�0V�B���,   �  +B  `g  ��  ��  _�  ��  K�  �  � h���w<���q{������4��"#ɈlB	ed�薽7�ɞٕ���̬�������r�u�y���_���k�M�Bk�����mo�>f��i��eS{+$�G})0��;�G�|��3��ޭ��]Ֆ!�u{`�g��M8��蟠H���@��5���ٜ�����ݳ{�_=|�Wv^[]�Y'ac�m�xX2˝C{����.�s;�ش�&>�*/.�뇕���:c�5��v��L��W�5�8M8acQ�ӯ�\��0�C-N�{�%��%���t�h6�j�X�{MJ	���E�T��F�\��xwE?�_��˒W��>[L���S��DM��〱�8��n҆���z��6����0f-�UO|ڈ�yTᢍV������0V�F���72i�S��Lp?wd{�js�|�t�?W&��k�/�����ZU�pP�d�j�>��̙�R3J�+EP4��TjF���wы�X����(5|��q�\~~y�a�c�+J��tjm�RI����1�eQ�/�,3*)�_�n �-^懱��
s��9�k�e�cz��|Z��ā���y��\z�e�-O�Y���T0��3��u�qjf�l�;���i0V0sR��=�옼ץ�jc��S�I���ۆ#���d��7��M֭��4jOG����N^!Ϟ�1��״nil�bO����૴����ݰK�$���k���T=�U�Q�����h g�ܣK��٠cj�;Eo����dC&͖��*�"c�"�2m׋���I/ru]����Sb��V�o��ϞTH���S�cj��7�X�$��)-�a��%�:�]�)�����a;��U��lV�pk�1O~[lʝ�:�OE�*L<��j����ꓘ؁1��U[�����ˬ#��[��.}���Bi����6b^F�4)�Q��`����l��l�>��� �/:�#_a,�^�5��L��s��1�u��{c�X㫏'�:(x�\�4Q����`��~�3A@����n�qּ�'�>�h2�x¤����e%#[AS��9���U���íwj�M06���i���C{dOd2�ݭ�ƞ��ӊ��_���N�`�%W�5�)�]h�*X��m&�qV����c3�/�uu�4j$�#�~>UI#Ƃ1��𖳯ńl���R�.Ø��e,[�ώ���҂­�	��_a��k�H��G��>Eޓd_?��XH�G�}�R�43��^B��TQ~Q8�LI߳c�MX���`����41���ps�������7`L��%���6)������-A+�����j�Ы�34�W�w��T�c���1kl�$èm�s�Y�/�aL�b%.l :С����Đ!�k�0f�ܐ<�Q1����=�j����XV+�N�|���;_i�c�o'�}|�A�v���z����i+Fn�Xc�[d��L�ߕ8�Ƃ6���j����iF�l��*�RV�1�y:Z���vu`�<�c"֩����=H�D�bb&���>c��^����.�h���:����Bw�"�W����DpY�ma��1�Ko��(K������}�>�c��6\��dH ��������b�]�Hp�lߊ�RMx�-*[\�fc�D�P�
�&W���a��F�'j�`l�lh�^g�u8�qȘi�,�M��I��t�����	9c�v������|�h�=���s������0�0��X�A\I�Ep*��=�$�Us"?\Lm����c~l��";��F�x�(i�b���d�p��Xv7�=��ܩ�25�a�r(�u��}d��U*��Д
�KyZ'�*�K��^-��BŵrV}�=C~�����W2K��Ņv3`�^t�5���/L<�ogg���}�-MKX75����,��[/">�9~&�����J��>��ci��m��/�P�P��a�#��9t�]�lL�q�G��0v�u�}lt�|��[Y�`F�,�ؠ�,W���r��'��r��y�6����L�,]b,a��Χ���J��V���.o��O��!@���#��qv��F���e���EN�2!��ˌ{���x���r�Î5���HG�����z����#F�L$�1?m<{���UpI�w��/V�+0���_���.$ۺ��lt��Fȓ�� z^l�s��Z�$/�)��0�f��-3Y8��,>}'�p�������uG~u���޾��>e���T��+�ͦc��陣5v`LJɳOTA%Ὅ �Zg��z��Y��>������[��w�]��2��B;#��YCPj.�	d�<�a����
��:m*g���\tu��+��aO���y�������G�+��{�"5n��絪�*K��3�"Y��e����yL��d�Y�[N%=l���Q�J�e��߻x�t^�[��_е�$~����1R����ʽ�xqK	�c���;�/Sċ;�?,-�Q�#62�.�q�xN���	�h/�]\�F��r���!��������CSbTI�oe�'��Md��(�ѿ.�a4�@s��ғڗ��%�ha�Z�'x���泓jM��3Ȋ9�-�0����w��і�M�YB�`���H�y0���8���	:���@[=fc����o����籏u|x'��2�7��r_�vQ����BUr���%�c�d����%�,o�]��	cA1'b��"�rb'.��0�}�1Ƴec,f~���C|���<��`�T/>j����B�yn1�ޅ���0� ��4NN��@s�Z��`�c��?X��B�bXmw��F�|�̈�+o����f,���}�4�
s�\��G���1J�|>�%܏o�����|ư�&�^����\>�p�]�7��gb�|�X�9gl�6L�cg',V_�D>T�9sM5�E���'�q�r�Kms=��D���"<<�e�bņ��^왻n�YDf�aL̡���o��	!]��Wm�s�=y��uqf�V]�=��b��T,(3+�͹���n�(w0�3)p(ۂ�Ⱦ4���`��:a�/��/�%�u�p��j��6l��;t�6x1^�����fM�g����4����_S�`������U��hɪ%�ʭxӵ�c���U�u�O�rf�eFHW>���	����_&�(m�B~��i0��K���8��-o�E5��B63
�ؓA�>�M���H�k��v�ha�)(s Ͱ���������1#/*P�X���wԮ��}qh��t���njM��c�z�մ����\�������T_��aQ����Er��X"o%��6�p�$G�o�z,�0����KPQdl.R��t5���߬�ۏ�|�kOϮ��/�o	���z`��ŉ�oz����,�O��5=+`́�ϋ\;��I=�y�[�Iī�b!������g2d���3гr9���`�c��q��HcSc��R��M�Y+;�"O:V��rPM�R��N�/6��7
�:�'���D�ᜳeP���I��ݵ���>�l�T~JhP����G.�$dJòuv��M�0Ƌe���;�X�ah\ރ���1�0�|'JsMϝmB��j�Dap��Q�t��{F1��im�{~�+Nb��D�/��d�P�ҹ�=�����0� 8��D`�C�-��p���D	��֨��y�z��2�<�V
�wH����w��Qq�{Oj��x�l`��0��8+%A2�ۂ~�=��Ɛ�k�ͥI�2����i)��gTaL ���k��5�xVl�<ڢ �V��J)ǒ�N4>�A[�^a�V�=�D�J�A���~���s��.�����9��3�<��t��Ez̀Bhd�$�JC�m:�/U>��	*�J�3�\�5h�}AN��X�&cB?����U��k���˰��Wpy�KG�k.����+ډ�XK긳���l9ytQ����f���y��k���FS�k�<-9��9&_p�&���XMR5ad ��߅1WI���4�J�����Iei���������s8
r�����Qh�-J?`L�󵍠��v�6_��	���c+a�o%]��c#�U3�'�'`��C�u��t��ߡ�y�l����tB�?V��N�=�al\0� c��C�)y�l���p�R�1��/�������,�7l�{�,�csze�I�Q���rr��Qg��aL�:�!�6��'%�e���d{?ƪX�knkl�?�<�{�^z% �<<��4:ȩ�e�.'�/��C����ޠA���bꤻ�Y�z�a0F�p)�F���gs;��*4jo��B"��=I���w�B*�a�WdN/=�*����eJ(��I4���B1K0�6\̶*��c�H���Ů9�[+"C�\0Ə�t붛9sQ�/	w���"SwR�zS/���Gt�z� ����k�����혚E��lF�6�H`���= �,
�;`�M�6�l�ʜ�Y7�O�Đg� �	��>�<`f��{ X
0�2�p�/���r*��+]���%I��������i`E�8���	���67�%����CL7
؅��'�	�
��4����kv��U�|��\g�Y7���bI���:��;LX*�`��h�9C ��"٨���&�+1y���ݧ�̥�%# F�10{`1�X�� s�,ؚ��*�]۽k?�iƙ�P�=`��ȁy ��X02`����}���2�rp	 �
}����5�� ���n`F�ƀ9V��8�+2��5#P�d�j����[m<�DvX	�3� �vX06`�� �H{֣mi��z���6�i|G�`/�=���E`/�=���80�>����H��edIʸ�=�耝 �X�>`���Y�6 ��	�CL�d?�A�l�h�Ma���{`v�,��;�	�=0#`�葃�n�-s�f��N�m�$����VLX04`;����6���� խbٽ|	��'���H�y�lX��~�� Ur��D��I���!O����[V|d�=S3�C[�R=XZR��!��Z�sJ�s��I�X0��S��S�ƿ,�+�ݭu�%���d_�f�Wbö~��c볎�0�#��C���C�Υn�G�o}�C՝������o]�@~���Z�<�|�R��g!�̛.�������.ʏ��o������9�ɬ�yqD�B=����+;��~���`�0r[oLK��Y�ޫ
^=���>;fqd��L���;L`�nW���xJ�nk�qm&�������.Z�J`�VphzSлCR�^g�=�SE=o9*��2�=W��5n9y�{��l4R�𼮗r�¨"�˹\�����F�L�����;��(f�W\�b�XL����u�*��N��f����[Ceeě���
� j������LX�jc��It�B�,��O0�uj�xԊo����0npq��?����p`�ҁ��g�<�q|M�֐���]��<���cm�ȸ�=9���}w�玡�w�K,ͻ���m��C+����0;ZKoG���]�1M��r�A�~���.�zd��2�>̿-���Y��~�C�d�d��4��hQ��J�-�q�����A$G�S2�/�'��Y��e��f�9��L.��X�I͖��
W|�u��>Z~	�ڭ�h���e/��dǐ��a�j�1�*J%}}cFc���FR��Kρ���&pU2+q黃
]Q{�e��"��G�,���~u3dE�9����ՎB��ۢ��>VƔ����1���AǕ�l4�(|헙�m���ԗc�rj���������:�^`�+���ݑ�+&, �I�'Y{�n��.��*�6l�Ȧ�m�0"`�Gݢ�����v���=<�ď�'���C������f�q�����ŏ:Ǵ�udeK�E��X'��Eٞ?����x�g�l���]Q�1�}�(���9�`s�:�M;�}:�><J���f\D��-�O�q���z���V`-|�u���ǡ�;����PVHȠa�c�rEE��(F�ʖU*W��2#Y\�������<2M��4��@�I�:�6�f���;2��a�!���:�Ƣ����U~7�:�SM��k���P�K�[ͶO�k*N���zTWĢ�r��,���b�
s���$7�o�,5���CQ�ف�ˮ9���m;����PG��!#<��۴��b�E&ʀ�"��?�P����& ��U�~0ũ����,56��oh~3Q�Csv�1�CT��ZɛŽw$rIVq�N�e�q���{��щvϏu&��[=�R#˰�&�W�6z�>ao�tZ�k�l�"��?t���n�*��ՙ���$��`d�|w��CC;�%����������w�e!��E�"�b�c��9���L������2?J�*˲������-����>���9aK���3�#;���� c�, X<��`�r�[�@�^��l��h�Ȧ�-X �w���u&*S���5�g�r'Ɛ��@��+�7�
�]`I��x7�b��ߢ��\_R$8m��#�n]�\7�E���yT�틘�mM�ud!��p���(��}y"UP�E�!�@`���;���P⡉ ���7�PŲ��&��m�]qW��zΩb��f&����i`������̕[}7]
����Ϫ[�t�����2m�GI�w��:��?��h�m�w8V܀q{�2��ʈ����"�B�U�jB2�C�d���Ȍe�=�)�(y��s��:�����\�͒��Hv�ێn=����1J+�,`�``�`�`r`�����9c{�~�L���q�[�ۙpl�,�5�{�pG7g����h/�9���N3�NO�	������u��N��1��	9i՜a�1�����}���V��r��;}���i��a6f � ����TD�6�໓�Q�\.�`�`����������6��fٓ$��n�ofj;�Y͋�L�.j�`�DF�8)yR��R�HY�s��~�K��9�Ɠ"��3��S�ܰ��1_Ru���0�nl���̡+�`{�d�,�����9k��mrD��+��rv���Ϗ䝼���1fK�#�D����X�����~Ŷ�y$1at�|����"�R���~�s'Xx�U[�#j�H>c��#�N��R`��3^�Ӭ�o#F���1X+�X9�v�=X7)�I��H�勣�jt����^.�z������pb��=��w5�P�;�-�&��V�4`-� ���S���$�d�5b��ׯV���j{����+:E���؛��QO���3%̐Nl��n�Og�g?lh�q:�TM�%;V6
&6�ٲj��&�>��$�0�vs~��2�R�Tc�~��n��\�Q������"lOd�N_�������ٶ��`9[^�_k���-����4W[��"ؒ���B5�o��s<B����)^�;� V���qF��=���ui�b6�,��W1L1�K�m�䌖'2��3{B���ݢ;���}�ݥd{V�
�u�p��i����(���	�)%S�/�>��*L<[f%ikHI���3��;&v�l�lG���Ly�����@/�#�I�v� �*Q7��Cq[X�څ���	y#*�:�Q�FId��-�ߚ�vw�rR&}as�Q��EAr�cv<o0�5��(����r1���7m����O�iTN�.鄁y�����ŀ!�:f3c�5�m{��E��D6¯��۝|�k�	�.)��HY�&j�`�`,`e\V���#����Efx����_�]P4tV'����r� �<�OW���w�gj��z�g�&�T\G,���L������||�����%�����>H��� Ss�.A�fݖ���q�W�R��#�s�y��1�߁ɪ�\8��C�o�CFW>����\�jFF��J.a3.�����ʾ~j46��R7��l3����	�����
�xoɸV�v���;�e���n`V�Z�/�}��X�e6ʽ�A�U��<���D8�:�?`��Հ��̓]X�KQ7b�%�Qn�r�A��lЖ�m�GEh6*6�1�
]���`囬8s���B����ɦ� �I�!����&�X#X0������]S!���Cg����oᗱEL��9��D������nC/E��#>̶e'��-�5;�1�Q�v��;��Ϗ\i:����\���W���<��%�"k�ِ�T�J̶�m3[3s�:Ω{��%~�C����#�V�����m�\7v�e��|g�J>�"<�5���,հ�h4	��;�f�*;��80�aޝ{�!��*��Ǟ.�1���X)�0���8��l�2�ͫ/�̤�Ⳝ��[�����;��v3;I��.���u|����SL6��!��*��N|G��6�9�H='��K����^���	�.� �]}�1�P���.�ݣ�N�ZL|�#0�����^�׊T$�"=#d�~��
�lL���t���U&�ڗ��z��?b�Gdiŵ	�	jR����x_Jd�{��m��g±�ִ�w*����Cl/�]�u�����'|ܔ���)5j���l��;�6l�]V&G9��7�^g�YfHg	� � �V37��(���ּ����7�0�v5&�x�Nu�%��C<�?~z��Т�B�
�`3`�8�wFB&������|��SHڷyPQZ��,M�LC�vg0zO��af�9�������2��C�vR�v���������t��-�����ϯ�P����cI�m�]�Cm�q+���YԨ����:��^����{a�w��3��E����I��Ny����������K�~�r����'��Nn��6�UD,�l�X5X�Q'�d�Peq���	�[ן!u�k ��B5	��O��<�Y�碤��Zu�2�S��9�zp& V�t����;�����繤d^��'V|r-���y\�!tT�#W8��?���H������ނq�W��/���)�����ž����[�,@5	�%���X�!��W��VQ�����8A1�LG*��A���g��i�=�bQ]�F;���o���̘����&n�8�b�@0��s�g�8{`�l0����>�η=�f�O{v����ak�lPu����J�F������f�f�XĶ�ɂ��jf�!����Ձݺ�L~�Y�}lA`�5�lx	fS�ç���T~�Y�):)�c�ŝ���������M�a�s�%	��`v�,l�X��}Q��*2id�Q�\ٸ�;1큚�U�t�>\�خǳ�����6����h��#ݠ��R�t�������mb�5N5[EL��q��[�^��7����;��GSڢq}=9l�)�V13�3����"����6�u���{����N���ia���;`�`-`M2�ԚW9��˽��u�}/G��"s�G��	��8�t�'��uX=C��I�˭I���4W����a?3��X(kݯv�e����ҍ�%b�B�飍
�`B`3`6`��w�2�X��(G�8o�<��f_xɩ �j�``ls���D�������׸zފ��x�yx5�#F�6�����r}�`�M���u�g5�xk��\���][���e�R�9`�t�`f`*`�`)`�y���fKz).4wv����v'f$'Q � ���u���f��1���tj>�u�H���� �h����q��L���1��ɻm����Mt�D.G��oU�*�G%q�c��Yf�-L�̼Ͳ��f\���;�?�l�l�81ӮF-l����������
��a��M�,�!�i/~���,�Pc�L����
�*q}�V]QC��	4�_�P�_!�������YU�⺣��?��׸��&21OHX�<~�:b�``�`�`4`�`�D�����H��]�J����&�;���l��QC:�����]8[�:��M���t�ҕH�L:��M��q� ��t��J�/U�G��zu�e���;Wu꺱n���mV#U�?��Y3f`�`�`�`#,*�/��3��4�_�m��	���=먽{VƁuZ^��::|	Qw#�&gW��n�l�m�r�f��qF�d��G���8��b�^q|z�g^�)?i��kK6'�������?8��0T6u�1�9Z�����w�u��`�`?��]f���ȶ�!�����}&`,��)�C1J�m`
s!��D<��؇��2�n��3�[td{ƕ����1���h!ۣM0r�a�;z)����`Fi=�=���n�"��b���%b3�������c+ ��u���2���Ͳ}#{�z��yg�IP� �{���#u�;����7�|KN��rՋ��e�x2�Lg���a�:��a��;F���9��ګ/��;�5bg�����q��Ł���Z��e�Z�K��`K���������ʠ��	�fSa;Tq^�#e�����m�׺;"�mF�L�g�Je�R��u��P5eeƘ��������Q�i�����g��u�^�\�R9�%�L����z���*��`�`3`���!�곸N��?�I+�H��4||��Tu	L>�;�i��uJ�V4����7�/��o[��Y?w1K�ݘ�U\�
ip�E��e>����]�.���|S��N���_CZv�./�H1����c3�����9����˖�+=���zK��c��Z��*0o\���rS�~ŏ����bX�L�tHv�h� f �3|�X.�Wx��|r׎��El��/������m�'���1��/XM��0+;8Qx��E��_i�R�TL���`G���2�����5���پ��_r�5��VR�훷g��nl��Y�2j�`���?P=��o��)�K����uGt��+!X6�TJN�~��s�|x��Xp�m� ���2銵p6�������������u
�1ڒ���"=E33/��������FM3�=E�p��Hi{K���h�r���n"���qf��t>�P֊��̵��v�@Aٵ��y�Y?^?j�TC��J)�lY�gT�!�!X/�(Xn���'{��Q����j�^VL�S�ƅY3j�`�`�`cXS�ӧ���7����vC.d+kpG�l�9���=���6�7ϳ�0������C:fd;�p���`Hdh���L$�Ͷ�����O��41޴�t0U00:0|��Ge�m����È��;:H3%v��� 6���<���DF��Zس���j�fˆ*"�����
e>�����YR],�J0mU�峪;�OwE{�m�w�W'H"R�
o�ʣ@��q��`W����uW]b��%;��*N�u�8�l>w�j�`$`��|��_1�s�[}��S�ۚ(m�9��*�R< k3����t��R�cĘ�6^Р�ݶuy�����	��>������g8��l���#�S��Y.5˔�|�S���`�΀���c����<ؔ�K���7��"ZCX3I~���Y�Ԩ�
��p6�X��n�b-��,q{��!����N�6�<�'���O����S_ ���6���m��vt	��Dyꥁ�M���僭�G7 F��H��%?V��YP:�T�v���&j�Ud$R^'2��������b���B�-�=�;[{Vv9Nx�r;�^^��E%���~��\V���_��R��^p1n�YfH7��
vL���V7e�������K�OV���Y1[y���0Z�\�XW�RqP��So_�/�o>�Kp/C��v�����q��Z]���'���i*���Em��S١9��U3*ڞ�����
�
0��j_���}��/�\m�K����`$`�`[�L��N3a6���		�Z9y�J�[�N��s[bm7y%g����<��`b`��Y
�v�Y�B���L"�&��������ks#ݔ�Y�����Uxk�['��=*Oto0��]�-ߋXX9X<�XX�Q��C�%],�]�V��f���A�E�l�D��`>k�!�}�e��^83��r#=�#��a�� 2�o�8���tb�I��k���?-���yk��<��.|jwy���_3�3�%`�t�`5`�`��6�:L�����Fr��wy�|���f�n�]3�{�u�����+)�i��wO��|1����`q�	���I�бo��*�^U,�g+�{6�d�&ۦ��S����C:�/2`e��8K�"s>��-����{t_S�ԁ]����a��K�|ZF�|��� K�ཪ{�Ү�e��c���*�Fd��Pc�����P�!��$gmC�$���nx>ؕr�(��FY'��(���v�1Պ6_C�Ml��6�h��h�#v��``�`Z`��&�n`��ة�Oq/��N�v�Q�u_�,�-�3``��v�:�$��B��d�n|H���Fs��E�Kc���`��fq����\�mC�8r~�X�Ch��6��L���\A�t,�!��l+�'��a�t.`]���:2\��M��T2�ϫ�� {6��YsjC`F`�`��_E	�ntWeI���1�k��D�d�a�@�#8�]��yNS0}|�r���@���v�}��nX��(�0Y��濐��T��M��$e)��n��Z�<���L���u�������f��<��;b�����ˇ�y������;S��"AdȻ�ֱQ�K�� ��p��lJ�y+bM`'1�J��E�x�`��$)U�*��k�{[�+B�B��V�:F�cMOD��lf�`�`�`�`�`#`q��ΑUX�������{��� �D�����MԱ{o7 ����љ>xm����f�;j`�`8�w=	�55�~q7,��r��:���,���.�̿���h��?��<fC�a�׾�*������ݞ�6�L,	�0c���8�Fw�����>�@nz#-�m[W�6�>���"2_3�����!�������CB�Wm�s��X:����Iߕ�L�%�醠��������7�ܜ�vB��]�:,��� �����Q�mi�@�qM0AR�υ�U�kt[�4X2�� j٘	T�S�j��/+g����?on�S�"��7`�`H���a�+M�'&��C͡z�쾭//�w�M
ʍ'�՛�L��\�����!]6X;�X�g&���X���{Ͼ��K�� {։Y�3�*�:�t�r�.��~aS��5���4J��؟����03"#t�~�f�^����=�пj�ۙ�S��Cj��]�m�;i�0C�$a�6J0c1[:��HJ�4�d��|��Ɇ�G�� �k �w	�UTR*������ے���_��rC���9��X,�܏3��_��y��v��75���vK"��1�s`�`&E����"�������D&�g�D��c��O~8|^��|Yb�0k�S �v,���>-�bd���w[���8�Y:� ͟�̀���9u��A���]0�Jc#|�$u��a�R�7���(�~��q.t�D�QD�]���c�R9���ɺ>|��I�b�޶9�K�`=�q��Y	�0c��;8w����t����[�z��8z�`4`�`<��������O����ˠ�^����\1��\8�RF�����'�VNd~�;��!�/f�}�eb�`����i�|�l�,:�c`��`k%��a�r�C�����[�J�x���
vL��?��`�\6�I�������N��iǖ�Y)���C��=�!���/%ß�TY�S�J���q�5���Ӽ��k���`��,��rC�yP���W	�z�R�V��XM�W�0:�]����v�m�;ƖS��9���.�eS��-:U�T��
v ���C��U���̬�V�_s���~FW���Pc ;vg���{��b��P�~*/�;��%+iz���o��U2��+��?��Y7f�i��5�S�u�r����{��m���tQ���@M���w��ؒ3:C���X��8���;b+��55�i0�-(�/����Ry"��t��HjRhp�X��%^�-�|� �s_\���>��r:I.�3��1�:�HG�L��,L����$e:]}�/í�V�2���#fw��������P�Ĭ<���g}���[<Ȧ6y&Ǣ���_��'����!�se�{jn�}i7�w���]��fzT��_�G�*��q��g'q�ҵ�}��R��?��l+���'Y-��V��`$`f�	�Fvl ��|u6_��4n4���� ���`>5�������!uj�OP����}!��Е�x*5�c��b���.<���^�-l*U=-������~�|h��w�q��N00|���C%���v�6r_�F5���z�oB�2f����DV��A0���k,�S-ê��d���:`���K���Ɇ���Կ�<��v�׵R}��ު(�_�S=�!�X2fw�l�����f��b]��Pk���Y��i�U�YSτ��G-,	��.�C,;�L�fM�*��%���t�8��c�(X
X��]�P�Ǽ��S؝�qJ�t5����+���!&��թ�&�*Whp�3�S{9��}�r��n����;~���3�K��,1�(0	�@��ƍL���H�T�?̎�\�=����P�� ��3��)�c��=/ڟ��Mז�$}~��OGm?7k�߉�j��w �I�i��&���M��՟q.�e;��0=0F�0��趁�x�ˌS9�I�;"l��aFҶ4��K5K̮���t���Lr���)eȾ|2�̾P+���``�`�Jk�Dz[��T�7��SY�5LF��������ؚf)��[�=��8{���k{�,�35��W������:UV��s���0�F-���י�-ky^�/����c�[4Lh}�z��*j�`D���ݖE�K�[+ۚ�1�
LX_���G#�4Y3�	�ˋ�`��t8��,"�NSp�D��Ǐ}Sb�ϩ'4K�
���:�
����q.�B��ϑ68ru�l�Xa�D�����i0��a"��Z?�0-0�s�;M���d��Դ09�&m�\B/���/��ڥ5�/Cקϋ������;w�XQ�-�,��C���wv#6v L��3|�#`�(�8n�q���Lꮯ�k��`R``Ir��`�v���(������s�0��u֌w�?M�lg�`�`H�r�X"[�CK�����sRȺ�q�|�!��N�s��ӊ4��O��c�t`}`��NWSE������|͢.��8�ϥ5K�2�V̊�Q+kSKǺ(˟/���n�t�m|ԥ�8C0n�^�-����	T��!W���=k�i~[�{uT��1g�!J�A��?fH��>����!Q����۸�T���N����L��߭c�F+J��$��L*uc&�i�
gp/I]b�1+��<Hd�VP��Y~w]�Z2�pȇSҞ�������Q�)}���teS�v�-����`�F������3Jߍst�[8j5?!Ǝ�y��`�`G�����b]�Q�d���1_�c��4˄Zf�`�NL�>�	y����RZ
��߸q�̓r)��X>�u��G�'�^XJ؂X,㹵�̱�����͒ό�AL���߯W��=�0�{V"Z�W���[7�Q%ߊo�jݱO�"�z���&0��B-l�!؇�&s2Ǻ�[%��g��PT{;��U7�J�N��j���m�	��K%<�����`�K�nZ��qǐ�ױ�X��Q�ʸ�w������-��}�	�%k������6�.�G��}��g4��0y�B�҄��g}�`�Q��Ycc�'"C�澊��w�>���?��3>��"w
1n0I0o����3O�*�	��S9_�]Y��p�����ۺw��˪��G�r�lf�`�`����Ƀ��)_��S�� s���܅�����1�bC-�������gy��}�|�yo�7l���Z��&�vg����4��c��e)�J���Z�֔%e���Ebfx��J�����L��c?j�S�����o(%�5� v��.�ia����`_�<�s���I.������f��}`�w���%j���a<l��f%/w��Z��W����-])W�*y�l�_���t۸�q](�RʴGr�G��k��	[���=���X.�6�3%�X0�4Q��.�c��w=%k�t�Ч������������t�`}-�d8�q�3�qӈ鏺�]� ^�v7go���"�n��,��ƌ�X�k���UA����"��ڸ������H2�yv�HgƘi�I�1�т���5�q� )n3�5�xC�"� Ɓ�]9Ԙ�8����b]nw�Y����*�$mop�/ ��!���D��qF���y<����?��-�j�q���`��GoR��is�A�!������]8{���O���7w�2�����t��`��������!�^�+��%2]��<Gr`��񝥻��~u����|��G���50օe�G��9Q�4�\��L��w�j��*ړ�	V��X�����QI�b��������:�奡�-��q2��k���L,��^���__�쿖0�턤��#�6���@�_�q�9����u��O�"�Y��~��O����%o䰣s/�:X7��]����[����.�Xh���w<֋߀q�B��]��d�M��Ȉ�DE"�2
E6��g�&#+;3�Y�eD��x>���s�y�Ͽ��uձ��%k��k�0!��X�>��E�,E�_���B�1�B�=kc�����C�)�=�bj���%��
0�'�%����1�4X������߄X�
Xs&%�
�f<1h����ʇ�͇��x��������q�4^.27�oZ1F�>�QWb�;�e`?����
Y*q���w����2���&6����i�U�����U���e������ģ�بa��}�����q�Ӗ0QK���E���N�����%����}�i��}j���Э�b�{r]�6�Z�?)��~�-��%!��������.���{1rN��Bq2u	�ự�ˈ9<C�"/�<F�2'���ph��[8���z=�� �&�a����U�a���đgҋ	V֟^ţ�I��_޴����{�l�C0lb���	���i����J?I����&Fv��F��m5`�4�#�������[�>t�G�ECj�m6d�60m0O��/Y՚\D�o�N�.��.[v#��u�۴��d���S������Vf�*�Ku`�$���.���
�<����|#�|�j7G~�g�M�����L��K���ܸ����3���
�gT�;ݛ�����Vs@�O���^���T��RKe��VH~�IX��8�Q�|�6��^�ƅ3��Ť��g(�~�D��Y
8��}���gK������s[mp\��R��|8�O��Y��,��9��w��,�s%����>W�S��yR�����ze��M-K�eN
�g��;HO
��F	�܅�e���:6,�؇j��2-�`�)}���b���?����6���M�iK3-zҴq�2��J{�T�w�RO[:�	0b��������0�fZ|�W�t�WKEMY��͸�ޚ�Eh�.���F�.)X�_��QV K��N(�kq�JOe�YN����?ڜ��°^0.0�7ml�G
BT���B�N2b�&�a��10J�|����S�M�/5{����	m�_
8�
��&!�&�a�``+�c�K0.����[z}Q����>��h��;f�x���Cwf`?�/�ߨn�T�Q��xz:���$���!�Z#����%���R�y��׌�(��0������W�``�;�� ��#K3�y���e�)����j"���߉���'+�����`:F���W�(�r$���AӂŻ���x�~ĸ�<�
X�T��傉{�M��x��ԣ�����A�NXNl��pO���=V�Z��f�t�st�7���W��	�V�tO�$�#[~ZU��,�G ڰ#)<P�Z�G��^ˮ�D���P+N�uC���|�Yֶn�3�3�D��Ͻu7ip�Rz�{��L��
��"�
��a�m��㌓%Cω3��?�,ن�a�k݊��[�� �5�KV�"���WE��'�fz��d.q�d����m
���icXV��d����������c�1}�E[�������l l�_��6<r�bH��ߣ�+��w;���(�����0~0=�C�H2��O�*�K�����Dː��Qg'�q�q�̀at+6��[)���;��b�:���,O^*��V�BL�6�9��3�yŘ�aa8o���ֲ����K�Q�6��6.�`�`�����j�n l��g�|����r�t?>��O�-?#. ��0y�|0�{8�O�a�1&�>��������}e/�3ElL�|��{���zi��m�c�v�T��D@Z�֞�-+A�L�������ou���T[���u���by~"b`��w�(�;,�=`�^��hI�s���;�uQ����wO��*Z�DLl��V'����,<:G�J�Q���u�){^�G��£�`k彼s``n`9`�[���g�/*�m9�K����O^��	��&�mv�&�t�$��e�RE�9��i��4{.�k``|`Y`v�mv3���\�=�<V7{Oۗ�P1�׌Rn7F�?�0���h4�}���B�F�T��,N��J��`2�19���m�6�p�cL�~���Z���C�#�﫜�L.�a�|����a&��'���=�3�-�'k�uۙ�k �&��d�"6̰R�b����X�ޞ�}}�^Q*��i�B�1�,1O�"7�z�.����m�v���M��HK�W�=�����#VPp�y��^ocb;�`��E/����m��5�|��t�����=�6}�4Y�z������T���޴�m� �1˗�[��'�1�յ95���[�C������`!��#��t{�����Q/Ӥ,���G�);���-�cC�MΛ�&Kknf7�z�e̩�N�e��h�E��&�r0�GE#�Z�n?�+X��MԒ�W���ʦ���v�����9��Zb0=0)�+`�l[�,����L�S�(e���!��g�������
���fW�l.i'{5a�_�5]�{U3:�:�i�ޕ�n�#u�	�����Bz�J���hs,�韐���v�ږmvJv�H�,v_t�s���qfa�������`��,�C''�	0���*�_����c�XO��s��Wa��e�e��n+�N74�@�|KKo��<eDj�a��"�V�����y����o�v�������Oު�C�n��6�vsݥ#�FG2%�^*R@R�!h?�Ja֭����[e���l���+]�DGi5���M�l���$K.2�=t1���J�4���v��@L���$�;>A��X�*\�8�~=CkJ�<��a���`8`�`%`D��:���_``6�7�ID$d����k�Q��|Ք3��l�x05��˨�bi$�"�RbFG+־9���#`��*�]�2X�X/X$�sb���;X��mJ�T5���]��I�� ��O�T�^�HՀ�!fv�u\�ya����͹�\OrΉ�K�������\0b0n�B_��S`�`����ġc��;�`��VZ���ٰ6�����5�6�]�4���@�y��FGg�9+�����(+���|��0:lRl��
L,l	�Lm��g�f쫩��r=\А�K棥��6#�8;���H���Ɂ��t�D��e���>�mu��x�AG&�[�a00�t��!vgÆ�F\�o�{�G���I|l�Q�N@b��^���꾀	�i��p�h��di��C�F�)�n=�|I�eX8�p;ڮ �
6��� �m
|B�FZ���(��\���^�)�:O�2J�ރ��vt����j��e�ŦDi�r�#e�5;��u"v�b_���΀������=V���I�-/`��>���Jn��"� vh[w� �ͳ<9�M��[ �gT�v�pȥyĨ�"�S�s���Dۻ��{qH_����N��U1�m�`�`�`s?���7�nLdo���Q=%2Q���/=vYG��R��F���/�� z\�5#��h�}�u�t�U�z:�n�����q�Z�����#Fg��X���V����|�����W�㿯u��s��.�h{
f�o��`������9]���9Z��^��F�`���<'�`�'`��Gp������݀,��IO�=�5G������b
ak�=#���L �b���_���b�e���e'tp���B����m��.c�3#;
���u��$o�o�o�[�=Q��q�J�b3
L޸����1T��	�Ƽ��'(n+{s�&8�	ã� n�"�`]``�`uR/EV��������P�%bΌ�so�I�?:�?B��m9��Ő��4Tg��Ƒ�R���)���� ��WL+C7�b\j��������`0f�L�P臨�/�g���gݭ����F�r[֦�ŁI�}�G,�ˬC_���{���UK��
}���:P�C�'����#VV v	���&N7�C�k��%���_dV�*�
DY;X)��0�1��Py��:^唿��G�;n�l��~!R�r�� F��f��%m���X2��Qg}��;O�&��C�7�m�<�P]�kt�>��Iov����麪�e�˯�;�`-���M�倭
�l�/����\��y\�b��'�皪�w���Dl�?�� �v2`X�}nxP.��Z]W�^��o(�v,̢�Q�4�����)ܺT!4mK/���Ɏ2�N���}mv�<�#`��h��4�F���Kܪ��*}LC��=�)�I~+��v`�}i�����3p��y{1�od���Ds󜁃9��J(/�3XX�E�y v�����"���<��)�5�O����vK��B��
b]ۺ�`c���	7����r�2��7�G���,L��m���0KF�2��f�)�{��ӥ���i���LbZ�;	�P��^q�3��4^-O�P�d�S�a���F[!b.`+�G��-�S/��R�]ꖾ���m	����V&�օ�y�\�"�b*�_��*覻y���V��16���̀���
#8����
۱{kß{y��Q�4k��`�`4`���j�����(�s�V�}��T�x�����X8X#bw���"��{����Z��f��2�i���ǃj�-h;��l�e�{R��V�vѴ6f	�U�����I��^�$����F�X�$����U�P&�a�������|���x44"��ȉ�<�	f��4�x �3{� V�O92[q��ջ�E-��%�!��[S�G�c��FLp��Q�����F������Z�� �����k	��������ި�m���l�F�;O�)�}�{6"�H��&u;�6�����;������d�/:[��j������`db�����= �<��K�����d5�&��\
�W�&=t��L̮��FB���!vj[��G�����U�{�X��q�������s��``�`��[&��g�.ax+eU�T!~�A���*"���/���W95��Vw����mb�5_��=w���M�=M�yu���1��L�Ӥ��0���T��<�-�u����ʤ�֣�ςi�`+`�`�u����V��>�=<k��~�;�B�ݛ����Fƈa#`�`95�Z�q7,���yIRRF�S���
�C`>`~`�0:
T��[e�c���Xy���3Ҥao&Жv�Ò�΀I�1Ԣ�ڶܭ�8r�ϯ�uj�@GxD��8������Q�ouw���R��-�WM	3��l9�H�d'"�w��,1z0a0c���羂���d�����:9��]T��d�/��L�A;�:Xb�`����S`����[r��c����J.�W* �t|׬�e��(��e���1�e�{^�kJ��J���a�g=�B�s�(>/�A,�zhvN�"��[	ٴ�� u����#:�ot8rG��W�� +˙�n�°�?:�2)�E���ՙK��k�De~`a�N�`j`�`�`�>[��+��W6��師��Z�<m#]���"^�l�1�E���y�]��el�����Ho���x��c�
=�=��'���-sS�0�q庴2w&b�/��oE˩�U0L��ce�]3�=���:���^ϱ�试�,�,���K�� vL��O�Ɗa(����F>o�^����K�[�ڌ�>�,kEL�"�*X�_]U䔯s��ѾE��t�E�Iec�nN�i6`6Ff6SL�����R��V��|�T�����Wq��#�����DP]1�cɵ*OM��1�t��_���L
�=�y�I��=��f_�b��{������fn!�'h�#s[}��M-ou��.�Úi���\��O�c���hu�������n��]��æ��x�=ܴ־�G�h?#f��?ݴ�l1�ك[��?�J	�͖�.va$��JLޑ|��ǟF��+��m�{���ʿ��p��C�x�u����#��"�v��R��x�[m��ǎC7'��Chy����nQ���3}̜�%L#���z+ll)o
i(5�ѡ��Y4g��bPh�ςIB{5���������Eߋ�{�lF|��wd�UV1�!�]�y����qs�Uߥ��ه:�\�5$�$�E�*u�5�E��*Q'�����&��3h:��s\ "�ԋ)�S��Ջ�u��xl�����]ԣϙ���Y
7���p(�CK��ltDSB���й�w�����-��P����-
8���F}cӘ>V7V�
��X?X7��ڃd�*�Z�N\)	�����a�{�
DE8���o���%y̏ؖ�i!�r�L�w�߰�<��E�ݔG<���՞�e�'K]~~�ʞ�1­Y�at�ĵ��� ��6�X!�d�7�i������%��5(�vb^q����3\���6��x�rO��ٽA,ﴀ�']��m9Ջk��t�dG�|w[X���l,l
�;`�`��N��\����=,����tm[�	O��W,��IJrR������1�q��N����{����|�����ɉ�Y�ń�JO��ԕ�������I�~�j��r�k��qo$���?������y^��G?��S`:������G_P��X(<����m-�-�z>�������bhSB:ݼ憨V����K���O�Z���e0Q0N���T�̥y�0�R�!]��ªq#W���x�gS�I��,�6K���ј+\mv�]Ồ%�Ɖ�ı�$/�c�=:��7s�ɏ ;��s9��GW���͇���?棿���4����R�^k��|�G��U���U^�2\������v�Gϲ��I���GYU�ڙ�0����`t��b����'Jxs0r&V:g5+��K���wHG�HEL�z���!]ffZ\�N8˷�U@ ��"!��Z��ϸԛa�]�W(ǏU��:������v?�3]�[V���KvyYb_k	v���at�6��A� ��G�0���OH���N,�gu��b��Au]J�N��e�����m��hu"���s'�|�$�u�[�J�'ث�!Ƈ_��5����!����{`��]͟bp��߭�ZYl�3kf��W�Fz�3c��j2��)��}-X���i��I��`���pħ۬��q����-H�h��>�H�)�.O�0�1�b�"����n�y0�U�$�W���^tO�MG�N씋�zG�t�nJ�j����>m��͎1�}���{]~,>|mE�˭\�P���������,�р��1 �������̱�*�|M�R͔�|���Wgt�K��|����|�	,+R�z�d�r��I(��TƐ�H%�5��B���gr7鮃с�M��y�˯h5�����|��+�x?	���Q0"�ֶuo���Z�2W�s�\�_���1db'V�'�+^��$�Ļ�������&�Ԅ�Ի_�į���*��p���%#�Y�X$���罉��n�8���1����oR����:��9�րt�<���{"��$z?���DD��Y}��.q*��ߵ��*�9����g�M���,ZClj۾����羛%qQ3��(,��`���h�ʐέAi�q�XQ�O���v�XfD ��m�O�>���}]g����xiV攏���ͬ��R�d���%����;<$&Ct�$�t)�:�wڀF:%��1�U��S.�}�,�����b�+�դ�SG�[Jk1����hr�M84���k��������OU�%�%�)��;4��GodS�X>����l<�p+�WO2�����^*���Ʒ��LĔ���R�?G%���鑉�E�j0J��<XXr*ujFg��);w���i�u��O������k�+#d�"�9���g��=�Dۍe���D��J]m?)ɗ�u�|��k.���M`X`��N�������)�уa#�&	����>��6��ۊ$�G&wèV?��ƕߩ*I�Yry�˔{���#ϕ�?��yWFu�0�c��Ur��I�oء(vr��ao����Q*d}g�,{0A��ೝ؉7�Ï�LU���6̔��s�&�w�ީ�|������+P�8��YfB�e�}̀X� �#X6b?���N��>P.�'�u�-�Zo�SK��K�k�i�/��	f`� 1��|U޴;l��m�.����ӣ�F�������IF��'}����s{��&cC���O+�	!�
�x�mv��j#�e�0�QƱ��L������ջ�z�j�3�m��:���#�����e��h�,kYX�Xk�������n�h��U'��~2{O¹����(�f6
��½~*�k��t_WT��4Y,�?������U����w�����0^$O%�{�������R��Y�a.���D����wN`��77y1O2��j��e��3B'g������g��e����r��͍O�*�FcO�V��, ��-OeC�+�-�nl� Y��t��.�H�{ͯ)�v���89� ��4��n�U���]5ߣ���G�;�	��1�����:����V���W��[H�NKX��-eeZ�´��\u���2��jz3?	b�u�Į���i\��_��Nf;��ܩ��,��n��=s�<��J�u&�}^��b�Q�؉ѐ咆8j�5�b��Օ_�|�6��+<4����5��5�/�W-N�NLaF�*�#���h��v���7�;�{���a�yR��6�;,Sb��u�5�B��1���]�};�W��~��v����)�Ҳ9���;�w��ao���6��� ����X����)u�nVH�񼆯�ɊwbBg�;+�.�.��Lm�O|��՗�g�*$�1�r����b?����e}y���K	ޭ����8x�;��
���_�t��[��m>Y*AȳK��#�Mo'P^�@3.6�V�D������UiY��y�W�s�U�N�ԏK�����J�p�]ڵ+>��;1#��:���~�Y������ٷ;�LFh(�$�U�9F�R��U��<��ᬚ�tG��-�Β]��-؉M�O(��d_�0}l�8�,�k�p'FtW�u2	��]M*ץ���I"�߉��N^Te"TВ=��{��n'���n����ѹ����)�W��������ģ|#���(�yr�LRމɯH}�Js/�&�(�b�ɩ��c'�o@$FwS~�i���/�C��D;�Ja)�eϳ?���K�u8;b'v�a�=�9E����E,秲� �᝘x�����oaWM3���ic�[�vb�v�,8�c�?ƨ����4�\ى��i#'�\vt���7�/��I4f'�ok\-�'��i�届�#6�;���S��|��,(�꼋~��م�;�g�y�n�9oI柗b�����?w�=\h���eXh�@Q�$�;D�[A�C�4R*�t7�*�����- ���]W'��3:��w={{��QێA�u!cq9l.n�@��7��?��~z���ATo�Pb��٨�Z7�.�g�Zla�U7C�A,��ύ��{���'�%d��p8�����(�e�٨2y���>�/g�X<������gw�K
Y]�x;@L��/�sbf�m�&8�֣� �T�'w������E�hO/,=�l�jc2z�s�SrDWH'��bW=@Z]�����R����}fj�� �!3�1ѷ���,'y�KbG�o�����x05�ix��A�'T�Ֆ�?#KB�<9��ߙ���a���Å�sW�Yc��fbf�;��;��� ӷM����4��J��̘˗5&�,!M�"O��:s��]���E/J��>ВZN-�q\w���q(�l��C~��u�7Q��%t���X�I����A�nު��q���BP�'��I����	~���ꯌ�Ib�Hg�l(LbnzZx���F�%��9T?概�KC��6�",*a@L�uCuH��Ň���%ϥ����1�_�C{S�/��ء��^�Z���)j�`q�S� ��q�l��(IB,o�I��3�	H���f�J�>!���}�; V wUg�Lw��C�����8�bPC�4w�� ��U8u�� �X���.��O�_���Uq�cQ6�uc���P��efz�F����yc.rO�.�_a�h�J�s�e7���/� P�.'�.jj�X
�������C�/u?��G�.�mQ�1y�a�'����������A��*] P��d���́�o]u��� �?�iԴ���i�
�Wc�cW�h��"q�)0ք�'v�2����5b��������Ք7#�r��;�mF�O�^�j���^=�� ə��k�S���A�s�A$����jӤ�?���գ�u)��`e�Xa7�w���b��".X
�WA�AA5[p����@4s���~*q�/�aj�2�B���ޥ�B���Q_4����g��߼,u �w����=��j��2f{�~��7���-��_�93��=y�zwQ����ѯ����f}-#|8�J���?���~���`�3
�9��d��{UcՂG��y�ױ�`/{�c�f�����F;I4����>���g���ش-3v��]�ۣ��^G�9���;C�ɁJ�����׶�ߢf��4��ߍ�3�,�eNҸE~5�(�ʁ?�J3
w�1y{�EM.��c�n��ݳ��T� q$$���Q:�eB��s��+;��u9��%,�G���9��9��%�#_�\��)�R"T��@+Yݖ�Gva��%�h���)�a?�������l�ۍ!%.���/��w��/����o�Y��e�n�Ȓ 1�OӪ�ݪ�f���b1U��jv�_��רG�9';xg����6J��[�­z5�LEEze��s�Վ���ܮ
tq~4\�oo�³/�9����Q\�B�n��2c(����K��~����H��J(�n�_�����׏��*�ӄƥ�;d���+������*��N���x;��X'�-�=���O��1���;�5�<!�d��Z�WK�^�5M�FӸ�[s59�s�a��M����u�|�RW�o���]3>F���鍄L�M~H��7K�e�+����o�U�B�UW���4��<{o��J�)b�P�5��xa!�)2#�^��߆��E$���n���m�s�־�Q��iu���5��oo⋁0I���Gq4�R����0�,�<�"�DG�u��Mӻs�K?���;O2�ě��c��������f��,���J��K�T��^_.*��i���O��8F��/e�ϊ��͈����t�`�S�iE�n�|��x$����}�񵍳���~f��6'����w��h>$=y������>��X*�̖�=�bF���3s5�A-�G���%��L�Ű�����*A Ǜ�7�0����]U-��0��eu�z�bz�?��-}{�����M�m�Ԣ߲~B���=x�n��1���w����<��|s�M�kK+�/L��N:�2�ZG����J�a|��|��|$�)w�7���#�Q=�?3�j�͚'7���)�w�C�B�˿�r��7�q��ηh�b�s����0J��@g�l<BtZ9�&�Tdz������yx��l^B��c:���o�-`�MO"��)7�""������gV�5�~6���ѐo���~
��N5�6�}��ڣ͖+j{��hl�+�-l%X��>������0��߻1�k�Ӵx�k�TA��1���4�6�R?�1^��bA����\ܳ�F"r�ZM�kc�#]��yI7F"�s�~�ƍ˻!F:	,���?��s�e�	w�ݴ.��y�w�
�e_M�+��<���"7`0�~�)m*���m���ҵ�t�
$�
gw�`z�~���idw|��r�D=��>�����fô����G�$:lu�������{��e��Y�XG#�˙7�ԅ�S'�(����{w��I=}o���ı?7�v�3ED���=-�>|�V�?� q�x�7��#!���� .���:��ż_zI*|�)ҵl��7���y�P����P���R��^vS�y�L�t�˙�"G�;f�<2�����W��@Q�����Éю��M�cĒ�k�v�υ�s/{�*�V��7�'�D�/n��ī	E?\amϩ9����/�\�:yNc7�L�Y޳-�4j�ûb�d=0�zR���R?~s��;��CK���w;�%����LyD:'�m4bzZa���Y�}`q�ㆮ�/�c_+,�v��ej|V��T;�ׄ�C�V���iG	y#����7 <l���+���t�)��Z������YH�-1�+7��(gs�¨
?�ub�eW(;���x�۵�x~�F��W�w\��oK
X]�V���X����~<����Ix�pPTn��`έ��9���#𖥳�Q-��fԡ@t��kk�2!�p�"~+2�G�����W�u����آ��.=Q�*���
�4��Μ}���Bl�iU�kxi�������l�#a��d:II��ۿ����,w�-�M\���I56M��|sՏ]:6�j��a�#Ow�I�c��>.�ԏ�#�{��&��°��͠P���,{�A#���a�<z柎�}�Y��6K�Մ���ԧ���;0wpB�q���!'D;�Z�̿S��`��ES�~@V1�ݫ7'��]�ɆjTjV��_�a�E`ײ8���aP�RH��?����X���$�;�G��и��0��.��,>ZE\f{�D[��U���[�6�5�j\�\��MV���3��8s���D���Ԕe�F3%D����w�w�o���V���d�����K#-.����ʐ�rk�~�:���\�O���y���B�{'{4+NM��
R�D	�۫ѹ�Nywh��H�ϱ���翍���qB��c`���]�+c��͇��-�YͬT"-���;�Ҭ�1��-�Z^�V(�V\��|�b��|��tQ'�sK�?M��Ռ���M2պ���B��F:�{�a@�JK��+�-�+��^�D�U�6���6��%���xZ��+i�����d¤����C���q�%��'��~�����&����1�&%����B؎�85�w�� �]�-8_����&�8C�������ꞻF��}����~�������"��7��AfC�RP����zZ=��.�7;��~�!|[�g�"��KO;��� Z�9��Qm�H�����Lp����h�����O�:���U�l�T7������{�>5�-�1K�� ��z��� ��*�g@gQ�{����1rKҏ��O�6~7���[��w��!�&ʡ}�NA,i�[ٛA%a ƽ�����s�u�Vb�.F��lɞ�Q�{v�������Lu>IQ�f��kq"�1��pM���r�Q6d�7{c��_{���J�_�տ�g�E2Yn=���9gv{GAK��~���nZ�ZA�>Y�@��Z粭_��|����2/�W�Ċ��/F�-E(�{�?N�ZnK�����)�d�WJ�Rm���| &�!�*��`��ݕ�+x��>�(%n��)�"dh�+��:���ԑ��%�����&� �]"K7�Z`�����[,�Y?��,�N�%&s2Y�G=�Ҙ�Tb7��R}X��o��Dk�-�UE�XyS�h ?�!�=��'�Vg�E莉jE�+ݾ<���~�<���
b�0V����|��u����&� 6��V�B1_u~�N�hq��$�q䇄G���3�X�3�*�ȁX���T��j)zT:_���y���/�2�8��艬��ʐM�g�1�!}�$�fs>�H�s��[к�k�x(P�y����P}�ΦPT�ͭHvmN�LO��\[f@,�l�hIe 7B����4!Q�5�E��j�*z�.��e���.�p�?�+)��+�g�:�G�R��g �}fN#9	�TS8I{�4uN�İ��h=��u�2��%{�2>�br&ޭ�O^/�Y�K���c�@���������[^�%L�6~��T ƶ��M9:�v�vu���}�.˙,���?5`���y��̦��	b.�|#J�(���E�W��HrR �����ډ>_��6���*����§���^\�L��j������ToߛU�>�h;U��FlJ�>���>��T��)!�K.$K����R�N�X�]��s7Vu�g F}��<K���UC���dѥ�1���Y��}!��P��_Ԫ�6"P1q��.�e�G�~��dT^��4���X�@9�s8��h�IAK�r��?�u�輑�����~�,�w:bL�ڛ�fo;B��f�=*t��@�i��Kn��d�Z�=���.�22�	|�"Ū\�����t?��ظ�{������x� VhZw;#��,��V�/�����r�^�Fb�g�k��4��\�D�#t�
��~/�gw�N��l�GU+S�uk;�I�=g�m����bb�A��
��L�p�4���&[@lVrR�����t�J��{�N,k� VyN�,Kl�-�=� �#�s_b2s�Yӭ�Ўn\����z% ��u�� �%G{2�	�2�$	Ħ	#�ߛ�}¸�ږu`�}_�Ĭk_��'J�D5����(���1O�{�Wa�.��`�uQ��X���L�����S��W�u/aP@,W�6[�"s�;���!.L8O$�5W�kQ�G�W���e
���8�����]xT����KOA����}�cfa.o�5p��i/�Ģ9����"�J�6���L��=A,<���L���]�K����&�� s�@+J6�l����NK�'���6.Z�^����8�j�z_�"�|�ػ,<�Ϭ�ma3,
�	�?���&��D���ʥ�[�Hy�;��ȅ��U;�����'[�^b��I�>tAG�O� F�B�3��F�u�����ֱ���EJV�ŶU�m��d.3z��K�b�Z��$����ZN��m����竧�n�q�f�g>�yRXP%� &4I�ŁTu��ډ2�@��sk�H���l4X6(l��Q��a��X,2S��1^r,��?����� ��Z����������C�^b��~�0nX�X��΢B[$�|� &a�z�ˍF�������Z��l�u)�kM&�+���壗�1wA���$���s�o"�&jP�*@�P��t֨ߢ;�{���sK�J��e�G3B��s�V5�1��M��x��Ca���b91T:Alc*s47�[^���Xv��ޫ������s�^�����.^�2�bS����_|d�rͥ���X�k�HR��S\�$����B��Om����3R�ʌ�|i5�YG ��!�1��/̸=�jZ���م���2���b�u�x=��O�^T8 1d�@q�ꀘ��×Q5�Z�s�b==�R'�� Ft��-�3$�l:�,y���U[�)/)��������2�j�l�X1�3��}ҟm���9�`}�^̂X�<����5�� Ol�;G�u�A,`����-�a�����D�G��z���6O����d�6}e?(sG�?�b~��XBm/��7�O���u�ɮ�L1���W���I�D�X�Ð�'����Fk���KX�����<�6?3S��࢖`����r_�b��c���ak�d�O>X�X�mr�>���6��,�C���/m��'ף���;k|��OUYD@�qq����A��E�I0l���|}� v�VN�ؓ���LTIU��3bH+'�	�Qܢ�Wzs�2�ȲC���I���JZ1,�MEk�W"C�"~�\� b����u�����F33�KN�@l�5L��eoL�`^���"�#��݈Q6$@C��߂�C��}~��7���0�w.�~�+�H��� V�_��i��t�/R;Ix*�b��R�r�S�eSF�Ԧ��R v�꨽����}Ѣ��L>{W}�j�$zG���⭚�-M�+���a��PP�P�ۂ,�.
�+������n���Ju\��"����D�n��h������x��R:�R�6V�G�ք�l	���~bۼj^YK�:HY,-D��C@�S1`��8
zy�=LȏʴM�	��O�8�cԙ�}M?8��+�1��!��>5��<U�Y��lM�m�Q���#C��ɩ���*����A	+�ݬz:lEΥ� vY�7~�l��8�Fw�������aw�[�M�j%<��s0�1ȡLk�W�%OH��iH���%�O����8�6�E��IN�|i��{ ��)���~g���$��T�(6��њ.�h���UT �(`�C�ER��ii�FA$�7�%R"�!��H������R����:s��̹s���wמ(�{C��O�G�vxO)m�]���jQ����㶷8.n������c����X����b��?n��e���X�*���/�jf٠��R�H�5������8�VN˚���t�����E&|��H_�\��Fa�VH=���q%�
7ߊ,��>�tv�ף��-Z�g�nZ�[TlAIf��!�|S�^^`�5�엪-����%�/�[�xG���ćk�����!J��U��"vE�kJ�[�P5b�=$gεn�5�q$��:���7�BxϞ-���&�h$ĺR�
��>�	\�G��IvC�ː�B����`S�
ok��={v/Ț��u0�>|�D
@�r�i����~���V��/��!&J����_�b,�*.�2-1� b]{+U�iN�{.dO5�r��L�Al����jbw���p�fx�������D+;'���
%s@�B�R~d�fɔ���c�� �h�Q�a�L���]���k�֌��]�[���l\���e]6�6@+��Mi���"*xj����,Ϋt9�]�(a�o�:�Oe ַP����(���������f��b��*�%=�[#����I՟D��Φ��0"SxU�m4�8�-��}k X��]
��3�D��id*�K�f�gܔ��IT���V���rb6���m2}�b��r�2�ҳ{�ѐ��m����/ӹ�3��xb��u�����/F��K�B�O|�[y�4�p�Y��61s�b�k�xo��~�����I��=�X���֖ z2r��ϝ��)�k'��J�J�<3�*��>ce�1
�)[�
�#���f/nԸZ�ס��!VQiC�.�p#V��~b�J����o��Ȏ���O���2�gOe¨��h���B�m�����:{�}^Sȣ2b�r�f�w�,b&Y�l�V��CL��IyS9�p(������@�a�be�3W�������~š#��u��	�4�֚n�����P��x�x�_M���y��ݸS�^���p��صC��c����� �'M���3��y�so��>��Y�:�߬)�T�y�b%VZ&d'A�?�e�Nq��[T F�ff���_�ܙY���O5>1�o�4k/��&^xvli��E���C��%��D�U��QqW9�) &nJL�u.h.Z��R:��nY1N��1q��]�;#������+�_ڦ���ͮV؛�-�6��d{�<m��(�λT����Md �o��)���w�ҲtC�\>y�b���ý��,�ʧ�M��G�AL'��x����J�np�����%�
�V�����*�_�YC�dŴE$pP��I��2�<�o�b5
]ׂM�Z��곩�����ve�A�ɢa�Ω.(���w���(j�{|�.��*�n����a@@�B�^M�͑"�	���h�9��3�X�2�7/V�.��.�6յV��Ӂ��n<���rn��D[�'R�K�tf����3���ko����1��U>S	��W��ëǨ!&��h��s�<��D�j��b\C�9JG�N�o���CLڐ=qa�/A�����!\`�	�~f��&�)_"�^c�i��]BW��l4=l~J5�(��Mr�aČ�^�s��mpwo��&�d���b�X���Lݯd���ܙ� v=@.<!0B�A×���ʨ��	bL1Y��$5�rH���� 9��3O�!ƛ~�֕�� �m}��1��w�d&k��
>՜��#��A���/w����&���1>��C������廪�y��Ή�����x>ٽc�C2F�����>�:W��ɱ����,&7Go���ɞb�X�&����+�'\�G���V!�u�ypI5Ir�HR�G��w`w��o~O��g��t���V`��iD�-�6%��#0$Y����)]��y�b��q!�ÄI�?S�n��^F��)��s�qc���gmOV]��֯!F�/H�ؔ:��i����@}
��E+�&���.�կD�t5�Jp#!�;���?:{a����������e�"����8?��MW��F�[������I6�i�K�b���x9
:�;'�J��a"!�=4O����'L���8��:G	bb���Eˌi%!lB�ؤj��Bx�8���"F������y}�76��k���4�����'f�Ҋ�^C��1�e������G���l��[��Fj?��X�ݵ���΋���9rG'�B;�˖{J�>OƕY�b����Bw�C��TUcR���+mż8�X�ݥF��
Ek�.)�X*��3�;�y�Q�.w���٘	��O���ƎX��]��k���0�I�{Gq���*��r7翤��c�M���[�G��G�nB���<4�N#�rg#�oxYp5.��P�c���}t�S���x�bC��r�������f�l� 6ۙ��S��a<C��t�Ş�>�mB��<�����s��[4��DĻ�ϖ39�?�0������p@L/��$O�Ӕ�P���q��ھpͿ�/x��^�<c�Vr�b��n(*�7|ǹ��}���YC���m�|�<��k�((�nIb��3���(}���lOU�n�K2+�}�����ќ, ���A�i��tb��E���[���0�ڳ�1Ղw &+�א����{��}^yC�X^�E�'Ӧ*��ZZ����1��w1��zn�C�'/}VF�e�\\W!�[��j�IH`���ĚK�Q�?��F�:��ސ�fd�ݵ7�ЇXP
N��1��B
�����Y����g�!@0�zaq��̫�B����d-����w҉��)I�{� 6(�ֺ��GZ_H��}ab�bb�*.��O7��S��mD,�!�^p9���t�~=������&�P*��rM6
1��#��>@L��H�|�H����A���Í�h��9�6+0d�\��6o���jC�����u��b坎Y�ꃇ&�{3�n���[ �B�����zk*��-)�.�h���ZDL;��Ǐ���b2�����ߙ���(��?�/�i��Lv�a^����
����
W�=�X���m�K�(�P��zR�C��5$���z&Zb҇��)�B���>��~�`���X��'�^�k�u�u��q2�u��I����iHEJ�mz��cJ�a@�s��k[���bw�K�#���(�,���a�8I�Pt<��.�؊�dр�!��*�9���`*�~��nw=��2� �N����I�p�e��m[�I�ޑ��-�E�_�>��
��23Ugd��y��%d��� b~C�*��2]�P���`9ɀ�O�I��,�U�*�!�uM�8�|��r����҃�k&Ů��T1�L�<�s�Q|�����g���� M9@�8w&��)����̶b*��Y�[�W��,�llH���~[��p�����-�� b�/�O�>mw,�_�=]y�X�d��R�>����%^_�/�v�w>A�X��*�s1�?���O��U�]�4��k���S��nf˛���uMPW���4�����_�W�b�H@l�U^�e��9��"dK����lP�,	3��Z�>�!Z� ��9r=��є��t�r�Om|b謿�����N��j7����!6�"����6z��kT��H#$�V��j��=��	֠}�o�$]ʇ�ƒ*�C+;��Q���>	�P���Ii�Qo��c���{Âi71����4=�Q��t��K��h�A���8��*���6�h�Y��X���1#/#��O�1�����D��ߚA|t�~��n� 6`=�;��=�ot�\��59�[�?u@�9n�ZG�f�N.��[��w�Ć�z����M��d�	��:�x�!�ܘxe�q���C�����.��˫�XQSxx��\��4�B]����C�m�J�	:��c4E3� 6��C2�{]�z��x&�xm 1:�}i|�P]vM�s�G���˿��7"<I(xU�4����g
�<>}+_N��-<��N��N
1�'���'v~T��4m&��f �v{��UU��UuIڶ�&ҝ�b�ʜ�߶i�S�pE%)�{���@�l��Lݖ�����I���~ s;İP%��ԝ�R(|�$n�|��l��2��n+�z,V�>�|���n�֕��ۖ�+���G$��^o]���'62�K{�F?�X�Wr�[�x)��>�vy�h�6%iA���x��S���x��B1��[nO��.�1�w�:�v-4b9��$ĉ��r��|$�H���b�b��"U�6F�x���
)}!f��/�]����=+��x�Te�,���jA�t�\���ջ���(��{����'�:�+��������OѲ���Vmh)���X��ֳ+�5���i��EA�k'[H�3xw�'��mMhQ�d���7����p���|�h�1cU��6�2Ĝ�N��jTE,���QL3V�b�κ�19?"~�bDpls�b�6��E�ˈ�w�K���,{_�U���׸�3�ʽ�$�b��M�F&Y����q.�gMPB����%5�ӯ�(q��2�0�!�"/���0�{���W���9��"�l9_9E�\�#�|�� vt�f���ǯ�֛��s8��kג�e89����3k��س�M���z{�`�5I��8t�mU��
܌��5!����Rc�M��Q�
+~�\2��b�B���M�ez�Ǻh���J� �"�+-R5pV�4k\z�/����+��O��2����y7_�&�C̅�[l����v��{{X��!�d�Dt��j�L�r�6m�P=�6Īq�q��*�ɼq���*i�쉇Xp��O��p������T���$�hM��*�g,<�*�Rdֽt�v�K���;�ojr���h���OBl��\��ѣ��ӡ��4�>	#�ma�,���W�H�h�y�T���d���]tv�wmǾ�~��)����/�/�DE�c����_�g'��u�Z�SĤ�e��UǶ�rgH>�z}%*|1�=��{x��?�,>����\�[�=�����7�e?hV�%�Eic�������1�YY�ؖ+��/��ɇīw��!�J%��I;����3�S��	bLv!����餲|�
"jo�?CLH���, ;[X0�%�Yi��*�v��ؤ�z�
O��w����V�Z�'?Al�y�ȡ�cN�<�;y�{���{��lU����9u�o�eT=��M����Ѓ$��DwA������1�/o$��[	��Y�m�-=��XD&40���
�A�,���������m�??��q���aoŻ���ڤ"c��~�����m�u愲rb��n'8ϫ���F��A�}6�1N*1y?����Q:��19�$�Jiu���-��1z��������v����^Tku���W��p��?�տ�����gd�>�dU$븋��������~I+�ze��EF&_�!M�0
�H�C����~�Y_����hg� �_a?>�h���w8|� ��Ȗ�B�Ȟ����K8��7�ޔ=8�{df�M�&�=3��w]=�����������T��>���}�����b��N ��1�:��
��p���곷b�**R�IzkZ���]�"R�� �������:yE?��i��y耘�G��&������G��dL�� ր2j����M��q>��B:6b4���/�&^�£�e{A�>$q��g�)n�m�=q|a6܄/ �H+d��=ߟdw�dM5�׏��FkC����G��
^����e��5K��2����أ� �_a��dbޢ��=lES�X+�\��0@LR=U= ;A\�d롥�����Kv�߬H���Y��C�<�d^�Y�Ěb��LT�z����Ia:V�F����S1󇌸PaJ�Ms�l�o� ���a�~L9��B�bT��on��a]2�˯���4�aV՝{���'����o��|t�u�Y��،�`�b�Z���&H��J����;#6��ߘ�A�Z��}ޞKo�7�[A#��=\0EU�S<r(Ιs��Ф9�P�U���'�I���a��
���(']��l�Q�3���=����>�:ME\����6���e�2�<t�|8/Ҵs���G��\:����Mg�/�lSdԦx��~`1i�ȅ9\aW=�3�/���lj�nK.��&�� V���9��3orn ��62O b��	�N0w����h�P�h-s�ALNiC)��v���Au�^���)�U��עqw���BZ��F-�y��$�֒{z�g!g%~�c

n����@��q�#��זU�)`F��1̱�4��vc�d�d�Ⱥ�5 �+���sc��	��:2w'ϸ(2��
����Y�ʻ�D�Ԗ�Ob!w8tR\#bd�oQՙ{Õ��X����]���e�Ώ�t�$ 6u3����M��z�Uq�̊Y ����?�Տ��`/HK�̹�S�f-W�<s)^����@�����X��R�a������Les9�-E}eYK 1�2*�R���7��M�z�u��r�ժ;b�"m�H��^���"��)^a���~Ҡ�Wbm������b����PbSRg�
{^%!�=��ߵ���bfy�1��Nyڼ�p�ᇲ�K���r/l���}m�=��y2�I@���xmk;S,�6�]f���`�l�����\M|��Iԓ�����:�I;��>,��d-~6��'2�b�]d�Ă��	��<���j�g��g��0�_�w�}�^�{��e�!�H���^�'��JV٦������%	��lX�1����f>���+=�t<o'>!� bB��"*��=�^���,?��,��A��<DkǪTP*�#kN_'M�<��^�YL�~}�5��f�����JH��v�����n�Cͧ=
4��-v��`5p{�Y|a��� ~���8����U/V�����/�������+�<�ݍ����l�hԱ���B9�zb�Hz2������mZT4tSU葅@l����9=&��;S-�w���d,�����}�������%6�+�0�^���Zf�P��4d[��)���Jޔм��H��{� �DkRV�$�,:�8 ����W�O �1�Xl۸��6[5n٠~�)���K��e�0d:H�kvp�1��Z�	��5�s���֟7	n�؈#㓟o�^�%�D�(-��
b�J�x�$8T����ee-��@lZ��/��41�wP.7l��ʣ��\��ߟ��Z���"g�V�j����$9�%9��B���'����TU���K1�&�`�=��o����bs3�� ��=�v�T&o�_'�����.�����'y=���V1���9M�t�p�?f�&�jh��y)�H�xO�q�U���Jn��sHGƆéha[8����L�
��G��U�fa����~t�K0�D��p/��Y\��5�|y��qٔg��٩�ok V���ece���H����i��5��!S�"���@���T�G�"_U����z���g�p���p\sAln�p�d�nVl3!5T�N,�^.����2�����d���A��ؐ��c��	yL|*C龒3pO�,���-�Ͱ�BVy&X��f�`8��b�h4섺[�(0Ͳ�N��>���6<p|_B��g���j�b�
���):�Y����*\��`�Fz�af�}�����zo�I�Q��X%���a޸I��>���,O�Z�.bb���O�\J�"�C+R>:}|b�JQ��-����J�P?<̴Ĩ7x�����ȯ+�C�o��X(��WsC�6v��='ѩN�_Z����%���D��"�Ե}���w�@��Q�	G�>�u��S���_�@L:ε�=>�EӘ+��w2���������ZDn	S��S�>�����)�-8i����3�U
�~���ojlb*Z�DnQ�}ӈ}&�;��KkN vb}� ��pT<��T+�V���v��y�U�3b^�x�]��0¿�(ϱA�n�H�.f�^���/t �_���4O��
�����(����
���%���ks�P��k��r7~���)�:�!��q��g17��Z˘v� *��]��P`�s��y�4b�tx_�Z���o��5���i�O�Xz������g��|_ߩ}qza�W�U��:��N)�iT?��ċ���b��=�j8��ԯ���ie>�خc�Ϊ�B�����"�0|c��O�:Xb�"	��5&C�uq�Al�%k/ /���l����|�Dh[��Ύ��zu��R��\}Ԣz� �Q"~�Òm��Pjk�K(�[p/�_,���~�/���
Ǆ��R7!kSz�p�z���R�h�c#:��X��]Yn�al��"j�KQ������6�R��������.ۨ!)��@�؞g������Muc���u!��y��B�^���q/L�T�nµL"հ7P�G̢[ǯ��?=3]Z�,���%��]0����|�, �b%9]�{���b�nj ��czR���1[�j��{�`{9��0� �r� �?���2��}��za�k�޿��Jf{��~�����q��a=0|�d��0@t{p��D��c��^[�?O��4��,:��1U:�ɷ���6�J����Q�d�re���������}��Ψ��t �p��:�$â�%�#]K�'� �fu�m�vZ��3S�S��"I�zS��蠅��,M>��ɌF ��ﱨ:����܈���%(� &NTL��&�a��r�O./���#�J��q;2��,��x4���i_�����P�nIN�B�u,猄5�����T	�s?FP��Ъo��J��L�w'�[��8�E�t�怀Xٹ�=�@.��/�8����MTA��l����q_�,�>�D�����i;5�]-�H����A��R�L?�d
V�0��})�����qa��jaS�;�|M����A�d2����I����҇	�=�i�����M�A��n5� m4� �䂷J�� �h4�(�9+���vX�;�Y;�Yϼ�4y�f��\��R5-qW>�=,	M±��V_e@�x���b�b_ۖ`|7<��X�"����@̎�-sI�lL)!v��6b[~2�,�Ǒ�Do�X}��' :��LU�Y���cl�����g*�M�E��<�|�����;��D���U ;׍�t����f�>?�J�$^W��P�e�H��j�3��8,��;�s+�T�����ubdK.��ӽ����u$�^k��؝�"�e�����LX������zsV�� ���&�1�)~��F�Y��ȩs�׬9�n�J{b8Ǩu��C��~�e�\_��w(b��V�9���y���9����®zpa�w:8�:.����СӒ�@x��$ld����'��v+�q>��Xko5Es�V?�퉪di��_�?�B���w��m����$�A�
����B�����J��=�4�Ѓ�B���~�� ��P׆ẅ�C����E�cHHb)ފ�,�b�Ч��l�ˢ/3�@� ^%c��)��C,�sO��Ĩ�F�Q��:�VY�D�����V�l���!�;O��6���� �}8�P�q�rh��s9�$3���A�r};~�V`����A��]�V}c��Lt?��%�4�Y��yS/�y���b���$��F϶�kU��(�秂X����k9��z>�7D8�;Z9� �л�v��ݤi�����'{+��@L5H��;AI&���S{#!�����H$����nQ�����2��� ��V�@�z'w��8�X�����b����(��z2��,��*��W-���FCY��=	H��b,	ĸ�';�1�U6~v�7�E��o�(�
���R�*ݢ���+�=C��������ט�ߊބ��]azY"�q�s�}�[��׬�L����+���c��|et��|��:ʌUB[q4�-�$Gl9�p�I���E'm���F���<��'��bה5Ƚ��Xgl~>6�C'<��IA����m'��������r�@jA�w8�!�:����'����d�1�ߍ!zb�%�}��]���z�p��u F���񼋽^Q.��>�h�q6��$?�ئ3�T��Q�"�A'��1��\ވ��G{�I�ORÓ��[cALA�p��}�FpĚ��ҋ�6w�� ��<��P$t��Д������S ���F�IG�b"���`*�Z�A=���cň���%�K�>���Z���fU�7�nJ�+��Eg��- V��j���+:�B��NUīb	Hc%Z���;��zv�s���O|a�-]M��f+ߧ���b=èY�a�K�`4�y����S�jFq"G&��,Xmh��8/�-��o���!=O�>�*?n�h��e���J��b�`h��x0������L����W�"���}2M��۹ί��X��}qnE��*���Fa6�>þ)Kը͢Û����b;�o1��~�JF��+��W5�F�C�$��g"���rrPٽ\��Űě��<���0�+��a��"��B�ֻ>�XGR�x�n�ض��v���-p����zA,H�����X 9���E��|	�m������z��/2������-���x�~���'lm���	��=��1�$>Ufe�}�n	�M?�1T	���y�@���i�<�GqX7�/����߻�|��=����8+����k����o�xWQ�9��4����-�RT�)��!.�2륧0�Ц��H[�;�b��[f���	;c�;~�*ą�O�A���\\��v���;-���%˩]�`����`j(�Iՠ]��"�X�c%(�dݴ�SO�U�}�ؕUO�dB�'����1�S�Ej�GVB���v$8FA,�Q1����ފ/�t�L���
�:�{)�-ǝ���}�ȈJ��8Jy�B����ӽ�����w�̊4
*��y�f��m��,r��t�7Wt�qx�{M�������X�%�,-Q��$���ZE�a�8�%2��z��������� ��lP�~̎c���8Sa����`a����Ѵ�?9��H9Ȳ�jٟ�������H��/�On/�2K���(R���6��f�Xc+�ItW!��VR��E }|�%����z`tD	؋C
�1��ㆯ��?YŪ�bfX�n�����waP]D�ѓ�x(X��G�V�!ΏQb��b���;�x�?�d�k���.��^#s���h.�hXZ6�c�1�������Y���� #�ia���;���h���eTl� `@�)�F`��AJ��Fj��F�P����$$��P@@»?�s��oݽ��}��D�=�o?v:ځ`௎8��0�}�J�	�A<�n�+��6c�䐔=G�j��2�[��fQ����:�i�&F���?�j���rA�S$yw��!v} Y��tr�?��KSU��_M3��Ш5+s-����%,W����MH*�׳���@�X_�`�6�T����V��.��Q&��e�е����˪������A���e�t'�eF�hߜ���md��1��y.��-C��AL�^oGc(ڤ?��b̆�B��~!i��aW�%22�9vJ|�`1�"���5��b�����:J�_�ز�yEDF��
�?e#sA)���eg��y��9�="��ֻ1>.*�&�)�%c4���2�mcz�b�/Yt�SKCl�c�ϥ��LV��Z�����h�7M�A���	�c���ɾjN���K �KRS��>�17��?M������4�\(�Μ+qj���0ֿ۬W,���G[�Zf��$<ԮĜ���(
(^�J_���_��6�/ ����_��L^x!JL�YK��)� �1Um9�ó��bؼ�-�o�b<$�L!���w<��	M��= �y�%�D�q8�o�>��"���k�v������P�	�+Z9�Pk؋77)<���_.Ifi�E�$�������Jz�(KOף^#\Al�R����2v6��~J�x�=n�G>p�����o�,�� �� ��t�F}���۾�`d©��"��D�EC��i�-,,>t�y���L��g�7c�P��{n�O�Y�@,�.R��?/ֵ�JZ_���b���vib���C���^K'� vY1N�a�H3F`İ%4N�"yĈ������lJ�7%�YcBGYA��a��F��_���)�_�V��� v,U�!{��[�W�j�R��9�1���#_oK��U������Fb�~��bF����k�'��-������7p���UK�l��j�������ܺ	P6b�Q� ��&��������dE��K��ږ߷�� f�\Q0�V�'k�ȣFI�W��0b4.,��b��vD�)�zC3���@�`�/Sw���1�1���n�>�%<�4���|nyuk\l�u�N�8:Wҋg�l����3~�"$�5l@��,<�*����<詑�ڋ��Z 6�6|"��{��5+%��;{���bw�ײ��nI��Y�ݟ�����n8u�*��(���wW �5?W˚U��kG���x�{
Ė|8�O]�x�e�)1����X�w�~�T���Ă���>�ٷ�+�إͅ@��H��W�E@���6�YrA�-�@Mwo)
b�Y�<(�?��z!��+��atnc鑠��;�~lJbt�I��ڇ�L��L��ҰU��zJKv�	o�T�d��^�k1��16ؙ��ԘY[M�싰�@L�z/�L��q�ﻵ��e-D �a�a�`XF���W�}�����SN3h�4"�;�c�~����b+d�'�Oͤ�N#�e|��B#� 6��;���+�+�q��$���3vs�,�����D�U���D�1�_�����U��D�L:v�p����D{ݞ��܅��6��w� �myv<&���i�e"��YV������sy�$��ba�cOX���q���i�}Ƚ2q��I�L/��B���X�!Ɉ��b�ͭ�XY(<<rsD�(:�d����wko-I��Ţ�4����ͳ��� *%%É]�tC����V���m l����ʛsʡ�z�	b�5�{(�u~$S�`d�|�� Ƥ=b�{^\���w{��qy�b��^~�s�4q��E��ف<�1�o��};#�(>+]B��@��p����3>�d��%��_=.���&�n���TfΓ���e��#U�rwK�0i��mY�u4� t@l^��w�>���^K��Q�A��Pi�̸�0ۓ�@]�\���@,�B���]\9�XtS��*Ģg�i�;H�N��6�v�/�JKb,37��~`�G"c��dc탘���E�EƇ*��ie�`��n�%Te���քR��_�9�[������Nk.��{�3�h��q�Q�F�+�'�`���tR������L�P���y�o<W��u��s��q֘���"�坷1&����;����S&�/�Rw���\d����:V��3�#֡�6���8�� ���Xw5d�{�}g������� ��;]c�y����x?�&15���Nx���4j��U��� ��Z;Ib�U�IN����В�b4�溺0��W,�9�����	u �>Y1�d�����&y[���P�T�2��{a��eY�ܴ�Y���|$�"vł�M�Z�(7�b�;��i��д��'��QCo��)}�!қ��Ʒ��r���] f��*x�mm"�BtN���S1�m�E=��薡M�4`�&b"���+�wvZ&�H`�iD��"SNS,�8�?.�`�z�� �G҃�0<@�!�Ow#g�:��3���w����;B�s?��#9�(|��y�eY�c~��^Dc�7a��m?�ov����{��z�÷�cr�B�H��sQN̡_�[e��%޻1�U���9�'�c��1��+�A��ԇZ~1=)��WL�m�#e)z�	@��(����v�w���3�9�G�L�r�RX��f�����N�7�/��/�J��'���O<^DE�W�ByA�rG�}$U����3w���M"+/-Y}O�sY yv���P3��qS�,6ӛ���ub��2RA��I� d6�f���Gإ�F<���r؉��(�?=�U��J�bh�)����y��LB���r�����Z��R��,ͨ�e9Q��b�@�/��$����9��-�SQ�ϣA�k�\/Y�!�u@���|͓/ ĒGφE�U&"���t���@���>?��K��"?>����Ķ�儽\���a[_��e��X��zH��EEzR3�Q��ۋ��d����tUs��P#W�c�O��%��r�A��B�e�~M�B�:]z*��[[�n�)��vZK�O�|1����,����Ý'Y��M��� f�����]i����Gi����&db�c&����ZNԂn��a+��X$�	�6ݛ@�\4դ�m���/���˓'ϙ�}�+��L���|gĂ���68P|�q:�8��[S��⥒���ۃ&�F�.�1�]��cv�_E^;�>���>���b�D���?�+5*�B/X)�@��ׇG���Dz�� �����:����O�n�%��2l�Y��@̪����Gf�,V�+��Jt) �>��b�d�����Š'� ��/|�����.�8�p��1���cN�8��U�us�h0�a���1�刚92��1��,ZH�q<v�!�-�H�2tޘ	'[0	z=��a�ˆ�`��*��c2wh�q�\�C��Ŭ�f��Ɍ��,���eQ���j�ȇ]�Y�����[��n�M�k]�@�P��,�
2uqɋ�	�4.��4��c��WM�X)ȺH��1��)D2��gk4u!��Y)�w�D�DRE�
����G�ׂX����|_����gqo���y$
AL�G� u��[X��q���Y2��n�͘;znRx\�v����E<��x5��u�X�b�hR���ߍ���g�f������uk#��@,�è�I��ݗ|E,�'y��|uĖ!�+;
Q��}�	ˢF�^mx���g+#�d����٫�^3����]��bӰ��z1��}�����]��:�d	�A�����9���]�/��@�pd��a��`���W�P5bN1�
�v{�i4骊�+A�hR
A&�$i�m�p�S�w��1m9��M�;�����l��E�����`zW�An��C���H�}v�˯K�Jѽ�n��Tm����bZ�B��֙:��!Pqbs���ӈ�<�R�D~ګį�sҪ��FY`"�ZO����ZDv�_�7�>�C����!3�ʊc�AM4?�����݁�5�M��_.?�cC1݊b
�L�T,�Ky���h�#�K��ݙgE��W̨�X� ��Z���P֬�'����+����@��
�7uݙ]@8��;UR��E �����/��N|��!0�+�"P����YCZ<?��\�؞��@LoI�,6��(�]���q�0���Pd�h_}稜+:�O�̑��bΓ5w�R���p*-���A�Y����`#)�����|%u��	�G�ה�[�Z��BE]J3@,��='cˋ
+wV[t�/_o��@LLv0� ����sNb+�g�����d�0֦G��Jg���A�)8:�^�s��e�>���bi�7��6d�J���2Im|�XU �'U��w�+�����Y�������O�j�����v�k0WP� ����+Hoqwq���}�bn��S4o'vn�}�È1�Ş�� �Q̳�<b��MHHo�b���������~ڌP�b�c�a�a��U�ŃX{�Q7�
����l�ʘ���q�� ǣ(8���=A�V��I�K=
�Ii����\��*�,_�1~�o$%��z�t�V�ڌ� V�O���B����@��0�.�M���r���MK�V�q��쁘��/�φ�q��ʢ|Pzc����-zǾr��%Sљo��3���{
�%坹PI�!0��k_,|b�ů���fJ�=Ktl{�Q"Alc�9�C=�G?Gf9CWb�Z;y����o	h�g<rk�4�bv1�j����<�M����Q%<ރX�u���{oI�̷���uC)� �$>��w|�aX�er�DS�E�L&�u�w���%���0�>f�b��L��#��J�!f�c<��UC�"�~f�(-dЅ�䠿��1(g�d���ܚ�ͫUa�EtRJ�F���`�=l�Շ׻�{��@@���<���h�mC�W2uڗJ[/r,�%�k�'�m̽#e��b���Ũ��g�<Z0�ı�U�p�z��^�#���8jyb],���N��
��Z1
;���A�ݸ���u�WD���V�1G����ӯ��bQM��w�ݑ?A�ח����o��~�a�m�$�F��P�ŰBd�������!���B@�~������+�\m���pC��`=���Ƞ����]�[�@5��Hd>ݬ��M���4pʉ�b�4���XX��D����jY�	��]I��^&��"���4��j�dٯ����;�)/8�c V�����ԼU�sxu�EG��|+�(�P]����xOF��%��d�d��IهX{i�]I� fzI��Դr��ynz�C"�5���xΝO��\7]6]�8��>-|<��R&N�UZ�������Ger����0,�%ym@�I3V�h��F��C7��4��X���+q~_.�/v�M�-��Hd�x�ov,J�P!�b
�7!�S�aC�s��E�K��h�s���:�j�k#�^.qb�2.�?h���eXh� P@B����[R:DJ��.AiP��[J���S:��F������߿�9�1Oi�����R1ĸ�-��,0"u�.��Y�
�m��]+��#�ܷ��lYk��/��:�;@�1q<��}��[d�AL"�T��.��@�Mߓ�&.:ެ:��I��)�XpF��$�����1�1�g���r#X���*�e�i( �v�\��#�EF�.��4���a��g�����L5'U��U4��܏;�q�n]�u�`��0�F��F�C_r&S4k�RJez�&e�ͽ�l�ơ�"O��� �Ã]b���E�}KP�i�W��lН\ v����Ub��j���s]:c�|ӌ�H�++����!�2���
�N�>/������N�&������$1��)J�{u���VG��� �0�� �8xp���U@E�^���ى�T���#��d-�
|D�1K�����2��7�)�K8�1������^��f-V�<Ir ��o��a��g�W�D4¥�b

��0�/�t�dZ�&Ϳ1�g�&:�~&��B��i3�Z �"_�-�� ��y;z3���7�$����zӑ<|�����0:��PVUz{}0��!)�y�`-�����l��A*4��I�2�U[��:��rZs�'}��{��b}�+p�5�b��řA6��vqc ���Ւk���?uN@U�r��0�ݨo���֢Ĝp��oR�V�Ĭ�r�˛P�˸�UDJ3=��1K3CqaLE��y�I�(��޲oAl_+��k���.�@d�m�'���S�^*U�D�+3�q63� �Z���T�-wqMX�%[K��cի+~G���O�2�U�Z�|�Ğ�m�V�6ۡ�p`�%
��1���C�"�͡X&;$�n�sj �v�j�C�O��d_H���bC;f����Ƚ�u=�0� �@�����S��>��a�<��Ģ=K�����jc��g����Al+p�%;$��Q렷��睘� �M�g%�F�Up�1���
��H���Lw'4�������a"4�A�d�r2�V��\|?�����Yb1��r��'N+H#�4��I�yb�l9p��3���iK�?O4y�X��nȊ�j���Kc�C��S�ݛ�b��A�q�2�\Nc 1��}�8��0ڏ�n��w���1����O�B�j���C�[�G1}��f2�z�/��#��L_�ع�G�t�|����}BC1E��>�=���!{5@�D;�Ffe�S�/�b*Aϣ�R��<�)��)�� 5��pb�SV[]!�P����g;�mc."��e3I�xy��L�ٽ��`�[L�BC^׏l�Ϸ˷�G��X�m����S/���}�7|�>�XV�����מU��)#�B�������h�K26Yh�{޹Қ��ګ�[��'��uDs�o�L�B@�����X���ҥ7r���ˤC$���`c���v���fmt����_�Ż�i���8.�r29��}G�����#I1��^�5�w�逘&�uvn��k뫙[fqn���\ �K�H�-���q��.O��"�ĺ���7�:�LJY�K��@L	18����T�2f!�]�/��l\mܨ/�Kbt�$��\q1��,u%��������>/k�b��Z,u,�L��pM�v�<7�Um��l?�&<��;��z�b����R�l��(G�T��ذ�AlL\�Q����Op�N�}�W��X���tP0;Q5|�FX�@���8+ϯ�U�����N���	�y����ˤ_r6���P-r����J��v>z}}H��d�^��b�Z�Q��Ω'�z��7��,n��	��JV���i�~�(.���X[�10C�����kVߤ/˶V1�-���Ʈ� 9t��j�2@L�}˾��m\+�(~6"~6����S�8�'y$�EfK�M0cȃ�e ��5�UM��"^�_�F��@,�$MQ�{�]�TqGE&�h�H�K�Wg���˓ᵆ��#J�Xx�~���)�Pz#o�zh1\��������Xy�H���ѹzc �Y=����;�l2,���57N���V�s�����]ê���hq:C$��r�{k�a��ߋ��O�5Ķ����)5��z#I��`&�?��ag�>�|}]�d�5�.�"�0��.��0��$�,GDD�Ŗnb�X@s˨��y-�����9⯶H �@0���l�hMK	9��N����/Ӧ���W ���L��ЇJl@�k�=�����@7iH�TW��fM�*W�+<Ƚ���dŠ�����BĹA;��-�5��au�^t��mlS>�;�78̖y�$�b$e��H�	b��bƣ\A�� �P�Z���ڡW�TZŀ<%�b��i�������g$`����X�V�I�����1��.̜���y0f#��YGS8�/F^Kc�b���תI�x�����uC�U�7�o������f2�,�&��Dkb]�����q��y�+I��M�Q`D�˙�THɓ>&~�����ʇ^�d���O�=����W���Dk���i��̯�`�  f��Q��r�5����g �ҩ$�mdw��ڻ�em�<wZ\1ĸ=_��V9���\�R���� ����"�kQ</�ZI���qE&xbj4o߱��
j�����o�ʇ�X$β5�ꧺ����'��7��<@,}k~y+��+0���!V�u��;Xw$�t�9��/Ȁ��y���2N�0i�_:$�s�π�J?
��i7�rH��Nܧ1��2���G�X�MD6D� k�N�^�f��q_8s;��b��������D��b�o�0d��	VY����g�`�c�X�8|3&�Ă�j�6��(�2�M���}�̛	l�M҈�����T?k�z�dc/�(��9{�o�\���M�1'��R�[����&���9��'�}Wu]��@�$�Vu��?>&�N���&��� ��aO~57$��r0_��p58�n �0�އ��_NZ��GĜl��K��Ɨ�WW\�yr��	g��X�b��L����fe�� ��R|+�N����!Ҫ&Y��������0R������jBZN��nV����B&�d�ӻ��"R� &1$x�]JMƎG��poHb�?#�3p]�|�A�^���׀D�X7�6�)�}���#���Ϲ��AL���)U�־N�C�=������|�4~��|�=_͚,�a���ѣ*Q��+��-Aˬb�ð��o\�']�7>GC]ڻbT�!�-�3>dv��&�#��e�w������a��g����?�45q\U��� �E��L_������o��-��J-�z)�SC,U��z�$�W�W�E��D��6m.��o�Ʈ{&�w{�(�/��\�>�?�b��ȹ��=���'�8��h���ۗ4���,H"K�C��w�?��z	̀�	CG�퓽�Q\JaiBX�\#�4��-��$�F�dm�]�Չ2}�k���]�Ni���*{���U�e9�������;�����ə��NV���F-�Fb���Vg|w�Y
�6�
b���*��g�f�"�J��� �`'��c�K�2�Ñ%��l! �
��7�g���N{���$6�c���_+�|���}��i��� vWČ�>5�z�>����7���`���S��Q�Gy��OV�?X��o,�#*�MI������(c	�6 �d�U���A� �JG�d�K������=�c�|���Le��ᠧὢ�gbo�8Pb������:gb�d���@,��U��л�z�F6/!;l[	���-#��Π+�^'e%����R�׶��agdWD���7�2��γV��>���`�M�u�@�`�v*O}Zh�'�ی����Ts�����E�<��E7v�D(�{�v�bj�4�޸)�B���I�!���<�$��%y%����/��@�k+���o+��.N�
�.a�{!�;���Ke�(� ƢE)�򉡑� ����'A���E￟��X�9�T:q��1�lϵ0B"d��u���� ��+��u�ۈ�20��=w.2�)�ݸt�Ip�.$a��f���R���x��y�T���X�Yr\k�KQ Sh8f��{1[�~�2��祙�b	���4z�[�������kp����m��r>io��'���ݝ����%9#�e�^]|��T�-�X��?���~|t��Y*�N8���6�`����.���������nM��*ӱ��Я�~qx�U���I,O�VM$�[��~U�u�>�������� ��_`DI�@(��1aV���;�n�X}]��+2�3q��6Ij<���?7?�u]�N��^�)�`/�3#��l�;[����DO�,b�B���?�#�����I��V8Ǆ]�#;�q�ƒ�� 
�Z�%�7�8�������|:iW��3E��ű`f!T;_i{�?�DwˀRl]ȋ1V�+67/�d�l�w�>E_J��&Y}���f�̈́��?7���� q��vd̒������w�>���_c?�J��ۼ`2(=^�~��x,k�ߘ��f�[���{���#����=��/��Ssͮr�)|*H�!�,蹨� ע���lp�>��/]!��1��Z:�=�Z�'�L|�vD(�;�$�	:�]��7ؾ�K�ߛ��/�;)GkV��v�[�ػ�hw��|�:3��'G�$q��V��_��т�\��3mўݩE�����>�3;�_X�uM����V�~s#��3��λ�{ �i���!-�Q���C�����b�g�����(z�OW������)6!`����6c���	�R���w��[��u#A,����W$�[��|��bN����G&wk���1�Å��e-jz�x���c�5�+;�+��+�Ѿ��-���.8�Y9Nu�����1����[%�&a���g���E���k������0ah �*�+]P�-� ,s.g��ç�4PB��ҡ�v�bZ�9/�h����ϰ^Y�|��g�������HW��($Y�{R�A}��F#��q��8}ye��1"wA,���ͱe�s4��6Ϲ��8��a��8��Dׇ*/�~����߆~�]���%RO�ٸ�(�4q��AA�L��S�]m��s)�~;	ļ���BU��`��$p�g"P>�X�S��,���i����h�;h�`�W����W1n!O��	bEv����PT����jU��ހV|�8Tf��G	�.��ޘo����wn�$���|Y���}���b{�5�E�H~-ܞ!ϻ�EZ�A���3���-�H/!��,SS�W�3�Y�٪ڧ���h�S��rL�u;�������]	�4@�
A�*����Uq:�&lR}�������(t�$��~|d�B,l4�o��+�2��.��M���N��w՛[>��5�-�b}����j5���e�A�ž�-����b'7`A������n;�����\�x�|R�:z0�~>bЪJن�'`K&"G��C��@l���.-��a~������,��=�)h�xEMb�g�b���2�Of��mR�Z8B�K!���������h�A,b	��P|%:�����3�_S�vx���%�w�J��w�}��Is�1!�遳q�E���(�K:;�����2/�0�r����Q�S!ca ���%b�6��C��Y��]��L��o2�@H[}�ɽ��"lC���Ǟ�m��{��`��h���eXh��aZ`������n���-�)����HIw)����t�4�p�93�9N����g�^��;���m��Q7<i_�Ss�����|����C0/�MNu�[OJut�h���f�7�c7�y�������0����YG-�G����;�V�u�����B�}�Zh�o�wf��j�U�B5��B�t�z����F�q�0FN<�q�&�N�^#�.��r��lJ�h�+:���z*)	b��o��:4�_"����]-s"��c��HW�I�5'�v�t_�c$�����>F��z���M��� �J�.��Vfpu/!#P������Y���k:��Տ�`q���X����Ϧ�W#��U���E�'E־_�f`/Q;Df	b�A�Gc���x�sv�E�������#Be&�H�p*�*�E�ݛh� �,������/W�+�e!)�t�'c���i���&���b���Hs,�DZMH�-A�Q��2�y"g����o�:�RW<s�obޏa�������Ik!Kւ3f ����$�t�.;r�ͨ�{!6�#"�U9Za�T#�rC�.N:1�]1�� XW��͛Hhκ�$�1} � I���<'��)]��:�q:M�mp�t��%"-��A��Z��@���w�=���.�Zԓ"^rC4�͂�Y|j��ߴ���!~)�b��	S�;���b��i���_/ȃX�ܦ2K�Z��s;���F�jU��B�I�+m�R�>ӿB�}��^;;.��
e�~��"Cb�|�l��[�0����4*�1'��Ҏ����B?V�R]�T�ؚ�h�G�x�k4t�Ѩc	M����l�2�p�7�V�Ҝ�Ĕ�iH�j�<����\�U�E���X1�4:&ѩ=�%n#�K|���bӖ��	�'^��)� C�l3e�1�W�3|��OΎyˬ��x�T�A�ѰN�Fm;��5>�4�n\��+3��-�lI�$��{=~b'����ԅ̢��Q�Y;o�A�+���p��1D��N�X�Z�co#�uK�!>d��w�
�( �b�7�1��9D���e�T���yA����0ܩe���їB+��k ��#�f@��Җ��a�Ni�ꢃ���5�X�|$Q()��3�7� V991�ƙ dFma�$rw��Ķ���I^�J�h.ر+F^�1��x���"����Q�B�S�}jFbސ��gYI��Ua'!1�,�{�,��)c�H���	u@�cHV��S��X�lbK��L�#�&�ݮ-v�r1�?M�lM=\ @'bz_��l��P�t�l6Plts�\r4e�
��Z2�RV�n����7,�(čz�Xz73����X�MV�����r��s�>�1��|����k?c+�1��=�ܭ�!�!}�.� V��_������E�v�?�Ĕ4��s���`��;;>
�O�� ���yń�nG{c�ʤ8�*8�Ĝ�3c�=,-���KP���U���{,�[�/����}T��Ov@,`J�|�O�5���s�u?�2�+��4�6=̟k}c��"uNe�Z�����KJ�rB���.����b�بΌ���#�޶t�bK���� F�+�O��0X�Q��4��B�:�(ᴋ���=]����b,�G�i|��{͵�X=ċ��O���я�4r��"�5�NuBA�	�mc�۩�99g�"r��"M���4,�=F �+��1��NVx� ��~�H�햼՝��~�^ ��50�y���٭g�|#�LL( �i�ڠ&?��-�Pj��n���Pľ�q�1h�5Wy<;9R�'b]��^�z�}��Yf%�#���� F9q6��9{��L��V?R���b_����h�"�m�k�/��B�I�1Qjqm��6�.|�>Z5 %���Ve �ޒӴ�3�}]3峍N���:i?���*z<#kT݂s�lĐ������_n�4..T�2N��+�m+f/��U�f��,��~[�>�L��_uR2aAq���&�`Lk�I<�eV�����V��~�����U2�g�o�Y.����]�{���x�������z����hEekE���3�icԍAl `���O��*a[����� �A�����P��'|WEB�"Dn�ǃ�5*�z��gO:}'�ź�/ fa;]��G�m�'2��������SND��QT��@%f|XV�  �~���@�����ݴ&���3^s��	�N�UҠ¿긑z�E�kİ��`s	�p�:HЅ��X��.�A���S���+�N�8�X����I�`T�?7�liT*��,���gRz��8�Kk��A�L���A,�(�s�����5���f��30��z[��]������
l� '�1�ȟ5q(����ʦ��b#��u�؇~�2�)Mr���~Ӑ�AS�u�h����H���؞��(>ZM�1$�����+ �B���s�\qV�XZ8Y��P8�@L���><�մL�����-Y��e4
ڠLL�!^�qC�ЉĐ��6�s�G0��amS杊�X<~ti��;�Z4}�4�;���w@l��ks|x�+�����h��bp�����h��������y�@L��ЭlP�3c�[f��n����ѵ�2,>�'2�Л-?LL�&51�ˬ���i�� [WH7A�3I�Ld�"u�÷� v�L�6�����ز@}�,�'���l�z2d�ZH����gb/$Sh��ҿ�R���=A� 1z��R�d���i�!&k;�Q����؈��v���D���Qjm
��w`@8Xݔ�S�����Z!d�׎�'��n��.�ea�%y���2ｦB>hi!5��)	��\�-��P�U��n�!���>/��&����Wˈ��*�I�͚Kt�_�2��+��	���_U������f�\w0�U/��)�ٝ7U�>_�����.X
;��lLĚ	7������Ej��m˓�9��P���#)�P�;��nf�v�b�U^�U�;Ӽ��.����-hL}�Ť����O��w��*3T4l��v�e'[�[�Z�o�"��.#X:lJ{SZnOQ����`���]���e������Cpwo!�q%����j~��K�s(�t(��>'xg��"9�,oGq�NtA���s���1�;Ef���gi��vf)��������ߞoq�s�$E_�t?m'�`�,[���UWIO�d/m�D��k���������/��+���y�*��k�i9��[�3��Az�X����d�i�.r�����ZoDK��O�"� �INP>C`�7�?N�%)��}½�OK��BG�A��X�fr$,&g5��i!H��bB8M!n�i�[������W��خ�������sXx�>_��,c�6F��8Ҹ��W�Ƹ���q�a�%�p�3��U�!�9�P�:��~n,r�F?]S3�5̖^��7�數�@/��sMht�W�'		I��`�G�hr���p;6��}%��B�R�"���ׂn���.)\��#�Q�]�o��t�t���}�Q��51�z���T>��q���Idv��n��qyTz޷�ҟ��%_�HM5Q�$T����N.�C1/IԲ��	��ਞK��o&n��H������o���9�+$4Ȥ ���K����w��s��8��6�	ﴝ]�%��ԣ߻ΏNO`�"UO/1Q^�yc1���e�L�K��A��/��fӈ!YWK�w�R�첵�J>7�WJ|�>׭%�ZeU���Rh�� �����ԩ-�Rm��>�0��65	D���W��'�Q�Ɓ�t���dc����ŕX�|d}0!�8eC�M�?���2���ۤ��;4z}㶺U�8��Ɨt_��1��h��B�ﻥ�gҬ��Fl�^4~�L9�&e��L�w�mf���q���B�%pG�=ٗΣ��4��5역nG���u�h��b�!{���61���~�o�X8���c�����!;����[�����u�<=�ö&r����1��ٞ.�ay�����~�vj����s��-�*�#�^iͦ5�ů$#sdDUaZΎ{�RZ-��_��C~��l�yծg��}gTg�����\t'�Nv��v/�K�ױ�ڢ��{�罔��fnY*R����=���Y_�U���ʸ�!1.�GCL�)0�?O�AXc�D��������KGZ�:kz�qR��V�-\���ө f�Aأ\���]k��`��(
6d��S(��Y���9�v�
�c#�K���\\�m���@8RPɄ�<3Ĥ͍�<�+؅\o<ˠ�8�L��4��8�bq������ҿu�n�Y\�:�֒�='���&E���0�J�i��Jy\t���}�E�l��\���/�"AL������JE7�m9.�}q�h��X�(iв�4e��?��K�>F�f��$rllt, ��H��ǗvvM������Ml��U$5�''��t����NoX���L��"�DӺb5tҲu����٩�PY��o&�ԼTPs�ǘ���F��f"��}I�Sͷn��r�?���g������J]�7}?�B��̕�i��z�� �ĢR\ \I�����s1+:�~��6ny��7,�d+jZRU��;��,�=G`24_�0#����g^���=^ˋ6��<x��{|aCQ+��8x1��]����j����\�t���Z�㡐��׸��=a��!���n�|z��VG��ov[��#��U��3j��n�_����O�q�zw��Y/ڲU��J��I�e��WՍ�ා>Z�64�,|�GP�4�s�&+���!��<���j|`͇���YH���c��C��u��_u�ɛ���֣���䇮���rkU��Q�ݮ��D�7�B:~��Z��֏OZyn�a�P^_(r`��[���>?P��;g2�!{�;%����NcX�F��>�a����0�N����xF�2��Қv��Q2�\�i�?i��_��,f�/ƥ[��~u&]^���9����YX=\�Ν�Ұ��u�(�0�2Q"B�������v�yJ��)O�Y�9N�p��B2tNz�#a�wQȶ����M"~7��q4pGo�������Ō��P��3k9��v�V���ޡ��@^�klkA�g�l��l^��sŸ�?�Ɖ$z܋=��>���M��� vs�ѯ><�%�En��ܽ�UK�v ������O�0w;}B��vC|�� �?_u+��~�iA�>KĲm�r;�Ż�u��2d�W�������T�����wQ_�̸f�A̵3j��(]�E�lm�:;�B��������B��b���8�e�Z���q�r��ë��b��A8 �y=6�Q�RB�_=�!@0D���[y�G�č��(�)&D�A�>8$b�.�s���^(ͭ K���󊥞�+�/&�Δ]P�v[̕kK&e#�'���F�QzW ֺ���1�V�-�1%7�3>b�	���汦�&��ָX�|n"��d���*&�=_"��M_٦�W ��~�&F7�M�b(֎@\n�(����Ϸ/�X��z�KPi(�`�����!��6�rZFh�F[�<�=3������-��Hi~��a��:tUeJ'�1H���^Qk*�Xms�D~�6#�{���\ذ�]�Y0<Gfl«q������ӌ1�\/�aԯ�6&'�7��`������`)�T����[Q�$b##�R�@�<.v�M���:�z:1b7>̐)]�U�ќyz����]��1�|��IAo�=(��ГA�P�=�*~J�A�[Q����۹b����l|x�CM8~^^qN����ri쫗i���R�}���H(��D+q��
;�B��Ƕل��؊	*IGy��K����a2,�eSzw4�5��uG{l�D�pAY�a�rS(�/�b��K�M�[DE�����R�!��<9��W�	Y��5ͦ@����4+f�_�^�M���+�Ą�jkv����VKV�P�]�� ����=���.�g��i�2-b4�DT����--+���X�OK\@,�MA���4ᝎ���F�˚�� v�m;��:P[���qR��
w�4Ć�n�P'�'�TEu�{L0��Ā�	;�5C�����_%���A���|�uf���C1ake�9���;5��گh�!ůtτǁ�qJ@�9GPU6�� ��mG8{��l�7�� �Ŭ����q��uČ�I�߳|e�X��w4y3�Utb��X�!��#�c�%Ɖ�~�l� �Kɘ͟��7%`$�L�`�x
bޅ�u�#�~�g*��sq��� 6% K��J��W6���V{�?�N���G�^�B̩�ݲ�(bA�!�R����4V�T�[%��)����-����N ZK�Vվ$b;Z�y����p�ݓۦ�?q��؇M_��I�Ȼ��n�:wl��@,�w��ӱ��0�@��Y��Lê��Y�%u��\]!�i]�ăX;��NXm/'q�^���8E�q�"�ZGAy�+���7�s�[����ƌl��0m�x���;5�=t�%��C�2��9V+lv:%�����k��h���g<z�q�w�
�{o��^!#��Dv�
ٛHd��l{E��[�Q���N��s�������|�]O�d�sT����p��d��7�&[m� �I G E5�Ȱ!-���q!�F�(�z��j ���/L�p�K�ت|�M��2VS��r������;w�wZ�v���V+�����(1��K���Q����*�Ի*Q �f����G��"g�>|W��j��/���'m[��<�Njb����4���AO*/W���Xd������R�|(������j@�!��e��l4�APcf���T-�=�ɠܾ;e;/C{���=��.��M
m=7:B8� �޾�C��+��`�R|4^g5g�C:���Z��gAL��_^e�N�i8�u��.w})�Ald�[1@9��f���C=�6���R�ʵo�[k��[]�Ŏ1�W�Q4�,�f9�A�됃�Qw<.�^DC�^Y�-GiK՗�}�+�Zf��[o�
b!\�h�i���l^E�ӧ�,�����nk�4���}s���Ek^<��A�ާn��Tu��<6�ab�.�@i�a�g��U_-��ܗ�1��n��J?d��[d���#��A��Hs1`�f��Cr')?ql�z�]RJ%|Vm��&[�<�A̭���\������)�|(F�����?�q�x��H�y�f)��S�����nE�9�k
#<� G��D*�c�E���oY�����F�� �h�.1W�'>{� �eN@vzG��!��ީO �H�0�$v�chr��"�.�9G�����!����!�,gv1��q6�%0A,6�E:OFH��Y����" 6$5��Iw�����&5��3'{�����4�6���b�A s�=��xMW�F�����)|�
�����\��D��&]�ڙ��RA�&��#3��k�g� A�m�*�������eA�����K�G��GB��3��n�˧�'uMU[(8K˚5��?�dc��e;�A3�兒�;T�;|�8�D� �mK��A�i�:@T���Tb�w�P`��Y�i�_�g]����{E)!�P�lv�GO❹��@�����A���ʚ�}��E��iG��$�z<�"��9b�Y����+}B��L����;�����6�*�R��=a��3�;�M�:N�[�~1�r�V�s�y�ob\��c'�>�GolЫQ�?���X�K�Ufzn����O,�DfKKt����UT{���1��z��5�I!��cxz�%�� Fyٯ�����״S_:�r^��1 �(z�������?	>������̛�w������e\а���in�����2%,�P��bH�BmJ�* �V���a�����F�@��%� �9T%_�{��RS���0l�r!b�'�g�y��6^��B���n1�:��6��%�`�I<����@�ǥV۟�a13�њ`��"�N�Ӌb5=�����P-���Xp��Q�Ur:������5Qr{.��C�T��1�XzS7����z����IG���6<����Ƅ+8oj� ��"���S��f0AL�7� ��A�K\��l��2Rx�#��0b�:��v�N!mv�� ��;��d&q7������Q*�D��d_������a�t#����4ɩ?6�5}�D9:�F��KO`ɮ!��a�|�#g8
"���m�deV�����yKU���l�q6�n��/����?3et��.��M�5^լ���mA*�|��=h��U���d�}�-Y��N��|FtB�T�|�i���*q�/��TzR����&
ŕ�;���t����L\� �;�bW����tlGO$+xR��ߙ}�ޔ�h~�4V� [�ܢj�W�$iBH��{�����{mվ�Wn��S��|8�K�4�U���$�S�3���<�8�qrC�\<�֖����*7�
��}y�ac�C�=��:'�o&�ekm�\4���0
�y)�J���GF��i��P;+��.�d5�3�>J�.Y�/�J����VQ���i���h�7뒓7��Wץ���OrI��]��`DK�N���;qӀ����@@�-��:}ʅ��oR)�k��/d�ÿ���Gt�E�JGJ��3�nҼN5ݭ��b��0���J¾���Akw�A����Ǎ� �^�;���j?�v�u�eC�����y�5��k�MZ�+l-c��E�|K��Q�a�m ��M3V�R���%3��79�k�ۦ,	�d��K�[��������£�:Jn�X�?�89^({�,��ߛ��0�5�%j�^t�R
%�Ӑ���`���,�n�$�-��n@�ۓ�������s���81�#~c^ԘW˝�#hZ�n�D}隩�-��4�&4q>Fm��.���ݚ�m�����9g�lL�� �Q��x��#����z��"��pv�W�����{��kr7׻���LA���f_"7,m�ծS��፸^T��6���S�͒zmP\ [�%:������# ��E]�1,�{{�z���X1���}�ɹ�[5g�g��τT%�.饆���5x^!����H 5"j�R_M4ҳ�|�).!��K��:�0qx�J[#f��:�6�=3�K��|�`��턡'>���Jb����5�d���b�lo�c/9F5�[�69���1'~>�n�� �,�UZ]~�>~�n��w�a�i�k_��sw�W�g+���A�qi;�$�Î	k�R��������ԾR#�E�Q��r�+�yk]L}�c�C�� �1��ZM?��0�ET�a�g�/���0^�t1S�s�Ϋ�2�����q��ޥ]~Q�Zۭ�x�0U1�
��S� ��L�Uc�����ݢ�}��Kl�t��}�Y���O_dj���e&���n�Q.*�	7H>y�e�� �h��m,�fz�o����L��}������9u���tx�2�6�#g��mwz��y���s�,��:����`�v���EE��>I��/C�=O�� �I�a�ɹZu�ǎ����ӷ���9c'��t6�]h��ɿY�I!n"���r�|~��*g�z�7��a�u��������%J�bN�(�_�HѮE�سl���m�Ew�i�
1Ň�`��|���i%ƍ4���R��H�_�_�wdw�e�R�%�PZ#x�����oyE���7f��u�3,���!�;��3��f�W�X���Q��+7����ήKS���Q��G���Gn~������/A�N�Z�y����;�#a�������Kc���3��J^�:����w��{�ݶ������v��*T_Kbc�Z+�/Q�󳽌��v�a@D��d�۝���k������a��B|*�)�E�	}Ȝ�C�n�Z�_5�D�/b_jSTUj9���f�J ����LT.�-�5�r�	ц�S��῱
b��bم�X��vbm+�-x3Q�뱬[O!E���@,�X\r�^����٥���Wѣ��[����`~Aj���b?֏o؍�.�6�U�bp܂��*��X�I��;w�a�mCk��a�/7���~g�7�S��\_���e?ѻ*�bq�W�8��b����h����Ѓ��"tsD�"4�g�jc����+�n����������G�5e�XՉs�T�(�;��8���I� f��V@�u�}IA��S�ʱ ���o��E9�,�'��:Ԭ������kA�I�pcN�"a��*���k�(���;t|�g8amĆ-�&��d�5]ҐV΄���@�j;� �����=cRꅼ��� f�_��#�<��2.f���$S�
bg�%+��z2��u
y�DU�S �+S�y�(�����&os���I�T����~��t�`nN�̡��B��7�(#F-��!m��@�S?��L����Q�+=�v��MZ�Z�*��mw�.�d���_��b%��$jx�O�	���z���@����	���-(���d�
i������"���P��RB6�A�s�y-������Z߰��N� ;Zt]���8�Ӫ]}6�K�
b�%��H�+m��zM1C/O�X9+9�D!�,��W�xCSO?�AƳ$JL`�QR�];���@L����	�kn���HZ����'�T{壾,��0XߨRB QḠuRb���
���q�C����Ʒڤk@Lk��FS4)���~�,U�#/9�-�ue=`k�Gw&ј%���.3Lk'1$�N��ws-� ��gP�{�Ĳc��� b�/VD�ˢ��J�:���@���J�(o����փ��#� F�'_�0�H=�<�Ծ~��.ĄBc���"�*��0�kq����U;5��-1D������ 7_�Қ��~�=��Q��k��z V\���x��jM��ISt[o��Y#���h��2ݓ�pZ�r9�X"���Wl�n
m��̪<�aSX���#'rʴ֫0�Yo1N�����-%#���we:�@f���lH���9D��G*VBU#SP=�T�5=���V)�BC���1���멺���%p��Y+,� �ec����T;C0��K�>�Đ�Ь}3fcT�&�{����˷A,>��.�����v��Ɂ���<�㛆NF8�U��Ԓ����O��Y��jw �%Wx��|��6�j�:	 x2���I�SΎt�D*"|Ě�;^�1yk-������V�2F��N��~`H��� !�WA�=Wrj��,Q���q͒��h�L������5��(i���p��b�=F|b91�,g��&�\���n%N�뀘\	������{��E�
>G�%E��i�&��ꟴtX���<���q�+zB-2� �;�;mz���M��ŘA�[b#i��ލ�o��uDRV�Ca�@��_�Gw��RA��أG���})�5Fa��8n@3Ca�-�K'�+%�������t�6m��Fp��Y�y��-� �D�|Uu��Ϡ;���o�찮�`���sQV4�����5bF���&~�
u�B�v� 6`�I�"��p.��ૡ���8�
����q�<?�[�tr��md��MQ.C�V<7�̈��z&`�K���9�����H��<w���n�RT�s��P�!��シo	�J1/,����XGD�r�t?t#ߺV��� x�I��ϲ��p���&��Ba�ƾXث7��%wc�ꪔ�8;�W�Ъ���o��ܑ��/&5,����AYC����:ln�Xz�!�-G���M,��W���G��X0`w�J��w��o���i�Lf)�F̩�8�8\�'�I�kP�4z�ۭ��ٯ;�L��X6�K�!������>N�9�F���a=��/�������3�)��x����?Ǣ4�/��!Ҵ��n��~�W�x����6���_����4;���9���eg�c��7o!� ��?�[7����a����0[�)Q��:�5j�m���~������uϙu��7�i�h�)��6��)��X�M��t��:�)�\%r�bg�R�&��@��L���̍�©��%���O���K���ۊL
���D7�l���wY�R�D����_v���Y
�
���Sʛ7bEn��8�R�]Q�`E�f�;�_u�U���ׇ�wu����&~�Q��cy�?��]�4�fr�M����T���K\���a�����?�|NuI��X(�kQ�v�@�&z�a�H��b��:!�d b�)�`�a`��M����C8���ڄsk>phAt�,��wG�%�CO@��tGhsL��s-�)�7�>����yec�Z\��f��K4��wP(��additionalMissiles
game
hero
perml00
perml01
W?MzUx�G�I�@����Ka``�����'�~d["�����{�>�����@غ���Rƣn�Y�ް�;}�J׿�L�_���i��Ϳ�V���ow<�n|_ŷܰ��Y�os׍�च�6o�<<����p{ߪЊi�G<�9�}�a! *<:ҷ�}�������[���HET   -   ��<�'�g0��`M<��|`��8a�h�y�^j:;�K��dL����0�����8�?�H���BET   �   =gH=0�� �5���5h���2R�6xexd6�oG�����3�\��)+W�U����<̚W������J��W-W�F��[���ZvBVt�� TSf ҁ\N�4�F:�|ܷ��R���4��L��R���"2jV��1����0-����E��k�jm�ḣ~�+N����'��I�H�u�U�tIS\�4����Y�"1H,�O8��:̓Ė`dEn|�-�d�M�O�;@7������#�j� �ѿ�Jl:��gH_Dނ3�Q��?�`�l�Q�ͣ�<����(�ry�ysy!͹�FaQ�6Kݵ�R�H�R3-�[gH=`����5�g6�X����$���#,�W��0����2d=���e�!ܦ>b	Ér���`~��	R+$	쌫���7�5��&�P�^x��@���9�;R�\I���4R