MPQ    H    h�  h                                                                                 �aI=��	��W�D<�lé��f�f�i���Ue�`��CWF�=M�1'���/�y{�%`��?���Q��KZyNZ����i�"f#�Hae�ψ*Dчxc�X؋�ZG����'�<^�(gcA+�ZS�M|���>B�T�~j�-���K@�����xi��|���8��c��A��9�}P[���.����V=L0ͷh��o$��Ql��ݲ`�1qOjq|�MJ�%��W�fN�'$�V'�I�Yh#�@�[��߽��N� q�7�&;�C��n�a�|3=���#��H�0�'�-���qGVt�)٪��W8�0'���fs~��9��!��L�.���8�����3R6%�R�E��?Ф>T����+����*��ؑ������g��e�NÏ��5]���-C]��/��gw����Bf%�Qɵ����Pqt�<m�BU� ��|Ml�����ڂz��7��%�r�}���B?�M���W����4l������כ��5�G��[��O�.%���ލG��B���/��ՀELG�X�9�Td��õ)v�ř�栻mf7�=�J�y�A��*/��N�O�D-E������"c���'R��z~�^�j/e�u�.���q��Q�0`��,�d�����y<_�qp�Ó8Z�f2��"��Q珅�j8��m�"��8�U]̘+O�����]���� ��R(I׎O��=Ď[���y_I�e��P��ts�xQyIH��kRZ>`�y��K�)������$�aqio�1p@�\_eܽZ��5Wx���.l*��f<��Ũ3,#KkW����؟�p��\gK� 8)���!(�4C��@��2�uA�xL�pCeW)H9�̼��Hs�g7��@�����ӯ։���3>1����jC=�䥟��{Bִ��#�_1�� ɭ���o�n���
D"w�p�/����Ӥ�& �*�9��m�[#�&4ɇ�di�Uk.��ŷA�I$�+�}H�m�?���N������_p����T�Ai��f�o�-�&��O�.�[��_g�|D\���w��=EM�h����_�W�V�2=D�W찻�"X� ٖU���h�5d���Ѯ�������˦90�gwZx���J�'5b�~���07T�;��;�0�|0�ܹ��/7�����W��?y�u��͓�����-�O�@�NF<�M�2։!%"��"���-?v���2�e.av��۹m� O_����,�=�R�*�z��cm�f��}bˢ�T�M�Dk2P�$�s$���;V�d&}a���Y��Y{��Nsx
��}9�6"׊���q��}L���io��͇��E& �稰�:��vq�)%g�GC�6�{2m*�;�������[��)9��1<S�iW&�����E�\�A�;g��Ic6�ܳ�XL�MG�W� �[�0���4�s�N�	��&ET��fSH�s��aȊ�m� 73����V	'j+��%��"��룒�)*̇ �?��x!8�#�0�d�}�f��U�R��F�)�&�}8��>-�b�^+f.r��1�~�;�o?�*6����F�0ݵ��dzr���u6�_ǰ�X#\�:Z���v*\>�1��U
�U���Ko�A<��������C��-g0��we�#�xz�t�wk�{}����8�nD���}Ю�F�jUFU���7����+
��6�d��%`��I-����<HG}ɚ�(��4\���뺣 
�۹�=��KP~��LexŻՍY�&�����*�!�h 1B�PLq%l�m��ǳ�@���<�k��'y��p~49�}Y��C�Hr��/�y�]v�^{�H³�E�'w(�$1$��L�7��qÑ�i�#�]J�^���ߠ�I���K"�m���3А����+���P�U���y�J��ۆ�"D5^��S���-���� ��5�z1�k�iOIhI�A��c�~}6�Z�/�D!��ÿ2(�w/��Y�9���}khEZ�W���}��-��Uϸ��"�~7^yN��+���cs�
ř��ع����Ce^!��^o�;��*�"ʈsw�h�J�!F2O�c�1ݎ��js"@�h/��M�.J���˧������6x�
�E�A��;��ҝ����݋���*5�����f:��&{n�����%g���0o�'��	�,�|��!��Zhe�[��x2�N-�������E��ۖ<)su��Q�	�e�W��o�ц���Q�xs�}��zR~`�hQUG*�������F{t�/��-K�߲��=����Tj�W�`z�7~��Ih�Mz4��oM�t�5M��f`=�\$m˘���KV�e�Q�Ӈ	�3�R������ `׆}����Lz&������=q�-�8)/��q�O��V7m]7���w����%�C�8y�"4�<s�*ݿ�.Ey�J%�6PHn�_'*<�
Y��?�,���p��@�$:���"'��~��A�e$k�Z���;g�EuW�c��H���w�b|��{ĕ�Y��}Q=�ws�d�F�%�[�1$�,�CR�b��imf�=�x^ fg��_�=����J2�.yn�1��rA;�p�s��a�F(�:��B�0Sfo)1��)�Z<K]A�B�E<z	�ͦ�b2
_\؊A��_�ь&P)J�?����F��}�P.�
ObFMN��� ���5K<�,��=�\�м�+m	��5?�#���Z �ֺ��s���"7^��*��B(���H��u�T_�K���Y�⨜G�T2���a��*# ���do��1���H��I�Iټ�S�ZH�8�(�oo4�'f�W��h�#�턉�v ׁC�}ŘM� ;�#��gV兺
��~��$�"�R��O*]	 �p*�lǐ�{�Ź���L��Ӝ�&�k�b�q��<�/���y|��p�z\q��ع�sǻ��%�B�7�l?�h��t��#��}d�囍� ���w5Z��H��D��0�= .���w��~��/2~�G:��=i�:�.;/���P����4a������Ǯ��RuSv||�j�����.U�w�s�G���d��o ��=�
�gi��a��ǃ�[9V�9j�lAs���t����?y"��Y������wO�����Mw]t��yB`ą~�s5-���K8p�)����]�w�����c�~bA�<9,�[m$S. ���">Gh���o�q�Q�Y9�X�9`�!cO�\����%��/�����4�VB��T�H#n��[עx�|����̒D�;��1����"3��%r����"P�~�G��)����`��8��m'�����@��p�k�.��ݳ؈�Ț-3�M��������e��!�����S|�q���c��Y����gyD�K-�i�@�p�%�	��hF�]"���bw'K<���������+'K-Cmf�"��G|��9�~�^����Sp��&)�) #r}(z��@�?�
�������}cl�C��ק��և5K]�V`�O�����oި�f��"�������E�ǖX��DT����p�o�"b� ��H��G��JV��y�gOi����̱j3�D��?��,�LD�|yC���'�z9a����?e%�	q���0p�0[��,����jlyWvyq����fm/y"7@�Q�OC���6�(JP��:�Т�����&D崫R]�{��{��R�~��j~�=�T[��œ���� �j����sl��Q��I�؝k��>�B���Z)���DN��p�a�,���ƃp��_PR���5Rd*�R��*���fW��7�3�{k��.͙|ຸ��3�bKvb�)�\�!�Q�C�1��r!��F��	���W��m9)���7�OHN�<7ު��>���S��1v�OEl>L��dS��ICxo��:
@�vZ�j��#�b�&_M���3�� �X�	}��'�wZ��/Nx+�-�w�n �"Dt|�m����!����m��I��2u}�$ǵf�}�]C�:#�������k��z���zT�A�T�H�
�P�!UO��~����zm|�%%�� ��#�E�0����_F��!�M.:�� e��Ǝ�[��U��Zh��d�.2��]��y��r�ˁ�Ξ��tZ���E$�'�X��9�w�/��T���˱��6�I�`�<�7�is�����Z+cuz���b:��Y��-M��@ډ�<?����T�<�}�rcp�|}�v�5�2$�aq%�6����ٙ�b�,g�̨i]�eO����m�7p���b����o��M*�Bk�)�_U���WJ�q����a��~Yz�{0NV�
=�9��������Eq�H��g��ăQog�"T�E!26�"v:hkv���%�uXC���{m�F�ֈ��D��b�[Y��9��1�>�S��9&�5F�]�$k��lYg�Y�I~@f�.YX'�eG������f��s��eR��N������i{=/S�FQ����ȅ A�[T\3������	��a+�4�)�5����$S��[c#?q(�!S∴�5z0�����}G��P���)�j�C�&�3o�i�:�=q+��Í��yK�������Hn���q�	 ֟I������p�o_"z�[�/�7��[��l�U����|oH6w�=3�3��9���4ǋ�ea�{xu��tA���6�N��:����
����7�j�=���7�H�������d���%��B�#-6R)���Go�Ś?IY�O�y�'��۴?���p=J��Py&�L����9�AܑY��(>��1�B1��q �k�gl�n�3��$<=���� �T��o}TХ���rIc߮���]��{��L�*�%;6\(��$G����K�q�u�iQ�Ћ8�[^1Ѥz6I�r��n6�(�>�����ސ���i#�o5U=��Ԋ|J[����75فS�h��h�9�3.� �����ӟk\WI���A��cs֨6ǭ��ʉ�!��;���>w� XY����E�h ]�W�	���-�Ѝ���"u��^6��Ƀ�+��c��4Zش�q�l=�C��)!0�٘o;�_�e_=�#o��c\ӗ|��O�}1��>����@��/�J�ɰ�#�ZC���@6��N���wLH;�4��=���ؐ��H�Y���(�����
~d��b��߻<os�]'��T	�c��ѱ^&���,e�V�s�P�'���%>� ���(�q�RԅuN
��]Є� ���?ѡ�-ɀ�$�S�8���'z���c�WGrz��_";�t=f�Q5��z�=C�ݵOf�W �N��d��d&���,�t V믈TMgJ_`8�\a���Sǩf�4��î�6�nb�R^���GKy�=�Az6�6nL�=BȻ�����W�3��/_�u�,
���Bmؙ���_��%��@8t�04dF�����3�yH�����n,XP*׀RY�������+K��[\�$��v*���?��o�e�!��Zn�+�V��E�c���������Lk��ׅ�{I�Y%�Q��s|�F�QX�k10�Ϟ�Ӈ-�i�|I�|Nx9	g/9�ŵ
?=�Z�4�+2��yn�2���;�$�s����>3�$p��kS!��1��)0�DK�W�B$�ལ	Â ����_�%A�fV�LG�PT�?U�睖3m N����

lRFh��7&^И�Kwz�G5�W3��l�+��	ʜV��d#j1p��gK�q}��n4��m�7�\��f�$(עL��u��,[�*Z:�c�Z�צ�g�f����#���[�U����C8}|ᶷw�7���C�s!��
s��"��W-D#)�>��*7 ���LjMp�=��)g�f޺�E���!���]i�-����0]���p7�l"=��6� ��ܧ�����w��Yb�6|���/J\t�4?:ɋ��\�Kؔ����G�%i�P�2��?@kV�/���>�}�5a�h�� �5���H�[}D	��������_r�
j^~G� :T`i�s���7�N^d���i4�Xy����<���iC�uN
���j�B��yU'�s��[��`N$� ��/�����i��a�������V=�'�An����j�p0y=��Ԩ5�r��w���rMr���u��BT!~��B-wW�K����d��宂��r���2c��A�w 9��I[H��.;�b�E�B��z)o��Q��o�ӓ;`m1�O�g0���%�Y��9��e�V]<(��#I�8[�������r\����;n�ϴBW��3�^�AF��~1C�j��uY�G���)Ǡ�۱�8p\'>'Å�����g#��
�&� ."�1�.V��V�3Ȅ啈���ޤ���P~-���f������N�"�G�x�UzgԠN]�ay��z{����M]������w���ʸ+4�Ű������	��}m⧀+y|���9�0��������`�|�dc�r�F��^
?;���GI� zl�����E�5�[�QIOA��R���==��ɫq���KS?E�h�X���Tی�+G�=�?��9u�#���%.J���y���[ϑ���kD#.��������{��L4'�7z������e~����/���d�n0V�",9�m�%]yr��qf�����f��T"Ҍ�Q�/�� �̧���]^K���4ׇע�Oc�]�&��ְ�R��W���I=�`[_P��n���x`�rs'��Q��/I>�fk��>����F	)�&ǟ��=�ua���z�p��_��[���b5Mp�׭%*P�fr�b�ș3�\k�z'�4��൏u܎�K1��)�!.�C���Z�ҫ�f�#�&� W�x9DD�̲�H)�7����9������c
ݨ>g����me9C�l��ծ'�q���<#C��A�[�[g��I`X���[� *�w��/	&������ d:���&m*1����s_���V�dSUŭ������#3}~C�5��f��\/oٕ�������i��Ə����H��f�OL��{�%镓Z|:�����LWE������/_bT�����h?x�M5e�����7�U/�!h�1dKh]�~z��uh�퍱�\�\����Z���@�{'뼂����J�$T������B��䵟���7Y�c�g-��u��u��9�=��˔@t-��u@��
<��^����W�����W��v3��2��alK���dQ�vP��<,�t��D4ؗ����L%�m�(�X��bA�5��%�M��Mk�����=�Ur���˃�S&a�zzY�,{ZwN�kG
� ,9�$��@d?� Ffq̱�B�����	oV�"ͽ��E�4�^�>:#(�v�O&%]M�C��{��W�qr����O�[�99 ,1a�Se-,&����dZ����S�g�,�I�j�ܩ��X��G�J�6V)�v��m���N����KVHS�	��B�]Ȁ��Ķ��3V�R��6	�E+x�~�d�(�!�3�������?,��!n���{0m*�ڀ-}�Gg�K����MW��&�	���Qt�:�+��ɍ^~�t*�%���)T�:	c�<���}I��8N�Rw�kj�_}c�,>�Jr}��� �y���U@?&��(o�J������-�ܭ�[���G�}e�\�xp�t������Ǽ��d�3۵G#�XGaj�U����7L�<�wv�/�5d ��ZE��}�Q-����ȯGʇ"���H�j�P���S��M�/�7=偫Pt��L� �K�\Z����P�����bB��vq$8#S��)˩�<�.X��$U�[��j�A}O���*rES���]l'�{����e,��d�(��$�;󓭸?q�y�i�
��^l#^�I?5��f��|�݈)�y�h��AƼ�
:�U� �/"�Jq����5T�/St5���=��Ν� �`��0��ke�I���A�ZcNN$6!��ed�!������w��oYz����@h�PW/�E��9�-����n�t"0��^Q��D�"+_v�c������دg �ǀ$C���!K�WT�;�ػ��ʾ���^뗗�Oo�91Q��`|	@�+0/%��d7��}Z���#�Q|t6�)��;hER|;7�9��q�ӵ��f� 	���Ԃ���N��E3ʢ��ګ�o��'A��	 �B�Gw9KW#�%e�f�n�zBE�{���;�S�L�Z���u�<�����f��0Ѽ�+�����.Iپ�w�z����^�UG�����4�t��u��v$�(\�=ތ-�J�W[wê�k��C�Q�O���t'M��`3�\\�����[��~[�[�É_4��Y�R��7�����������Q"Lpu8ȖF>�6"����.w/�т�Ⱦ�t�mS��ZRW�P�{%#�t8o:�4s�9��"T�N"by�����)sngp�*r�RY~����R���Q�v��$0	;�QR��L���w��e�!��Z)�ӖqKEk��cmw:�����KB���22N|{:�Y#p�Q3� sW@�F-T��21�w�����؋�i�����Ax2Zgj}��P־=��ߏ��2s�>n�S��A;��s4c �|u���-J���S�8N1  �)�Y�K�:^����{_E	�W֧�*_ҷ�A�]���!VP�}?�B&�1@x
���M�
��fF��<��K��mSK�|������R�Q�ǋ|+��	�i�+ �#E�����`>�ij�?cf7�$mk�����(����^uй�-.��zm���{#���w��n�#8����T��}���V�83���EٲY*��;�ή������tRWn�*�j��Yr`��C ������M��9�g������f�E��.��n;]?�"pdVl}	��A@��+ұB�Q�Rr���NbF����/�SB��!�ɦ%\g���o��1d%�o�-\�?��g��I.�Y��}Z���CuR�[w�5��H~�Dd<o���;�ó?�څp����~��-:��i�̜���	������4W� �Z��wy��T�uI.�2��j\����U��as�� ��Tp�� �]S�	�}zi�u�az�ჀC�Vx���nAiK�*d��+CyXT'O��M�w���l�MmG�����B��~���-���K�˗�����I?��m1��I�scO��A�	m9"�H[#�.v�l�Xm�=!ҷy��oU��Q�3n�N�	`Ha7O����%�?s�w�TX��Vx�sJ<�#$q�[M����^��#�H�;)w]���^�3��6|���������T�G�H�)*��V�l8KA�'ys'�7���̮˟&4�����.=!�ݩQo�~2�3܃�#y�}o�O�H�J�4�b��_UމX֚⌘��1�g/���`:�f}[VM��� �]XȚ�-.w�ym�s��
� �������m�a��f|^�1���F�+���IA��; ����r����L?��i�����xl~�i�h��L�>5�袭LR:O�G��D������~�Li���0E)�X�U�Tu.���O�Xn���!���͎��VJ�$'yܾ�F��L`��;D��r��Iį2������'c5Hz��#��c�e�㉃�P�T@����0Q�!,��S�༨y�Jq��ēɗ�f�D"m��Q�/��{ւ����-��ƍ���i�@�5��:t]��5�1�mRYJ�����=y�z[:0_�*��6b���,��s��Q���I��k��>�Z�U��)܇���.��g�a����sLp��_����+��5H�����*��f��z�3�e�kw����ఆR���K��)�I!�*�Cw)�Ga{�F���^����NWZ1f9_��-<H�7T�x�tE�M[��>Ŕ�>�P�ibHG9C�ps��l�j� [�#�Ǐ\s��8�Z�{Ϫ?����L�w��/����m!e ?r ���m��������چ�M���(<8��l��a1}Iא0u��_>;��ٰ!�p���D�����Ȃ@�߱�O���6GX���|���Re燫�E���%�_��%�P��p��ȉ��unl�і4U�Ah��9d��h�9�e����h-��7�۞V!ZI<C�;Ώ'FA߯õ�e��T�����-M�v�|�7��t�"��Ɛ�up�q��8����-��@�_<�|�c$�r\��hDs�2}Uvn,�2Z�ag����iS�1��"��,]@D�o×�[��km�9�Wb������M �dk�e���wtD}���L����a��Yp��{5�N�=
s4�9�ˢכꅏ��}q�:���ƀzۑo�S��Xq�E���d�:��v���%�D�Cv�{�S\�|`��E���[�ya9T_1���S@�.&2����H�I�R[�gM�I����$T�X��%GO�ʥ�5��Ie��*�ȌbN�H���n�1�S����7��{<|���3�=�ǂ	�+S:S������dx�j�T4?�/�!�ؘ���0Hh�zP}Rh��F�P�� ��%9& U�_���"�+ۃ���x�o)k��z�[ӛ�U�᷎�nC�Hz��m��f4�_�l�a�e>+�h��a���}U۠���Qo�~�³gr�H���/�k˾�k=�e�)oxke)t�5M�����^��ߔېܔ��wj&����:7�=��2Lu�J~�d�P}�5�ϸ4�-lw䥖��G%=ߚ��օd����j��js=��OPo�Lv�޻�w������3'���BgZ0q� ~^����70Q<@L��e˧�%�K}J^�T�;r�F���A�]�8{l�ҳ��bq�.({*�$���hE�q�AiG���� ^���muIz,�\g������,��z��C�|Cjݥ^<U�����J�^��5���SO"؋���i-i ��c��x�kҒ�I���A�	�c)��6=��� _�!�G��C�Rw`R�Y)J��;��h��7Wj&�N�C-������"��y^lJ���\+:dzc$E�j��تK��"�KCDq�!fE��K�;lqKۧ��Y�Z�Y���2�5O*"1.����0o@qoL/`f����5��+��$�a�6ɥ�g�-
�;r�۝s�ʰ����w��x��<s���1�D��;��ջ(o)��'��@	;Lʜ�����^�Re��/�ic`_|��6�.[佶�T�'�wȊ�u�����9�h�a�?A����v	��	��.n�z#W`�YDPG({���9l�O mt33�𾼣�c] =y���E��W�2تh�����^��*�w�%��M�Q�`.��\w���b���gʡִQ�d���pR��ہ��6/��׷��l��L�̚�q��qDBB~�)��/Q,��|��4�mξ�5D_Ë$�%�a@8j�!4�M�[uԁi��y>�����Pn��>*�
Yy�K�=�R���鑑f�$�A��,���������e��|o]Z�g�����E�ZcHj4�����W��]��6�{��Y>�Q���s2��Fh�e�}18G�T淇�
�i�J�r)`x�z\g������v=	Y���%.2.��n��@4;c�Eso�=��q��W��Sz�S�Ͷ1,)&	�K��T6��!_	�L(�s��_��gA�t��B@P��:?��x��l`÷a�
���F���-���b*K���PVL�M)��"v(+AC	 W.��3# Q�~޲�b��d�6�x�7���0C���u(�#�2ku�=[�N��� ��3>��]��d�#sT���k��i������	�����-�����J��y{�@��+W�9���2�t���� h$�.��M��J���gg�/�;����	���L;��.� A:]��p�Rl���۬���ᚄ��PR�-�Ϣ�b�Y��$b/ k0�$x��e�\�&��J&��l��%��F�(?W?�ϸ��ק�t�}�漛m�Ӗj�5+irHy��D���n�ؑ���U�����~���:�˗i�Ev?�ȿą��4�5��5���9����uDr��f�jA��!��Ut]sa���4i��;� ���u��84Ii�f�a��`�[��V��;urAd%�߅}��懾ys0	�G�(d�w ��ը�=Mh�3�+%+B��d~�h�-m��K��C������K�h������c
/�A�9���[���.����8\��ԎVo�bQ��4����`#�OV�4��TZ%�E��ңA'KV�,���q#�k4[�E��M������̣��;�r9{�M5[3��;��´"���_�+p�GB�A)Ec����v8&�H'��?�ҁ������z,�Ӑ.Xj��$���Y.�3>S���f:�xG\��Y�ƗL�!<i��\����}�}V0��. g���|D������1�����]��C���w8A6�.q�%�8��5Ӽ�_���m7ۀ1|�u�5��F�Q��پ���ډ`rN�h���j?�T����6�_l��,�Cp�ׇ�H5^�G{hO���ȗ������;>�'g�����E�	X�I{TС�á�4�s$[�����I����3J'p�y�}`���߱��RD�~�^�H��QAM=���@�'��8zj�-����et�ペ컏�A%0L)�,�u9��<My�{~q\J���AfH"�OQ�O%���X�Y
��HmA3☁��{���2]��y��%/R�莻�=��a[0$�e�������g��as��wQ�4�I4+�kw=�>L�8���N)��U��+a�5�p��p�k_�+���25C���c�>*�1�f���|K;3�f.kC�5�j�a૝k�Dv�K�G�)*�\!G4CR�6����Ữ�@k��]W~89z��̨��H�<\7��ȕ�n����B��l.>���<#IIC)Ǭ�X��gb�{�b#�*�w-q��5�5�q��z������2wk:/�����i �V%m`�A����)ڻ�A(�S�ţ�w�o���}�n��+N��6��%�˜Q�돿�9+�fg��IK���O�T��.��?�|0B��\�����E��g����_�f����̝C�I�Pr��Ue��h���d;T�����(�^���r�5J�S�eZ��6�'���j�Z��3T��iЧx��h�)�L�7x��݂)ƫQu�?V����
a�-.E@���<Pw��jj��YA��䦣-�v��w2��iab���G����ѡ�=�U,�+������� 	m�jcgJb�Ql����M�,�k�k�9?����u��*�P`a���Y�_{��N��
��9��������v	Yq��8mE�U7�o�*��/eE�E�6p:�Lv�W�%S\CQ�{6Uݧ�u��c����[�'9oސ1��SqA&m�D�.n��<����sg2I�^ܟ�X�X�G�x~�l5��<��#}y�*~N�:�gs�iS4��x���v���llZ3����	_�+.��ڛj�W:���A�l��?���!�-���0#��P�}��A 3�:��td &/���k��+r+R��Q���jH��xS���p�$�2��I��Pwz�����a�_3�D����*A���;����Uv"�����oY�(�nG�cX��m˙Οx��e2�xf�DtR���gh��� �Z���k�6����j�䍙��/7���A!�e+�d������-:���ԇG���pkS֠�������lu�ۥ|"=��Pji8Lѹ<������@b���䳖��T%FB�q\%ىZǟ�R�#<�ql����ѡ���}E�x�)rzh���k]b �{G�ͳ��"(vlu$X�#�Bq/�*i���ek^�'�KGIIu9W�ȟY��G�S�T���+�@�1Ue���&J��ц2�5J:bS*/3�n��ݺ �����zSk��Iԝ-A�c�6xgT�y�!�̿��w+�YD:�춋�h�%�W��X��$�-��$@["�M�^�%�:ߢ+r�c_���lإO��}gC�_e!��J�6;G*�|���!l�Ti՗�?O��1I��V!@L�8/�E8������Y�ko��e�6�A��1���;��q����_��|�yA�5��񙃞�����ѢU����o��'���	V�����������eS���d^�����I���1�!�����u��N8��P9��qH��\���T&��j�i��z�4��T�FG�+����J�jS#t��b�"�ߞ~�=��@W��#�� v�9@���`��M8�`)��\r}\˄4ѩ�p��Q���?����kR/�ׁྲྀ�%�r0W���LfDi�L􈷬�����$]�/p���]dR�*�mI�=�Vw��q�%YV�8e*4)����x���y��L���^n� *�?{Yt=����Y�\�Ƒ�$&���@��K%�oXe���L2Z��P��'fEa%c#}��4{����1�F8�>8{�$%YYfSQ)��s��F�&N)
1�2ϯ�N��i�~��b�x��g�e�ņ�f=�z�E�O2�n,����r;> Us�a/ղB�����^SR�16x�)���K��;q��ڱ�	�a���CL_HA�kԽ6�P�1t?mߝg�V @h����
;l�F������aw1K(����l�H�¼}�+���	dF!AM#�o�F9&�B���_6Z��*7JƺK;����	(h�64��uP����ȏ;T┋�N!5��S��z#�%��,����u��TM�� u�٨\��}�V�$V���=��W$�7TNp���u_A Cqd�i��MA�U�]Cgª(����k�t�þ��;3-]uFMp�l3&�gQ˹�)��8����0�
� b|�+��\�/[�>�eGM���o\]�@�%�Tǧ �%:�՝#B�?Q2J�`�eΏT}P�����}�5���Hte�D7.�)#ڑ�3���髛R�~���:%�Pi��K�\Q�I��1%4M�3�����:�:�u?֎�I�jҏ!�<�JU�]�s<���o�L�Y ��m	�!��7i�w�ap�+�6�V��֛$A_���ʗ��[y�,SEǍ��=w;<��CoMc�fBL�~�O�-�VK����*6�u�c1�����cũ�A�>9�J[�w.�{��3�,�/IMo��0Q���DU
`� LO�I��T'�%�k'�-��η4V���@s#چ�[ûe��ߖ���G���;;��� U�+13�P��i��O˓�>򏆫�G�us)`�[�L�8G'�k�m�#�П��]�W�.s��ݟJ��4J�3y�<�Y�S�s����O�T2�<���7����|�@@��K-g�u`7��վT�\����T;t]�Q����iw�(��C�@���u�ӗ��7Nem�����u|�)�j�?�a���?�k��W�Mr����xe?L@��x���Q�.lt����D��O�5���BĒOR�d������w�
�����~�ES
ZX�]pT+5s�\㾡��$�����M�3r�J��Iy�\j��?��Sn��w�D�{��9��8A$�6���2'�	z%���e�"��u,x����Y40G��,J��V��y�;q��דJfY�`"�2hQΏS�15O�5p�c����՘\3������ Jv]��y��0Rϕ��r=o�[�O9�����lG��=*qisXrQ �>I��JkR>������)ҩ�ǰ�n�Ka�xA��Ep���_<�a.�5>T�׾�C*���fû��<�3s�k~�J�k���ܟ��Kb)	)E�!���C-����%�|���B��7JKW���9��E�#�H���7�3��X=��"��g�;dw>�[���jiCd$ѥ�\o�b�/��i&#t���x�vS�n���8Z�u{����w���/:�:��cҋ �A�`��m�`e��K���@���.�����㐒�R>�}O�K�&G��Ow��:F��7��f����D�@v�αR�O]?�������S|����7$�����ET��#�_s?h��6E�2㝾�.�+���G�U 
�h�R^d\�ӯh��C*v�^�u�������Z�f�1�+'��4�%C��ST�ϥЂ�V��K�k��;�7jg���]���3�uf���G�E!c-��@@Ƶ4<��«�����v��^������v�i2�"�a]}���w��¬�Xþ,S7l��D�Q����m���i׽br�M�۞�M��ky�1�K�z��J�sa�]Yf�N{뉞NB�D
���9�yz�QWS�1��q���Y�0�o"N͎�E:X�o'�:T�v�.%Γ�C,��{Y8B�B����5�`�[E��9�}�1v��S�Bd&�����"�̈́���g�d�Iꨫ���X�զGŐf�U��OG�~�>��N�����sSo�-��q�'��	3�K@h�	��z+	�L�ʹ��/��7���E?]�8!�Nɴ�/�0�C���R}�	6�<�1�����/�k&JL��U�)�T�+�C��`�e���6��цw����m$��֋�N�#��\(�_����*@��6��{q���XmLU�c���o�Gd�)G��~O�%H1�t���`�e�"�xa��t�T��"�����տ��Ff�	8�j\\(���7]���Wр��d�J��d��.�-� ��
>G�y�+oֻ�G��T#�G���F=�
�PejVL,��|([���I����q�P���=B���q(F4Ք�Z�i�m,<
ø�nGȧ>�;�}@l7
��r5�G� 4]ݜ�{"䘳����a(q�l$����޾�qJF|i=i?��<�^�B�@�Ipf"����<O�bj������������U�\��@��JG�i�M�5ŷ}S\��T6�ퟬ� �I/�A�kHN�I��{A}z.c�uw6�:;�6��!�C���j�w�#Y_Jm�1��h��VW����ʲ-�tF���"a�:^� ��=�+�&c��4Š�Mؠs���
{C�n�!��x�~�;"{Qp�ʏ���OXN���O�$?1dd����@'W�/�D��5���K��h����h6��p��u�G�;�������ެw��4���Pj���m|���t�����;�o�`�'rּ	qPќyg��y�ԻHe����_y`Q�Ҭ|�d5ｬ����>�u��ˈ�4��p��t�Ŗ�l���y[����zY2��O�9G����Kѭᅦ�t)���t�R�ٿ�=�f��;��Wl	��?���^���Aȳ�#Z���M��q`$��\ͣ��?&��ҙ���-����Z��R�,��ϒ�vv�-�����L�ۣ�'{����x���:"/�)�l�E�m�c�뇟���%�j�8`҂4�Aԣ�zA����y4}`�ny�*C��Yo� ��i�����a$�u�������HZ�e�-2JgZZ�%����E��c��x�o	���c�O�CgV{kXYt�Q��ys�y&F޿���1�:�
m�	h�i���h�"x�lqg
��!��=�v�ߠ12�_&nGw��h�;44s���M����	�SW41Q�H)ȟK[w�k6�L�	��@�)�_w�A)��8q�Pp��?A2Z�&*�?���J
�V}F�X�#|�<�hKc�����C�C���ت@+�;	6�&�3#����²����Z�YP7��fSj�ɉ(C�o��u�x������O�i$��S���f��#�Ņǟᘟ�ꔯ�5i��"���#��X~�_R7�v���W�^�q�)��[2 �t朗�M܉��
g���8�r�����Ù���vE]�p��l�.��"	�ف��U���[�E��b���ʴL/��l� �F��y�\����  E��(�%���e�?���SgΪ�H}�I�Լ����5a~WHoSDu䝳�{?����K��v5q~3�l:��i���4Z�:-ۡL��4Ȓ߰�ɟ(����EXu:Z�CM�j��^�W�5Ug�s��������` �2Pd�M���i��a�%C��!V)z(q�.AZ9��;��\q�y�H�f���a�wv���� WM^�u���BӸ~W�-cA�Kb̃P���57�^���Z0Fc�D�A&��9��M[�\�.'���)�:.2t��#�o��BQk��<`ٰ�O�ԉ��N%��Kǈ�;�h�Vɜ��>#���[�QC��='�����Y�Y;Z�};��CB3_6�-q�꓉�	���NG�<I){��w8ܓ�'*��ɹ��C-�7gO�W.�\3������3��W��ŨnK�`��<1��W������:?���I��툶g@R��u�����F���T])�^���qw�/(ʤ6[.a��l�r�ur&pmm����|o���%"�|����j���m�P0.r�]��<?��H�3���l��l�v��uD��=�5R�I�=-�O��X�>�=�/���������7x~E�*�X���T�������_/�����nv	J]g/y�[���}����XZD�z����sP��
υ���'t�z�(�h�ejr܃Pk��/�w��0B3,�����y��qR_��Z��f���">�Q��e��R�~%7�u�7�(���&廁�]�6�BrR�k�����=��[ˏ�������3s���sw�QiI*�k-�>�aQ�&�t)�j��p�)��a܃�fg�pbwX_wlL���c59����*<��f�	�rN�3N��k�+͠N�+R��K+L)`:[!
��C��69�9W�d#���W�w�9�2̞�IH�Jw7�E�E���@�����{�>�K��٬�C��	�A���]�|�1!
#/P3�'��A�Z��5�m���u�w!ߛ/�RUg��Z� ����Tm�[a�(Ǉ��%ڷy���[řV��kկ���}���!`�p�U�H~�����ᬽ�����{�`��j�6�O��YgS��lL|&������8hE���|��_��)���8���A�9G_����tGU���h��zd����jM"�^������������T�Z-�,=�'W���ಱ���aTvn�]�(�� P茕�Kd7�vg�SX+�ᅍu�J#��Rˀ-T��@��e<���U͉ó�مr���<v��2+u�aX#���9��b��s�,�b⨰�%������[,m|,��g�b-i����M���kT�ۣ��8.�C�]�	��.*a0��Y�rj{�z2N}�V
D�)9��@׬=ڏ�L\q8�_.f'�OoB9Z�)+E���8":[>v� %I�C �{�Z#��X��}��P�[ q�9�<1�*S�4�&��R�d����(�c1�g~�IS�ܕ��Xnr�G ɂ���e��R�ف�ŁN8������d�S�V����w�l�G�"�93B�W"��		F+�q�P}��E� �"�?�!ڹm���0��0�%2}#� �7(L���J��A{&e������+ȧꍇL��`淜�ի���M�(\+����5�����WR\_�Hp�����b��}�&L5����U��h�۔�oܟ��fp��ft��B��OB8��zehOQx\EPtP�ݝ7�3��P��![
�D�*j��z��{�7���c�Eћ�pd��b����i�S-=R��`�G6V�����֌��x0��"�����=QxP`�pL�y�7t��Ȧ9��٨�L�=��g�B8��q��@o������@<�41�I�N�G���};#2e6�r�̮�D]XY�{�/4�Q��B_�(lP�$������qe�5i�p)�3�^X���ZYIk�i�m�)�ϳ��}��^��w-{��v��U�t����8J�%�h_�5@UES�y����:�� �,/���k�lI
�A�bc�m36�-v��3!��y�T�Aw�<�Yzz���hgK�W�<��^-��j��PB"ua^�;�0�S+��Tc� -�;�F؛���3΂Cu��!��~@H�;����O�*97�Jg�C��O[�s1Ui�Li@��/d��Б��%ɧ!�g�=�,6ڽ�'&^���;#�y�Dx,��������k1u�UHv��1H*��qj�ƫ�o:��'-1�	�Q��\F�	�e�)��Z�zp�J�gb}� �'+ ۸;�y�uUGl��:ʄy��p3�(M5��K�t��� z�O�JW(G9��͔��t�V��ON��!�=J�^�62wW�$ת�Ɛ�뼠�/c���t���e|Mn̂`c�\(����7W���ǡG�����K��v�Rel؁��@���I���2�L\�J�"��"k�{4�7�/&�>�ӓ�`1vm?f!�����<l%��48[��4�H��-.���}y�;i�X]
nS+*�^�YjC��N\'��?M���n$� ��1-�8r���dPe[��g�Zb^���!EW�?c�Û��]��X��x.���{&�oY���Q�s�wFy�_�A1�^�e྇�F�i����5�x��gV��żD�=�5����2_��nblw-�;��s �������K�dv�S�KI1lp�)���K6v��E���%}	����n_��iADz"Գ�FPKe?|靝���_��r
�
�a"F�e��!�K�}
�!���>�$�3��+r�0	Q���#�������x*��U�5�xo7����/���(����Iu�F��pS��;;�
�w�Gg��@5�Ag#$(��b�@���0�
�E$N��=��ٞ���3~Κn#�e��	zWڼEʱ7�Ŗ��kxo ��U����Mw�s�!gxͺ�l��� V�#!�t/���w�]�Xp�W0l�z2���f�2�̱.�Ӿ�����Bb�m���,�/q����c�4[\S�����e�q%p@���?W-��@���~L}F`���w�G�5�8�Hja*Dбm����/4����Q8�~nKj:[ܪi�p�P-��0��g�b4Cq��Ƽ|�c^��p֮u5���p�jH�@�rYIU��Ys�M��e�UΟ ޡn� :�i!_i4��af�����Vd�:I�AUs�ߖ��CyĄ;&刹�w�0��y�MY�P�<��B�i~'~�-�KuK=s���4��q��Y�����!c;�FAA��94�[�a.b����Ki)�w���oA4�Q)h9�:v;`�`�O����,�%�L��HD94V䄲6*�#�w[9������'|̴F�;&�V�4�x3:<�h��|��l�<�xGs#�)�=��B��8�DT'e�������
Ɵ�����.��ݕ�����3�xF��B��i�L��m��-��r�y�u ��@�u!-�Ns����g�N��{F���RGX�TX���G]�Z���wIWQ�_IQv�q�����M[I��m����u|�"��Hɗ6��5c)�u϶�3�r�����?S����ه�lj����(��8L5�~q�8��O)̢�R&�J��m�ǫ� B�r��E�kLX��TỂ��@���1��8��j����J�My�z�q��8�ױZJD��j��X���f!�����'�Lz�}��'T+e��z�+�`�@i�=�0=��, ��{Sy��Lq��5��f���"��aQ�o�������X��������}��,(��V�X]�]�����REaA��d=eW�[��S�>����I�'��s���Q6�{I��)k��>�ǋ����)�K^�fp���a._���Mop=-P_��:��? 54�b�t�-*���f�w�x3))k����;R@����UK�LS){�F!�\SC�83� Ҳ�/Ԧ	��,�WF$9�X��{&Hp�7@8r���B��گS����>�L��|���C�>V��ŗ�X�e���#���~�l�{�gs�pi����Y��vw|��/�jYpl �Y� ��:��qm1v5���:k�rR��á�J��F82Ț�}��������߳����:�\���&ƶa�����:�O&�"B��2m|�~���u��s<�E�v��w�}_)|��<
���t蝴ܻ�=��SKU6w/h�f�dgW�%R)�yBݩT�ˣ7�?�Z�Bk�'��'��VߛBc��AET���8F
�8�ĕ�{�7 ���s����'u\ ���˻-��`@��R<a&��O����T�
����vZ�I2��saS���X��3I,I�D���ї����S9�mw�3%b�$���8M�:k/=��<��������i��u�aKѽY\T�{��vN�
�B�9��B�D!���qS�������
�o}p:��+E���%jK:ʷ�v.�;%�b�C�f�{Ϝ��x��{:���[�X�9�%1l�S�F�&%������tV����g9*�I ?���XI/�G;!ӥ=�����44���iNS]������uS�i�I��g�C�}��3�<�=��	��+�������({<�鰇}�W?Ӿ�!�D���70��,��}�*��2܂�KX��.&��K1*�_�+,u�"X��[e���3xG�c���d��4ڠJ��s�Y���R�9_D��ut�Ѯ���>'��΁�UGg��֩�oj���"���n�]'�*��)�le�wxW%@tc�;�h��N'��j��o<�x�j�����& 7����Ѷ��dxRG��(Ϥa&-�A|���>G�R���������+���U$�Vo�=��P[̆L�zW���+��1����'˺�9�B�|q �����Т]����< �ո$�����qR�}6�h��r���6f�]�5/{؛���p��-�(g�o$ibe�T��q�nWi3��ZJ�^��J��If -���Z��K���hs�����9]hx��1�U�"����J����ٸ5��S�e��&B�ի  {/���AHk��5I%mpAsk�c��?6)A�l��!ҿ��e�wLu�Y�ʫ�'&�hB6WV�ܵ�u-����5	v"�8^�v��Z�+�[c*���Xؖ0Ԏ�*C0�e!���1�;�kǸ������E����
O�l1�f}��B�@ݾ�/L���k����|����3�65�r墥���;^��	谺N��-I�wM����
��#�m�l���&n��;Ro�_#'��	��x�orh��mJ\e$���UQ˥��"hV�����Qۓ��w�u���`]�Ԡ �+���C���b�t�u����z����EHG������ỬvtM!�*B�O�i=�'�1�TW"`l�Tm��;r�����������M	��`�\�P�˵i��LW��&{�ЪY��dR �܁�S_�y�ף}�؆�L�j]����]$�d/�TV/�����ۿ�{p�m��勡K �wd%*�`8V�T4:�ۣG ?�մ�y*���3z�n�Ɍ*yYe����n�����C$�c������s5 �~��e����Z�J����[E�Ϲc�u}��f�R�����{�[Y��HQ��s���FTR����1Ȟ��s�Eji*�,�^ϕx[�Fg���W��=���V_42S�n}�6��;��bs[��Ճf��?��_1S�`B1�)VK��"@xڂgw	�`I�� �_y�A_J�.FaP&/�?���8_�����Im
l��F
=T����ugKٍ�����9�o��_Y+-Zj	lK?�c#�?��*�����PX�"7{(���ܬ`N(���'u!4����L���Ŏ����I��|i#_YӅ�0���Y��e��ߤ��X�.��F����ժÊ�(0�GW5�������m��� �t��Mǆ� �g�T�'��;Z �����O����ɾ]F�p�$lD�ۘغ�M������ә�ᦻW�bMr4��ħ/l*�o��-�\��Cض���X�n%�ӝ�?b��N7��C}�����Hӂw�5��He�D+���Z�6�J䑉A��,[�~���:�!Li�i��E쿰T����4�o[���������u0����j<Ʀ�߄U	�s��J� ���� �0�o�$[�iOkNa�.V�Ƕ�V��!��KAPͪ��"���ڌy�������
w��K��PMT���vB}R~Bž-Yv|K픃��l�P΃�T����c���A\�e9��X[j��.�\��_P$�7�@8�o��3QD� �6`�0�OBK/�%_�%��(�>���)JV����5=#k�m[t�Z��X0��x��;С�q��9��3b����� ����1S��CG.*�)�����X8�c'�Ъ�>�������r�Z�.�����c��]c3*p	�*!��dO��_��J<�LO��7s��Sް#���@��b=g�jsh#&<������&��P]_���TVw����|��"*�x}S�(�L�6"m�����|%��l�ɲ����{:ゝ��VLr�RΡϲ}?]�����٢~l�[q����sz�5�t��3_�Oc񿢴&��e ��5����H�ʖE$��X�Y�T<��Í�5��<s�x2�E-5��ޯJ�ޢyù�̝��󰲱'{�D���,{�����W	��n'*d�zV�>�B`e`q��I��{à��208�c,[�қ�{y��qH��)gf
T!"t�BQ���B��Eu����k-	���Q�g�!��P�]�������R w<�'z�=���[�oY�Q���=�r�����s���QQUvI Y{k�(`>8N:�\8{)�L����:��aI!�\Tp�_�n��2��5/X���	*�LIfjhя3�k/D���u���9)ܰ�GK��)�z! ��C��.ne��M6`�L�H�VW�j9�B̔boHK�R7{꒕{�y���l�lk>	����%��*C���w*�S����1#��T�U}��kb��)�11�F�N���w�*/kؤ������� �i���m̰���#R��O�-K���ŏ]��!�$y�} E?����&X���e��7ɘ��I��0���J��G���])On���P��7�|(N��N
�09E%��r�A_�J���k�
Fם/�������R#U�]h� �dm`���v���,��*�~0f�?IZP�!�"'9'���V����Tl�� ��T+e�A����V7{���ɭ���ju�ՠ�_<E��!'-��@���<��g�
�@����Ϧn�y,�v��72az'aN����d���T&���j,���fu�+���60mrnqz�b� �,8bM�F�k
���}3K����i�<܄af�Y�U&{|�jN�T�
zy9���bj(�bpqn��$�9���lo����_jQE��瀻T:�4�vI��%?��C��I{
����{�v��q)�[v`f9��1��yS�x-&Y��� �� �`�g���I;�܋��X$QGv�W��s��H����o�Nn2I���TxToS =��䌕�b2�ء�3��XH�	���+����`���Y��x��� ?��v!�δ���0�}�<8�}Y���-�՗�a�`��&��Q�Ɗl�:��+>г�����Vm�G����/
�����T�<tĒ�J�Ms_�{]0IG����s���	�	<)U�h����ao�d�Z����𭖗��6dPre�6xR%�t��G�SS+�ii�F�F�פ���HHj-�H���=7nх��Xz��?d�"��|����<M-s�~�}l�G�0�\���g�nG@����ۑUi=��PV-�L=����kZ���1�v���Ȇ@*�Bn�9q�KQEwǋ�ͩ���<{w����l������}1����rf/!�Q?>]N2�{�'۳�wzxC(b�{$�c���q�2�i��A�5��^ΰ���IIa�l�#��EG����������ݬ��U�1�QN�Jx!
��sE56��S����O��p�2 vRc�R��kyWBI@�A�/cp��6dt��$�!ͭ��
w�3Y�:'좙�h�MW��U{�-�?�ϐ�)"�;^�ѕ&5+��acKs��q��ؑ����rC�Z�!�c6;�;�Mk��`���@�!��8�Oѱ)1����B��@��/�e���}9���J���a6P��Est�e;�|R�z���3h���ee����m=��d�Ӣ��,Ѽ�o��'�F	��H��6[���@e���P��&���ݍs�lܽO�n;��<u�6��̄/�X��tR�^�*��¼�P�ξU}z*��@Y�G�,��|$���_Mt�c����ߊC�=�`�,�NW}���4��!�k�%̳qv��L��M�M`��\��M�p��#�.�=�Cë�7��	R��9���O�*��^�Q���LRb�ȸ�_���>In���*/�^��IC����vm5�5�|�xò��%�h%8Q��4�����s���{y�66��vnɡ"*�mY`�����H�0�$<ܠs�Z����ڨe�v�CGZ�S���}EM�c��� t�����*T��{���Y�ҪQ�?syөF�K����1����'�:d�iE���و�x6ǹg̶���;X=��߱=V2���n��Imf;���s��>�]���	��i�S>�1��)�VSK��7]Z���	���:U�_4V�Az��ԩ�P�?�AC��+5���(�.
'��F%�����+�
/K�J�W,�4�v���E+�/�	��wC�#gP��2f���OR�KN�a�476��[r��ے(�n� Rxu�A���Ώ��"�zS���ĭ����#������G������E���s:�ٔ�����f��G����W�	T@����{�a� �`��UXM����$og.pͺ�~P�V~W��Q,�*=@�'<�]�lCp��l�s?�S��h���$͉�t=��Եb�g��|?/ǿ��Q�H�\I�ؑ�7Ǔa%�?C���?���L|��(�}<Q�e$jӽ
�52�H`��D��-�Fȑe�Z������~�g�:���i�{~u�k�_��Q�49�+�|x��ِ��W�u+�iTj�
𦨅�U�C�s�_0�[�v�%� ��_u�R�ߴ�ij�a\�Q���V�W�Bv^AKG�L�䗍��y�\�1�o΄w'�կ�MO{��ZUB8��~],�-��K󆑃����J�O���k�9c��^Aw�9?`[E��.�<�����c���r�o�Q_���0�`j 7O}6 ����%{C�Ǚ^��:�V�B,a~#F2�[�Ԕ�T�����jG�;�=C��4�E3��ޮ.»����mV��حG�P�)���8\?8m"'��G��#������H���C.߷)݋�E����3e����+�_!d�qp�m��� ��k�k�(W��E��&1���:gQ�$#��A��Hlx�@0l]��{��2w����Y�̊��j��u�#o�m>�p���e|��VJb��@5�+��]凶�YrU���ʰ�?�u��d��ٽ�{l`�����׮�F5#���.(O��3�o�ހ���c��n<���#E�L�X��]T���HP���ݙ�Kʻ v��CJ.�0y�/'ܛϮ�Q�B�D�M/�� �$>�T���z�:'��z���]�ee� ����	��=�H�"03�K,���B��y/�~q��r�fEى"%�Q��%�ri�  ҉�ˏ�N^��F��(���]�S��Sy�R��{�Bg�=[X�[\���T��ؑ���vݴHsDYDQl-YI�4�k�sY>s�\����)�m,��CZN�ad�{��z�p���_( Խ���5*DV�*u�*m#|f/���B�3�J�kj ��q�B���n�&DKN�)���!{��C���,l����ʊ꟣��W�ݱ9Ag�j$H&Ϩ7�����(�;��	Yd'��>$L�rx�j2�CP�+�� �N��Bv#`���$�b	�|�����y��ݾOw2F�/&f4��:�O�j aa�L��mgf���a����c�!��
����]�>w�}�
֐kl�����y	��R���R��f~H�,T-���α���OɌ����R'|�����G���DcE��U�m�A_�8ﲲ]��%7��$���e��3r�Uld7h���d�yӛ�㱯��J���Y��zs
Z�P��5'h�x������T������`�!���;�7�d{����2<UuR��:��1b{-%Ta@��`<;t�Ŧ��+�J瞣T|�v�z2�,�aI���*B������#t,?�ͨApy�=����T�mm?��،b^���G��M�k�h;�7���q����n�	��b(a�m�YRw�{WN.��

u9}U�׽��" q���K5����o�>w����E�A<��,>:@��vd�%��C���{E�ݮU��q����[1�@9�9�1b�|Sbʐ&��55Z�䅯t'�g�o�IVs�E�X��G�1�s���ܿ���*N�'��y!�S��S[�����]���3��3s��s(V	z�U+uK����^Fo��=�3&j?IF�!+���v)�0j{�w�H}����(�D��R�~�&�d��A��8�+y���X��Q�!��PQ�m`�����I,�(/�wC钏��H�_�D��=g��Ȍ����D[U}�G��3so YS�����k���M��ߕ�5�e9��xME�tt�^����й��$۲�0��8%j�zÙ��7����z��lRdnu�W��8�-�X�x"�GG.����'՗��w������[]="��PQ��L����h��9�����Ve�{;�B	΃q����B��F��٤�<�H��ڊ���Y�y!},�v�er!��l8']�N�{�����+�(]��$�M��1�q��i)Gp���^	�"RgvI\Z(�~Q�� ۡ���V���e��!�G��U�|�����J3�2��-z5��SqŐ@���+ q����f�k4E�I[��Ai�rcKH6����!Ȼ�e��w�FY�ʊ�-�h���W�{y��2-�����]"M �^M����+\�@c�܍��،C��D�ZC��!ʁ�d�;��=�e����;T��T�O�˪1��}Ľ@��/��e�xs��2���n]�6k.��OC*;����ǰ�8���qL ����F@� x��#l��Ţ\�qѷ��oK�'^g	����e��6���|�eZ���K%2�z�Ҙ���if����I�*��u&_������E�y���X���+%����Yz�h��;��GJ}�7�b��2,t�����q���=I�'�dW�6w��3�<�����%�L'`�j�M?g`X�\9}��+-ߩ>~N���XÆB�F��R6H��W�Q����
���L�y�ȓ֭�ӱM䗍��z/7[R��r��N�m�-�W�����M%`��8L��4�d��́i�y ���un��*��vY[�;�_�<���3�F$�4�N�i����D�e�4���ZF|a�.(�E�6rcj�B�[����y�����H�{Wg�Y��Q��sT1KF�d�0!J1�Os�v�f����i`��Tb�x��g�[ō�`=�2��<82��n����:!;�C�s�Uչsp���S�u��S���1�ԇ)ƼK�2����ڸJ�	��B���!_�5�A��1�$�:P�"�?-��ni�Ʒ�(
�A�F@�)��B��&KO9����/:�D�r+�%�	��x���#B���m�z�I��Fd����7�	�����v�(�y)[�=uWo~�곆����;���po�?�B���#�2�3B����5U��ᎨW����A��K� ��(��W�_{��!�B҄܍� �l���MH����f�g��&��+��q��w�����b�9]|F�p�kl���(o���ݱ����O��1r�b��2��Ts/"�g�Ք�c"�\�w��l����	�%A�j�
1?����.}���@������5�(CH[K}D���������7���� �~&:,wiz�=a�~�&����,�4���W���Z��AHCu&����5jy����KtU���s�ƫ���&�� Ϯ2Ы��.Zi��)a׷��}^JV7k�<�AF��ߧ��H��y���$��J��wb���J'+MJj��M_�B�Q�~x��-O+/K�@��<����0�J�"��-vcl� A���9�[ 0.=g�F^����or�4QzG� `E0�O�A%�[$W%v	v���uk�V5�����#!�[��B�����z-����;F�7���/�3�*�@�V�Q���u�M��G��	)�7���=R8H�'	��t�C����������C.�����s�{�z3���`>��Zz�̡�(���3���~�J�&�q����ټ�g�����\�d��.�S*r�{}�]�ص��D�wZ��ʐAǖ��nx���1�^Ǥm�^���Bx|��w�HU��������8M\�<��r�����/?S��X�؞�lۂ�e���6	5����),O�'�*.�ޛ���I��#��EZ�lX���T������	p�n����ޕ�Z�&J���y����:�i䴱]�D����4u�_� �$��uc'�V@z�; �x�eV�ރ��F���Uお0.ǯ,П���~yJ��q>	����uf�~"�q�Q��`��Q ���D���[#����[|�����'�]������Rv��]t�=��[7�T��)�s���K08�0s�93Q�%$I0�k���>�����3b)����w1���a���R��p��_c�~�h��5%P�ׅ �*(SfJ��^�B3�'k��B������f� K	r)�^�!��Ct|���҃���,��pWw��9��̊�EH��7񮰕�8P����de@�">?�\����E��C�ִ��SɸI�ȴ�>�#*t���3WN&�!"Ū|�`���Vw���/��;��ʼ� <y����m�����M�KJ{ڣ��<T�Ņ�S�� Zy��}V�d�،ܨ��4ͩ�mm��fK�A�1�g}D�}M˱�O$p�Sά�mD�|۝�~`P�$yAE[I��h�}_:G��m7��@H��%Y�r)�n�OU��h��d#�;�V ������	��4��Z������'�_
�̱��"� Tb���3�ʵ�����˹71�l�?���M�u��Γ�4�l�-���@�<�<r�����ĉ/���G��/�}v{2��aD���i�NV����e,�P���u�x��$�mh0�0�bs�b>�M}Zk�.&�r`&�l�s��J��	pa���Y͸�{2~cNiM�
��9xܱ�w��S�q�z��|�w�o.��͕G�E���6�:���vp]%5��Cs[�{�#1�I?��l1��'�	[��9y�1��S=<&��`�Љq�̇��gjB�Iq;	܁�X�%�G�����#��ؿEd�|�N�<���.�RS�����XaĎ�y3.���(�	���+P�f�<����|��c����3?��!F�P��w:0E����x}���#�ϗ\h@��|"&�:iռ�u�� �+�xM��:v�L���^x���-�.k��ֲ2�*��C:�_U.��Rk�"SO�i������U�,�Ǩ o{m���%R����l3˻�*�:�e�A{xH��ttQ��Ɉ���M*�<[�ۍn�0I6jc�����7$���O����-d�#��2�y�US�-�i�s��G�������B-��dޚ��V����=�n�PLO�L�[�#�C�4�I�l�³�̒��l�B�&�q���-�G����\<q:̸��J�3+�B=�}'?v�Ϸr�҆��QX]D�G{i�³=�P�Y�(X��$zƑ����q�-i��
��N�^D5}� IW'`�ٽ� ��Ք��@?�0\���kU�"�]�J���W5,SLH�{���� l���)~k�R(Iv\�A�D�c&�D6�:��=�	!��%���lw}�@Y�z���zh��W�u���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��z ��UWPdHh1�7�fWAl\o�婶Ej���(1j�Dd
��	Z]����;���4U�1�m�v��}������/;���ƾm3ң(�И����Ir:^���-���a�]���LEp�
O&J:��=�Ş�ѡ=	m�grI�3SZʸ彌��}�����]�˝��}}8@�Pr9D��j(.�!\�#��Z��q���~�j?k�ŉ���P��ՙgZ�LQ̡_�qްj^�=z(�&�]��z�.Be��k������s($jt�&a@���#8_W3�����)!�ns�om����u�Q����M`�,�L Ѐ��������5qc�g��6���M�a!h�E������'/����^���b?�պ�F�ۋ�	�4a~U��R't�,�Q!ym�����B(�84�����]�Ɖ>��(䙎x���l�F$�MF�!���|�R��ۑ�ܯ��JsY ���1߿�B;��y��3��� ,`9��-���L�4�%#����I�����z������9B@�I#+4���0�z¢ �m!ۆ�#��P�/Ea/B G�~T�e��������̽\�o�J�����p'� ��i�N�*�}�� ��A7��.{��G�K�c�W�di�����[;K����Ck:�D��L���ۙ��1�'�vP�s���O{C���'�!�|?Tu�[��^� �P��u�e��}BRA�f��`�;�gƘ��Z�b��Bx�����_�V��(�[�o�%I���aC�h�I�l��3b��~�\�adũBj�ܩxuչ^�Q���|�^8B<����{"զo���:�,��^���CJ0p�_��"2d����Y��ܫ���0�N���E���_� �/��3��	��?��J����,���y�K��S:�J��WA�V�6U_�<��16"�s�wlA$W�Iá�l�
��m_pZ:d~����#)9�s��fL�l_PP����	}���Ɗ��'Ƣ�9�r+~.$�ZМ���n�<Ǝ��jI������ ��$����o]�Th�eC��$���.��� ��E<�$� ����Uzz<�[�(t�P�$�q���q��e��THHЯ)z� ��D��<K�+4�@���'�qo"��ԛ��R�X�i̑M��:���͚6�^.e��{N|ů�Y}��TaΓ[�`4���w?��6N�<3�j�`#���]��B�I��B���� Q
���zˬT��u%�����#�����~:��U����w���uh�:z��G�;F,�"O�NQ�܉��< g�+ \��D$�\��}Ē�Omb�TZ���a�:�)�9���c\P��_%�����^���s�e�\()�m_n�{E�:�z ��K���@�gɷ�aS�����oxL�������<���+�U�/�ߞ��QzVX�5����j��=j3_�K��G�jg��M��&���Ѯ�._8KMj�%"�6_|�w�ĕ���0sηfPȼ@��	�(�H�c�?��R�ķk{i�?�V|\�5m�0O���޴�ֳ�{c����<�k��l��.+%:�'w0.@"OZ�xߋ��d�k�q�����|r�E ی��0xuo�'�H
w#.i�fh��dK��Z�E"�
�������~��ɫ����7�{b�� x��,�9
M�Y��$�vzqx��kO��cT��#�,�9�w=S�����@�����t���J>&���I��J���M���)�^^�k2�Θۓe������ �E�8�.�X�L�%��������-���F
�cKr��}����:�'��}˭��fr��53��~	���t��K:@$�L��L<m��+�A��4U�Y.��p����[��d����aj��"�|�ֆ�9���&�������U"6O��a����o3y�0���;�Iu<��&�/�B
 ��t�H�*��I�j;������!�^HL�(��a�V��H�1m��^���9�N��=H��Ԭ~���C�4�z��ݑ���pv�l�]�1:`��-S��W��5)IX����S�!A.��\I�'�B�]���t��Pc<���m8@�V�m!��zW�~Cr[��B��Y�����QV�n;�hDh�����l�%*&Q��󣡺�(�k��Y|���s}S��.�s���T�B����	7
!f��$��}��_BN�TOr+�N"n�W�X��tʠ
)��oM�WbT���Vd����B��W��\:I>����|G�1U]���dId�w�	e���a^���)�@�&I1�p�v�(
���#9��3�����zP��*XЃ�#�cl���_����w��]��^�̴���$&���SS�=���<��	8t�rt!�S�%����2׷9�����o��?@��=rd|&��e�K�#� ̢����իĐ��;Pq��xZ(4��L0�q�^s��=E��&(���nҙ�K�O�k�������s�t�5h&�i���8� �W~����w!�6us�G���1Š�(���MK�]��X���ҥ��'9�q..]�7ٻ�M����Q�q�o�P�'����Ɩ��?5��1����wX4=U��'oBF,W�y����fx N[��j�4T>���ef��G�������q�����F�ŀӖ�_R�����2��z�i��U�s�p6�γʿ��[iM����E��`-�����^s�`��	�i�a��`hz?�:ٔ�Bk�T#�Z���(�z�χ����������B+������T���a�Q�W�g6^�xzP��&X�# ~��i}�k*���A�AB�.�n�����WPOVit�K��;��ú#��C���D�X����A�$5v '��P�����/C�����'�T �F7:^�|�P���u� o��^Ak��D��"d���ץ��/���A��L�*x�@����y�e���=�[��\Qk�%T2b�����3�JI�j�^2<�j�������ڒ���Gw~u�4�^����)�I����ǣ��~"��Ы�����^��C��yp٥|�m5��Z	DY��ͫ8;�0Q�
��1���ȅ�׺�>2�0��JtJ$���xu"���F�Y�>��J3W��\V�f_N�����3�w�$B���h.l��э��_�N/dJ����I�9ȥ�����l
��['��9)ݞ0�Ƶjb'Q�9�_�~y�����q�@�޸wƹK�����E&�G�d �)�����B��zenE�$��� ��.� @�EG������h��z��q[7���;Ӹ���˿����?ǿcH�8zö�σ��'$>+}xԟS^�|$1�4+����F�BXo���`�b,���LyD�fZ�,EL@.�����&�D%,��*�s�����{3y|4�.�m����@�}�_���J)-?�{�F ^v�yh'�L�U����3��<��U��2�y�W~�o×�U�)�׻']�&AԵ/��F��3��1G|M�|%Ó���<��(]�ZQ/�(�4ǥ��	� ����	�t\�l�<	f��3��1��&���*����	j��N���ӚZ��%�&���Vb�p��{��樱��L�w� *E�!���l�wh�d5���޽{�u��^4���#Z��d�$rJ���+huѽ��+�a'���9B�L����(��JDꆯЏ\\B�������Q��e亗7�B�-L��<�g(@��q��M2q/����Iȇ�6-��:a����_���q�����:CcV�1��K��L1�Y�s����U�/;�/wu�X�J���K^�S�*kĝ��\Z��%��f�1�X�}���ƤI+t������v%�¾�[z��4�D�9GX��T7�H*�����^o�wd!c�����-�ax�����Q�蟐P�ٝ)D�;���x4�����}��sfC �ǒ�i�����s�b��*h"��E��2 f�2K��jx ���&� �aZm೿�8��C<���"�Ѝ����j��� K嘙�R�`��)��p�Xc���E�R�T_�^�e�g�G.�t��+G�� ,���(�It}e_�rTg�*lJ�˹���ЩcA+
�v��tO��AY��ـz)PjԞzr̰ AS�A��`.��: ��)�WƳi� X��qP;��$�n�3C�N�D�{7�-dR��F�GKF'���P���:/�C��~���H��"T˝�q}^w�wP|�u	;�Av鉪y>���jM�3&�b���L��vZ��xx��v�!�ZH���y�[U�N<^�%�����MF�>^IzLڈ)��ѕۥ�2�i��ʩa���KYu���^U���A>�t�1i��IO"+T����N�V7^q�MC���pӰ��A�E-8Y�2F��80\1�=1�c-�� ���_�вݕ0J�iq��s�y����iCJ���W�=9VS��_�����D�w�$m*��wL3l�s����_��ydU8��]i��yiS9��<�vl����4����ݩ��� x�'��9�s�~H��nӊW!��rq���$�׫�u��1T��Ү7 m��������*�ze�Ƞ$l�/�+��.�΢ +(E�Y#�6�Ts�`z�P[Am�f�@�GBT�����7�n�jH�0�z��vߚ�F�R$�+
��Ԋ
�Ǹl��H/����#�X:nI��[Mb�0Լ�RyZ�f��E�-.\cÏ�+8�oi�f�s������X{�FK|?y�.HwQ~R@�nh_��E)x${�*� i����Mڌ�ޙU�᫖�t0���j��U�0<�y�������b�DU�b��'��&��/L���M��c{G�D������<�]]�/�(F4Қ�t=�j^V	�Q�ʡ�
<�9��~�ζ�T���_��4����	���N9|۾)�Z 6^�F��g�۹r{QR¨�������t��lRL�hW=5``���@𽦀��`�𙵰�ſ���~�/o�Jg{�+3E���bY��~����P	\��Y�3�&J��/���\mt��~�F����Ű�����\�8c����(�q�A�2��V���\I{�6��ESz�"�_e��q*g�{��CN�[�|�QKP�_L<ZZ�������Z�D/�XX��H��#pK	��5��K��\%~�%i3fs�X�L�}'I�r�BI6�
�:@�s�H%�m��抷�o�����^�q�!���j��kBĢ
Vca3���	-��J�����QKCA�����ʥ�ƀg����ݞi-T}�Of���]Ț�/K.�M��*i~��K��!	fR�XK��kxG����T��jwa�8a�jĳ8Į$�����6��:i���������8R�����X~�H�#wj����RQ�w_ח.^)gwg�r:�!����\8�,Hj�˳�bth���Y��g���lUB6�^������AV���t:����Kkȃ�1�rΩ�/�HiA�ؽ�PJq��`����������5����Қ�W��� �(�[���0�<�;��ɬmr(,&�&��6跙(,�M
z�ur���%�1n�cD����0B�+����6\�=�X�1yLPN��1���d g�]33vs)�w.�Ut��.v��8!��`��éS)j����1=�p@cn�t�M��56�ȗ��婊�����s{�����k���#6����Hr��g!�쐉~]1���}��1�խ�L�ΚX]�B�JӍ���s����"�������T������]�(X"v�U/���.��7CQ����x�<�O�c���Λ��D��me�-(7(]Y<2_}��k���R�>���s�D�c���3ֽһ������ ��{J�o�V��k���b�]���=��uU4�L{��A2���@������Kn�.;cp��=Y����{�i���� @��<�8֕�q�R��j3���ŔY��0�8��5����Ě ;P�R��W��Jd؁PK�֬��~͞Zc��%���47�8��0�O�y�m�:P~άp��Q�
�>�]��<�pg�n�y���WK{K�ܪ�zF|S<�T�K�����]q�7fq�`h��W��SP��]W��tiGdol�-� �n_��`f�5��A�4Q��?����Ed�-d(�ZC-�՛�L����Y	s����}��=Gck]BF�X5�skoϹXY6��/o��U+�Jp��𗹽d���"!�KQ�n�����x��,�&:%�����2�"d������o�n#�S�އ�z�I�0���'$i[t���v@�r ڎ�g�ߕ���r8�e+r�!��Z��t����"_#�&������Z�D�g�	df�[o���="�U��r�4���ߌ�|O�����o�ڀtE���O}� ���I��
��|o��!b��U���9�"%I7`&vI�if���+z�p�#�#��l$���6�޻���wk,0���=�#�n�J��u�ץ4Ы��L�>4+�0��U~�¤��!�_��Bz�kv;�\������StK�3�/��_ X���m�����X.4;��/�T������m��+R])��h�R����;r����S��v#v���Ux�5>����h+Ǳ���N_҃�o� 5�[�Č�Gm>��A#�pP�Ko�?���9���Tx)��P�f3��D	e����[��KG�J)*�.�)���n��6��e*��*z��7��6�u?*���T���W�P��O�4f�LSzmp�?���D���&|`�^��t�v���SL.����Ǯ޴�M��x��ɵ���e�J^�����j��Y�TCe��
����e�V�r���/I f�?�[B�53�x���EB���X��L��ɣO �o%�qZ���n���ZY�J;g��g���dv�Ri��hU�ۏ�(3��Z�e{��x�l3����#��|��0%ìH( ��W�8_#́��&B���5��Y�oF6�G%e�E�oɧ���#whS��=�h�c[�h�\l�A��5�� P�?���h=Jw	��h[�?��u��b
l���5�3v;��hÁt�3�� $fY�x�����C56���U��3_�������>_�̅r'h����O�sI��=��t:V<z�a��t��܈���z�����H��S�v�'L���v0|^�!_6�u�-.6fݻWSP:���×��r_�v��z[v�ˈ��	����Є�Kq��H=�HdC3I�a��s�G7��!���O�b��W�\��*0<�	�2yXb��_o�%n�
Rw��i�?��*X� �`[+<��\��{p��!V��"w�Ȥ|%<6�0�����Q��`Y�����)(J�����;�ދ�|?�QKF���l\#'*��qC++��i,�0��'�~�&�O�Z��^8<\٥@�+z̚�¸�}t�I<j���-�FpH:8�ͮ]�܀�Þb)�K,�C�s���]��
ט�|���ߏ��`n�O�S.l��U�C5�C���!�B�/ߜ[�;�1�^p ��Ix�zcޟ��!Ǒl��~Zp�]P�FWx�"༹�[���*�f��
�G���a]���Fۢ{+G[�X��w�m�c5�A�>���G��1�f)�r��m�!�2.`��k���<�2M�d�Y�z��M�ۈc6m�K.2n �?�T�>��zGA��������_�+s)ƞ��_�T|ouYgG��}L4�gl���͏!�_�݋]T�~:� �����~����:����!F��f@��h�r:?���L��%BD��������%���C�b�×�>���,؀�a�M�&��tՇ=�eK�!/�-Ep	�F���\'b��C���*���ݳ�����R("��X=0��b��6��| t~@��$�P�n�JhS���봸]a+;S@�t0�T9J��ļ�P�aEˊNMZ�-]xk>��w�NΉk����L0[5 �F�wc]9Gd��6�v:�ץ�(3�|G�A�p��3�c�"�}�g���(t��=}s~@p�2�!��!�a,e��ૹ�=����Jy$4��e���B/���CD�{%�n$�E��>��C�i^�y���,����"�$�8��٧��n�A����~Yg��k��� �6"���;�BÈ��f�:�"�~��IcH�w��K1�(���y��y��˟7_P��>����+����V��=�o��m��j�%,��&2�4��/!�U�rjοw�vKM��L ��2�����Dyq��uߌ?<��!4����kS����Y���@Z����1�� 
d�i[���Gd�?Y�`���j+č���R3��k4����@��(�l����Ñ@a��kY\3��*k�ݦ�D�V��[`N�/t@?�%e*?���J�1�y�4��{�uF�@�wAM�͖���D��&	h�l��^)�b�M�h�KZ@	��q�
�����;�=9X�x"/b��9~�'�M�0�2�R+����e�=N�I����f�{�n�=�3�� ���G8�ߝIN�Ш3yK�`����Լ���-I����% )-�����,�u�Ms��j�~3��V }:�1�y7��L|��Fu@�:R�MG���F 7O�&�д\�hjgk74�߳�N\�,�}�''OE�7T�7"��\/�Đ)�l��^u\(�L7��r�6B�K�����)a!�n����"(z�8�#z�f��?�ś9D~����G� ��d;T��^�U�W��(cݲi���s.5����y�Є;jE�K[C���%g��>D��8���O��	8�-4jsc���.�|�1�O=��m����>�h��r	���Hsd��R옓ď-2i�<pVT�=5ESr'�����x֋�zcb����k���l\��kJj(�0\[O2�<x�����kŹ�uOd~|���E�N��Æ�xM�>���
O�i��ҞZ�[�E���
Ws�9�}@W[v�������7̄�D���v,]�"M�{��o�$��bq���C����F�v+,g��OJ�}��㪆r���-��{Y�>��j�!̍J�$��%�7�¤<�6��k
�����ķ����^���B���Xğ,%����uhԭm�7��3���|xPrX�%��MQ:�-Q�>�h��r���0>~�z�L��N�:ڝ��$�L����ޔ����1󇇁б��=���2�G�aB^*"q�~��hz9�ۿ&gr���%�-0�OΒ|a�c:��63Q9,��7);�Y&<�����zc�3� Ѽ�W+eHv���!� ;x#A���]�6�Ln��s��V� �H܎Umh����ھ9s	�^��|������n�Xٿ���0<"]�Um/݃C4�\�����]6	2'��Uj�<(,��2|���í�,��;���LZ	�U�N�k����Z����z_�乫���e{9���ǋVD�?N�� sW�KNqh�t�5�4��D��1���|�̓A�Zj���{�� lJ�C�+������a���̎ڗ�x���IJ�c��O=\���2��͂��d9�ݑ�����۠G(���q�ι2����t�I�k�6c�@:�V�X_�qq^�Ҷ/Q(C����0"�K���L�6��9�u0h�e4/��6X������CK=����ǝ,�\ِf%@�f'w�X-�K}ە��wWI�@��n��'os%3�Ꚏ��S�6�8g}��t ��c��U/xf��[%c�F�3�-�A������YQ�]�����}�zl'�r@��,G����}�T�f�g��Q�c���m���P/*5����K��;�f�%�KV3dx{İ�P(?��X�aY�M��k28x<x��Eġz�\�Ω;���'W嗄4R�=��`�h�Y�׵�����RCY_�G^�߶g�i�3�������,|s��g�Nt����{}g�SXl	,[��ӆ�O�A����8�tn�@��?2�����*�/z�A��|�b�Ƞ�y�/�P��ʯ�i�Գ��_��<"�Z��(�]�ɝyp$:�vwm�$,ڍy�Zo�6���(<"�M����ŵGO�e^Dc���������2!��q�e�jP*˂e�[�kД���3*[�ܫ�y�	��b��Կ:|!��`@�v���"j_��e��$Yn��M��	6Iq�R���X ��{ЦC�EU.�@$τ3	�6��hg�uH�n�g�[��8�1R�#�����W��d����]������a�`�o"Ӯ5��]a�7cˈ��]��N"*�/�-{.v�V7wP�@���p��O������\6FD+(�ev�P7\P�<�/�	��ȠQ��"�y��D���xS��y���&�$��������V�P>���b���	��)�����I�������^Ͽ
����v��b
Qpój=�R���x��5���UK�
��m�
�l�)�c��R.�3�N��Ȗ�����я
�j^ҟ�Q� ��R�"��y݌d����:�/n�Ro<�����|F��l<w0q��yҒ>:J��nQ=�&>C!�pgS1|y��-���K���.C0SC�T���?�71�~G7%�`��'.S�w��ĥ��#d#-�!Dn��`�1���q�u%pQ��������-FYV���H��Τ�d��_�׷����q0�kz�5�gM��%���Y@���6�3�����=�q��z.���sn+���{�6��4&�ͳ�62K׈���y�f!�nW��SH͟���_���ȳ	�i�ɻ�(@��74���Q��К��Q�ș�Ց�Z��@%"��v��]�3�AZ��lg0��f�.�oK)���"3���4G�zӓTC|I��[o���t�s��5� b�wI�,E
i%�|�I�!��6dF�]���V�v7YYI��@����A����#  $�]�j�?��4)�;�PJ0;zjу�#f1���Vu/l�4���E��>���0	�#U2Վ�ء/!W���v�k*�n���o³�eχ����3�?}X�-����҆����;�M��$<��ס��ߋ�)7.h�ɽ�
 MrC~��ʽT�*��v�EU,Ok>�Z����P-��σ�͎�Yދ���ci>��#��P9%�oɠ3�2�}9hCB��'��usݚO��\(e+)�z�.��/��+*2�%���U�ɮ����'e^�O*.�G7O��6��1?^F9�oj�9��W{UB�����L8�pm$�?� �D6�q�Z�j�5���ڍ�)Lb��0���l*�j�����n�O��^5k�<,�j@��󈶗�䖦�잋�t������G �����4�i��x�D�Ev ���̀~�}�� 8��%;6��#i��wZ��H;d͛a����[y�����D(��Z�Q8���:lg�^�头W��0��dhU������78
���r�BH&ƴif�Y��{Fj˳%�y��o}>�D�)��N[S,P��*k[�\ o�E����o, ���?n�hq�	��C[�^��)�����l]ˤ5F]v�b�h�7�����47�Y:���_�����5Iß�r��.�gUx�1�ސ5,�� *m'�
���)s�����=�DnQv3�8a���{��2�r����3����[;`�7{�vdc��q��#�.��B���g:i�������&�1vE�[*Eӈ��h��и�q����|_H:}J@ԅn��{e���q��&#2��nbޫ���*d�2̍��f��b=�<oE�nY�w�D��9�*�﨏>�<'mۯۇ��wY��ѐw�{�|�U��d7/d��Q +�����)���\n��ȯ޿?�\hQg��l��#[h�%H�+s�,�2Z�[����D���ӭ]8p���Y�#+�[ưv.�}�#�<m�!7�F$xC8���]�ɔ��!�)W5�w�sL2����w�\�̣����B��Qw`"�i��B��|��w&7C�ɑ�U*�����Ї����]1H��p� R�}]lzj �$9� V~���]ĕ�F�tU��b��4��^*C���n
R��δ����mF�N+�QX��	w�����]Ano	�O�bE���CJ3�&gm6r5����I�Ō��2�9�>[��%��<B�m� �2"|�?�&>�ӂG5p����)��_U~�]oV�d/�T5B�u��G*�Lvj��,s�t�N!KI����T�8.�Բ���3j�2�&����$s!z+f��`�IFr�~��W+�ٳ��2����ɭ�Y!-�� G/f��6�`3��G�MO^>��ջ�U�U��-�̎�z�.�3�vb�#C�]��^�ך<���+?���¯@�0ϟb�Hǝ�Bt��Yg���_O���C����l�u_��@��[����J|�ʼ�Ma���N�)�-.�r�w�A���*Γ��[iu^����c���d�������(g�cG�%Rp6m�c����1s�����t���=��#~���pDߕ�+��̃a�=s�Q��m$�=<)�ǭJ�f��haD�M����!/V�S�w]�{���$D"�E��O-4t��i��E��5͆���h$�b�ɍs��P��_9�~����Z3�4�6���YnBwm�˚Bs����~�čc��>��@ܯ�1�ح��yKf��Ӧ)PP�V�����y���m�ͻ1أ���!�"j��<��tC2%5��6�����j�Q�wJ��v���)tV <V-2Ք�~�nD�B�lD�s*���յ�����5�~V��YS�(��E�ݷ&1��4I~�D���;G�Y:H/���+�c�c��3ʛ4}i�<���t���6�w�@����jT35%��(��k�D������NP�*@sX�e��X�f71G���h��{^4�G7��+}Z�Ipޣ=��Z�h��X� ����R�K���Tw@���z��S�9I�^x�ճ������dbM��5��eL�N�9���}��$i���g3�tk��2����N Y�3-��`/F��+��~IdQI��� ��u��t����u1�q�Bꮨ����
=�:��-q����~��ut�:ХG)�%F��ZO���h
m��9g�kh	���
i\"�`}PLzOyM�T�Yѡ̴���"�)ޡI�:�\\y몑�.���ר���Y��)�JFn=��Fh�z�E�W�%��s?K�튫�����º�H��H���K�LU�������z��4�b@�5����.�vdj?m�Kr��+�P�6��Zڮ<�����8��=j�ϗу|�*�]�ġ#�����r���ΐ	��pH'{ �K�R�,���7�i?��V�[w5���[���(��YU�?��c������k )�l��7c�'*0:15O�,Qx��L=J�k���)����Px|�=�Eֆwv�x������k
��iJ����:���E�
lP�$1a��~�U�\�"�7�����у���,��-M��ܚ�$cS?q#���~b�(���*f�,����S&��ٶ�w���>��YpK����>��{�U��Ju���Y�f�vN�jd=k�N��L�@�������ћ����Xx�&%�b��)� ����O���0�:r��\р�g:��3�ݴ��|r5��?�Y~������t$:*��ȊLH
��'a��D\��?퇵���i������8��av��"%�����98�0&�I
fQ��a��O��a����r3�����l�;%�<M"�����Ρ. �_H���P$;���T���o�����~*pH���o>ygi�����S�%�����h�\�u"�%�iA@`����ɹ&���Z��,G��%�R��m
��V��4����A&-��*��E���(w�ٙdV'L#;.�h�Ή�7ƙQ�ڣ3�c(�f��kb��P��}�4��%���W+�>��Bus)����
3�Z�v��}m6�B a9O��+Nt�W9%��F)8
;�ho�Mz�'��r�DdN���kW>U�\Zh���9����1甸��d��p	���������x�.#g��S1&�v�w:`5��;W,�� ���������5��/g�����_ѐI��]� r)�'��&g�e��=���Ξ�	
M�r�=S7��:���$��K�ζ(| �z'@�s�rvam�G����#�$C̴�}�0�B�g���b�x�VP_*�����Z����^@?q;�^��=��&:U{�aY���!�|k����Lvs%�t�֯&�$�f�8��WPͮ���^!I�:s�ͻ�W�-Ųl��q�M��C�i�ɀ��-�G<���q 3��I�|�g?Mx���o���M+�',�R��}��!�-?`�������G74�b�U=�'�Y,)V�y�A��_K<�ݛ´�4f�H�/�`ƆP;��5��X�Ic���F���ӨX�R)B�ێ���L�{��s6��`'�����m	:����׌!`քK-�E��)�@��E2��V��s��4Gz����f�B};�#�%�z�ᤇ*D��e�M�����B=:���TY������ceڽ�n/�
�H�_�X�M6 ��ui�*�V�ݩ�A�Br.x�������W��,i^��{.;ĺu��ChFDSQ���$�v����'��PP�JD�A��C�=���Mᕹ,�TR�l���^�@�P�Ϫu!��zigA=mʪ ;���C�����A����s6���x�OF�Ⱥ;�p��^��[��Kc��%������8��MI!�ň�o�����yh���(�h$?����ur��^��ſj����dY���"2�;������5^f�C'��pkq+�?s�l�Y�\��0#�A���B���}��"��B��ݜ��J����74X�󘻠�Х�J�PW�.VZMt_����W`�ȖwI>h$�-6þ�ql�z�2w_m�dt��3� �9Z9y����li���q��Eu�pϓ����'��h9!e�~KfV�^��k��	�˶D�G��ؘ��$� ������l�h��e��=$��g��6.Ӛ RlWE�S=��:e�z�2�[��r��.���eY��=L�>�I�Q8YHm��z/��!�����+Q��Ա�m���/��qW̢>X"�X�Aߡ'��b�Z���ya2uf��E��.�K��������s�
���7a{�]^|m2.�@6�j_d�4�+O�)�p{}8� 0�m͋q�kwlU�іK��"��ڜA�y`8<�j����U;1����'(��&���/3��{���
6Gj�����SU!<&"]Co/��4��ށd���D	e`����<~ᅞsΝ����֖��o�c�w	��N��7���Z��-�v���^��pj{�ݰ�C���|`�2&F�sI���h�+�5�)�Scٽ�����b�������vU��zJ��+���M;�3M����W.&����lJV��"K�\�տ��d0��#ŷ��Ɇ������N�1(���q�2C�q��X�I�W6������+�_�Yq������3Cu�v'�K7>@LbP����H�����/IcX��M�פK�����c��W�\�*)%s�$f���X �'}.��Y-�I�����r��+P%f"��-̝�Fx��UB�E-c��2Ѳ#KF|�	6�c�˧�fw-ԡl�rS,��Q�Y�����/m'�p����a̞P�}��ifUI}���.ٖd4uT��t	�*pa���X��3yf��K)|'x�'ݗ�����T�a�C_�Q0s8���N���tm��HB:�<���f��xR�S�s�)%�1��Dj�#Q�R�Ҡ_�K�^0� gw�
�F�l=8/�,�_���)*t��E�`��g�!'l���?�"�A���H�Lta�	��;R�����P�/M۳A�Z�����Ē�d��$���#��y�������Ǩ(����ŝ#������mt�,����gk6/��(/�"M�y�\�vZ_���p�c����PyA�r i�%5O�D�����P��ض��������3�ܞ=4�\N���y���!�Q�`W쩺_Mj��X�c�w1�nÆ�M�3�6��@�%�b��\��)X�{Ã���С��	��F��60ś:�H��kgh�`��XG1��:�d��� ��TFU�U�s]C�ƞ�ۥ��Č���"������������[�V]�:Y"��x/��].��7*?(�S�8��"tOd���I�қ�L�D�eɑ7B�<���|&%�s�?(?���D��ˮv֤���Wޞ�r�m"vG�eV,-��Fb�����<����v�jC��y�R�!��:1���`��p�= �J�mZ�h�d�|��{G�X/����vOiR�di3\S���5��wR���C���2��R[ �R_��L�d?�|�Q���ͥH˟x�_���R���p0D�y8�:��Ȭ��Q��>�'$����g&��y�'���K��ʁb�S��wT�T{'`�
�5�)�7�6�`�2l^��S7���$h˥��d��F-�O�n���`��	�<'9�(5$Q�� �����Y�-y
!�:�;�W�!���w� ��JC�	l̤d�k�͕m�%5��R�p�O�Y�h��SY�R�Y�����:����\������in��w�N�t�A8;&����t�2�ȸ����y��nʙ�S0>��Yʟwj�Ȧ��ib1����D@����M������ۧ�X��ȌJ�(ɅZ��S}"N��k�fX�Z<±g#0�f�,o�M��j�"�7·m��4z��&a|<������o��t.P�� 5�I�
��|�+�!i�2�X�p@���t�7�j�I�>n��x.��Ú*°#�-�$�A����`��iw�n�*��0.���ք�#ʖ��ͻu���4W��x>>{[0�A?U����!j[����k�(:�ÿ��F��z�#�:H��u�X��l�q�)�$U��߿;�1�{U=�a��T(�sV�F!Ҋ٨��ϝt� �
 ,�^~��p~y�V��c\���EWU4uk�x�'a��&�wT/����n��ç�GC�����l!�<:u�]dy/	}42�ԧ��v�	^vR���<T��� � �Vן�g�p�<R�	��N���F�Z`����N�eB1�;�{�*�<���7cT�k��Z��w+thw��5���,yN������t���8;.C��o�o�JǇ�+��E�-�LFƏ86U���q��-��J�J���\�xd��fi��hl���B�i��#����(k2�q��2\ĳ���WIsI68�/�s���}_�;'q�+:���wC�[=�ܥ^K��	L��B�>���!����/b�JX�p�0l�Kii�Е󭝫�2\���%l�f���XYi�}����H	I�7���P����7%_R[�F����C��*���V��F5�ʍ	$�3�Onc��)�D--D���@5o��Q�OS�{3�(ol�&�M��wL���}c�f"$ǽ��ُO���v���*�@��)���B�f���K5�x����D���
%a�γ�X�8$�ڕ�M�ƍA�z�UD��(Fw�ChXR�+�O�Vt�����$R�7�_7T	^���g�Ƶ��w������,�����t��
��6kg��l������<���RA�q�a�t�(%������J��	�L/&��AɆ���N�%O�ZWY�JΕ�ճRk���t�Q�("���I����"*�mҔG,������6HHb(h��Mp2��զt�U��:@c��O�I�x�����^3�Ɲs�ϑ�P����)��ĸ����3�����du��\*ώj��k�!Bmp`���MGja9ܑ���Ј�n<�M0��6u����X��3��Bf{�����p#�l�g�߿f6�2j�Hҵ�g�D�����1�����������].�.�o]<_@���T����"�C�I�괛o�4ok]��"�Ɩ/��5."�d7�%θ�6�꜋-O=\��B
��' DW.�e"Vi7���<���58��L�!���%d�D�_��$���g��>C�P-}�F4+@4�VE\�Kh�b.F��52���Օ��|�CZ���f�k��� �C�"��뎏�po�N=����F���a�v}�\�6='A�������RHI35�t��=8��Y8���	�Ƶ�$�D ���R{l�%;�d8�A�a�F�����2�񙶤(5�� �0��y�X:��b����Q��[>oV�����6g�fay������Ky���n�Sop�T<�J����R���7�a�`����6eS��7ؽw �ԕ�d�$-��n���`�oŅ��k򡞪QFGt�KVӛ�|F-r�A��j�t���z��J����Ѻ�:~��̝�
k�����5KCQ�#�/�AYlfG�]��K:�����m8�m>�07҅��nWMC�'U��:q�&���:��2��F��p�n���S�v'��{ܟ�����c�i�<&�AK@|;`Fc���A���T�q����e�Z����KU"����D{�_LZU5�g\�fO�ow��G�z"_���F+�4s�r�?�?|u��wOo�it����	� �I	�
��|�S2!�*ub���	�kւ�7���I�� ���
���:�#2�r$Y4�֖6#�tf��g[�˜�0g\`�/Ft#C�(��H1u[� 40��q�Y>���05�>U���+W!`�����kַm��)P�_�Mϳ��Γ���H4�XF��*���~|���2�;2^D�J�4�w��;�܋)c�+h.��67>r�z��O�֫�vMU��E>#ԟ��`��Ө���������g��� ��G>Al#e��PeKouu#�^Jh9�y����I�U���Ӝ��eW���&lN�hG���,*^㋉�#~���Ӗv8e��r*�.�7{0�6HK?�Ã����e?�W'�n���6�Ld/�m�x�?�	�D⥩����оm��K��9#�L�1�Z�I��A���)"�A��{��^��h�j����w��5ˎ�����'��F�׏�� ���h�!�ǉxW�E�(�Q�ͬa�)� d�5%�Y�'�=�6kZ�,�;� ��ǰ���&T��%��l���;�(���ZRO�?�1l�?6gt�����܆2��ٮ��h����8����ᙕB�2Q���YOx�F��Q%ŏ���do)��p\�ƃG�SX^]���~[�4\���q �9 ��'?��h��]	-�[����3���wl	��5rȭv�3oh#���?��`XY�8���{I�gV�5u���F�Z0��]6F��^�,��'�T{�(�s�m�I=Y��J~��?a}�/�*�^�_�J`���.�����ㅾv�heׁ���>�.�v���o�:;�����ҟvDX[֖R���k�lT���qa�èQPH��R��u�1����X��}���R�_��Jb
US���3*�H�x�����b�,�oq�n�w�YC����*�����S�<.���[~���E��w��|��Tɐ����QLb<�ф��)����I��q[H���)?JJpQ�
���>#��ܢ�+�+A�,I� އQBÆ߄����;8����Q+� ��"�j}��<�2vM�F�Xq8���]<���#S4)�4��2�s��* ڲ�#{����y�����`�)B��ڲ�(���y�C~����)�eq������1t�;p`�.���z�&�K^�̄w~�D.]p�lF��ا�����_��
�h��BF
�o�����/�F;o�+��KX�N�wY ��1�AǬ�{!q��o�	�Ҵ�mbu���~���p�8%�2�򌑹��&ښ��{�mp�2��?��>^XGa�.�l�	��h_�}�J��pwTa�;un�GV��L"��Ǹ�� �<!w���=��T�������0��$����X+"~!��mfm"�uD*r����#����BT�^
�7���@�ߣ%<[ ���h���/M{.-K�H��A9��i���-��⚦�����b�ECI
Պy��͡�W�����M�B��0{�b��I�I5yt�fu���=ݪP1�݆��Z��|@Q����]�J(qG�Jaa�{N���-�X���PwC�k��&�?][�+ڦr�c���dL��°�7~�(�k�G^�pb$G�4c7���u ��W�t3+�=ݷ�~g�pp������av,H�}�#�n�=h��s/��wA������W�E�{/��ܣH6{�1u$p��EW�*Yմ�Gi��	�����a$L���$�4&�90��]Q���~��&��g�`�Y6�A��$��B#q��ƻĤ�h~�8�c��e�p⯈F���=Ey�U�����P�h5⮨܋_4�Bw��y�m���P��yaj��V�|�2Q�{Z�����jm>�wv2�v�U4U1� �C2M�*J�Dٵw�gE䌟C�s��/��Ul	�a��Y��Mqٌ	31>��`�	��~��D~Gģ9Yf���4]�+$*�CQ3@�O4)�Q�h�ˈ�����m#��@�����3a����;@�=�DT> �N��@��e�'��2?@1�����^S{
��s�����u�-S��O���]�hFk6�,K/���~��K�P��>�� ������*�9u��x������<���D��3߆aЋe��{N@�ǯ,�����WP����l�+�)�r�?��NL�Q3��`[�-���EIQ�2�= ����e+���u]R���������Ͷ(�:�e:����Hr�*��u���:��4GU��Fd��O(���}BȖ�g��h��H�|��\N��}�>O��+TR�������rܤ)
��1�\�l>�Z���U͖"���� n<)���n麢�r>�z8�=�.��[޶�K՛�w�(� �o������Cot3�����UD�5a^�� Q���#5S���0��jkQ^K��0�=�w��ni��t]��恷9�8S�:j�Ϸ�C'�|6�����ͩ��h@���2�x��	��HӼG�w}RL����)�i���V���5�s��rM<��=o��<Oc� ��t�kL�Fl�h'c�?�@70f��O�ax�M�Yk%���/^��P�|MC�E8�Ȇ#��x��_��
�w�i�A����^���;EK��
�xV����H�����?��N�7,����M�Qt,���ME�4��$qO*���H�T�J��J�,�8ѯ4��|�#D������&I��]�>^v�ˁh2J!M�Ӆu�"e ���Xkj�`�$E��z_��$�}3��F�X$�z%��� ,��a��e�Z�<|��`�r����,�i:�y,W��ȳr��k�~ANɇ�<� /�::�J��.�Lt%��c�Z�ۅ���I�ᄨ�~��"g��
a�B$"���~9��S&ǆ�4���YO.˝a���@�3���=��;/ι<����9���z�N 1a��[0H���pY;�����O
��rLΙ����V��H<+�m��J�1o9��Ƣu*v��C���{B$�R�r��?��p��$��K�M�I��S�����+�N��*G􋉕Af�����_[ъ;$��"ա��q��smp�JV�w}���4ɶ����)�P�!ʆ̣H�3�?��VM�m;�qh��O����]H�Q����F�(����U�6N|}H;ܾ:l����$�B]H����
Y���\ 6}�!B�BJO��XNZ��W�TtجM
azo�#������;d+"��z�ZW���\r���9��0�1�m@�|Vd�uQ	��x���P�>�߾T`���H1�8�vU�,`���Ơ����6�Ќ��냡л'���U�G�ڔAK�����]�����-�Q&���y=���t,�	p�er���Sv���$� *��q�޶s&� ��@�2r����-�d�D��#;0<��]��v���f��5=�PE���* Z`�+̄~�q!�^�V.=} o&`6%�G_ԙQ��އ�k��B�2�s�z t1&��IL�{8)�W��逼g�!/��s,�5��;����R�W�#M�:w���f��Xo�-�R>sqf�L�o쵻M�{M8"�a��Z3F,'�2������G�b?F��i�U�w�4�~�U#��'���,��y� ��E�8���"�4����˪�,Tʥ+���ۙ��/2�G�F*5z�� �R���4�Pܲ:x�'�sj��W�@)��w�����}�`<	{-$W��c�H8��A�
�݉��zw�A�̒�B��#��D�˸zE/�P>������HwoBc׉�� �T�`'�OU���%���3׏���Q�Ӱu ���i���*E�+�0�Az�k.c�J����*W���i�hĮ<�I;.iK�[c.C��D������!�\~VTp�';O�P�\��'U�C?q��*������T8��~_�^$�`Pɧ�u���� �tA���F�@���_�҆��Y�gUQ�������xf���Q�։�֊[k[��%���)�`�kJvIG���[3Ѣ�t����ĩN�?�#�u�gr^"���P
Oс�[��ͣ��F"���W_�/�I^>��C~Lpf����d����Y�:�pW�0��i�
d��/]�#P��v��hW�݂�PJ:�*����Zw��~��v&JJRhW��8V@��_��w�40pꭡw/��$z��$X�l��$��>�_��d�R��*����º9 F���blB7��|��P5��ֳ#��Tp'�O�9Ƿ~�(=��Dc�������*�-	��>Uh��� �'���{o�W�'e���$�h��8�P.9Nn x�cExͲîB�[z���[o��sSĲ�G��#�$u���?�Hӛ�zU���	�_\+�����y��I�l���
g~qX�uR��Pwbd�i�	+�yG�f�8�EE,.).��1PT�|�	��;s�B}��t�{:7�|l{�.`
��N@���_�m��QM�)eT�{#X� ���ͱk�Q=CU���k"����:��"���Zy�R%��ѥ��hhU�����'N�&yY*/ٮK�����0:2GP�q���s��8_<'v]�/6R4���AW����	�M�N�<A���ky��C͎�#JޖԴ}�I�<	���N杫���Z�v��zP�22h���{�AШ韞Ǆq��X�̑Y0n㤲_hDdN5-��9My��y�Τ��j�@��&���\YwJ4�8+�nV���O��N?�%H�=!N�*o�`��J|T �A\z�1�+lؤ��ŝqG�oa�e}�t�(x=�q�[2��Ť��I ��6e�Dr�L�_�wq7���(��C�D��i�=K�_�Li����<��./�g;�/�|�X�8�����K���bN��A�\�8�%qf ��XF��}r�����Ic��"��࿛%3?���lJ��qla�� e�N��7|p1`xį�Jc��&-�>��"<�lQ[Đ�����	N�s� G7����*�}0^Jf{Jl�����<G�ۋ髚-�*V�|�V���"f�K(xTP�I/��>`a�rp��;�8��t<��Z�Ѝ΢+�j��V�RIW��WK�������R�W_$� ^ێgd@�DUcQ)��K,UZ��`y�t��S�F��g2��l�BM�+�����Ac:���Dt��y>��3M�^�i�v�p/3%�A�B<����
�!��1�@�&�	��k�_���~U�S){(z����ɪ|��`
m?�,�!'�3z�6�(UGhM��i��a�	
��g!c��V���Z��m��KO!�*�ϾظP{M܂�s���P��j��3#�����B3%ϻ��8��!���`�>a�`D_jX-P�~O��]��niN�M���6�q�/����M���{���~���Z��g�6V�} �0Hfg�
Q�֊H1�Bb�
�^ɏ�zO�;_�]�l���f������(",4��B�!wj�A��]�7$"#��/��.���7�͸�Uy�	��OJb���ъ�U�ZDD��e��H7�g�<_�l��M��Y։�ǚ�r�D�c��=�J޵8��_��S�h�V����8	�b���b§�k��W�P����]ϸs��m�����4p<��=&?1�S���)�ʧ�#r�y����"��A�R��13Bwnš�h��|��)Ö�;��Q�; h��R�!ʷ2�d廢�p�3�G͋uJ��Ĥ��P��.0*}y�d�:�Vˬ��aQv>�7N���	�gU�y�m����K�Ǿ�g�S�.�T	_�M�\����j�17�`��:D��S��؊xԥA�)d܌�-�N]n�`��*�"l����Q�κ��}���7-OW��9�a�1�x�C�������p�'���J�k
���t5�c��U��qpY��D�j�U�����v �:��ʌ�]F�x��n���4����NC&爥�'�2�%,�E�����nn�vS�A���9��[�����iH��n�@I�x�_�Լ���}d־��Ȳ���2�ZH�����G",��׷�A�Z���gI�<f��Mo����N"̄O�S{84 ӌdE|bȝ��oA/�trt~�) !�I�j�
b�|�a�!O�1��6�֌���M�7�h�I��[�9��ǵ
�C�#_˕$&�W��u�������0T��Ѽ�h#pz��w%Mu���4=(-�V�>�v�0"�UUkk�1��!й��~k�I�iL�¬6.Ϡ2�� [��u�XX�}���g�:Q�e�>;ӊ�i���0���{�Xf�)�W`h;&���r<�f��p�c�iv0�lU��y>����̱�{��Ճ�$?����;���w�"��bf�}�y��@�у�0�JW�b�Y��a���N|S-l�*-�_w�
]��)�n8][�l�ڕՍc��d���������:(��XG�L�pq���Vc�V`茏c����t�l�=,'*~�iwp��p����a%���PL����=����*�>��f!Mctǘ�]��ԉ�/q!_��u	{��$EEEFR�(�.�fiM`�`>��0c����$�1�(\�������~H_��:����#6����3��7+�Cc}��&�h�pW��vR�~iL��m:�?�L�D�=O����(�~���#�L�����?޾� ���SAI��y%U�^�V��V�jV�R�^Έ����7R5�/�׸|��y� ��e���-�?(xA��E�[���*�VVO ��4%Q�'��i��Z��:;1���q`ܒ��`��g@��7ç�X (}�Z;�����l=�NQ�������F��:X������Cu�8)�e��]�B�kN��^GY��+F@1d%�-`�	<o��Ł*��m�BS�>b�2�[�o�\��H�����# Zjb?�%h��	�fS[����Z�>dls�a5�rv�J�hM�����
�\Yдr�u���t�5��������kS�瀐�$��V5�'2=U��	�s��=Q�=��%D�
�aG�젙����>�?7�2��}�1e����av��s��S��H�.����0:ܷá��ļC�vn2x[@�v����������q�y�R*SH�Ѱ�-�ԛ�,�Qv��g���|�P�Nab�7Q���*�}���<E�b�Io��Jno�w�F���vw*⾑�*��<�#��Es!�<&����w���|o��ɺ�DzhZQ��}��9�e�)�e!�J�[q��W?��XQUP���#�޳�;��+��,,3�ޱ������dF�i�,8����o��+�5ɰC�}�ʶ<4���F��%8V]�v���q�)�
�ͣ0sbzM�=(�T(�"����T�ߙ/`�g��Ւ����M�iCh��x��~ߦÇ䅕x1�lQp����S�ez�{ �uh[�6��~d��]Z�GF�����Թ����q΋��b
h�3���z���Fe�+r]X���wC���O�A���%r��噵;�<=(m�|�Ϡ+p�Ţ�z2WM����z�P���R�m��2�e�?C�>�z4G���V���H@_k�;3�y��N.T�T�u�B�G �L���yX؊��!!De�'%T=A����楩e�Ȳ��2}��+!P��fW���tr}l��C��o#��߱��-��/rߍ�(�Z���6����M��F��Ց'����y-��Pjn�Ɉ�bDȸC�-��4[K�����Y����%0e��b$, ǳ�t������5��N�ɇ�޾��`@�/�^M�JV�t��a�]NWc�-��A�Lw�3؉u 
�)�F[�7��cg�Qd6��ԭ���`(=o=GH+ap��\�h�c�����SM� �t�+�=��~Q��p��ԕ�c�h�a`T�ʧ⫃8+=��]nY1��0t>sИ�7��o��/lv'�Mj�{o��$���E�����i�wi��0�[^��P&�l��$�9ɣ�p�xNM���l~�V��5��
�6l,�N�WB����p���l��~��c�����b�r{.��yam^˩�WP�B�H��ϥ����c;�����7[xj��I�f��2{�lĎ�_�njWCw�jv#�IY ��2+8���rD���QX��Ɉ�����Q��?��ы�Ol��Y)�7�*�3�1��
���@��n}cG.��Yx�q+N�W�yL�3�4�k撕
��U��i�sS@����5��3���t��g�LD��_¥&N�@Ɏ�e��p�܉O1ݙ����_{t�gV���v0�Wu޹�)�0�>h0U�Vr��,Z�(�cK�J�h:dj������^9�Ux������5�qU���z�/t�9�e�.=Nj1��������
A�W��A�M��.2�)f�Nv��3CN�`=5�R�BIz�j��f� s�7�2����u6��� ��J� ��:��M��S�r�㔝�uJ�:��G��FΫsO�K���"��� g5�>b�f~�\xq�}f�OO!;T<���"�R��n#)�pg��]\��E��|x̀\Ƕ��oʳ)k�Xn��b��:�z�b�-݃����L/�C������n
 �.�*질�̝Un��QEݼ��;����5�2�������j�fYK%����ь��k�ӮRƪ���8=�j�nbϭ��|�G�����ͻ���=�H�&�ba�	�H=�!�R6$���iU8&V^i�5�i���9�Tz��b����c�8^��*�k���l����4u4#0�^O|��xA|�Sa	k�a�y�w|���E���.x�>��vZ
Yvoi���(�,�%Z�E��
�1��rG�9e�L��\��xq�7�����*�;��,��AM�I����$�)Tqy���S���Ǻ���,�j�B����ѝ�|�����o�5��� >H1˫�J�F��/>��a����PkԎh���@��[�����������J\X�%5�d�?�x�w�_�O#c�f�F�Krbݏ�^:,G��t�r31r��O��~��K�V��
	o:d�{��*�L���Mg��Fwb������������LjN� aL�"����8�9N��&q�����O�[�a�E��*Z�3��겧U�;�0�<��c<I��%i �T��JH 3����;�d���Q����L8�9}�GVxEHf�m29�ۅ�9�����v�	`�m�es�|����� �p��¢��@��L��p�S�c�����\���$�ui�A��j��d8�	+�%���ѡ�����mZ�V��ҷ07�`�E}��z��4����$Ȥ) �Vw��;e�0hh����t����Q`�J����(�<J��X��.�}�(j�$���՟�Վ��B�	��ܠ
����ƪ�}�z�Bp/�O�C�NĒaW�jؖ��
�	to��9�f���dU6��]�W��s\\ ީCRh�o�17y����cd	���C���(�7�~	9�11vN�v?zy��n�0��|���f���i�UV��eG��I?@�D�P�����g7]'��yz����&�G\��=[���	ZS8r��S��=��$��ҹ��V��x�z���@��rƁ�ח���0�#%#*��D��⿷�gĲfVgc�P�����`�ZJت̮X1q��T^Uc�=g��&�a��#���<�q��k	bN�w�su�ut0&�4_�/>8�L�W�����U�!�o�s����qw��+��AM-�Y����с��N��GqPڙi<����Mȧ<��������A'|gI��~�q��?���o��%�4$qU�̚'Q�,y�y��4���<⁧��4�������֜ ����� �|BFx�����Ry�	��Iܜ�c�Q�s��y��kv�*��轡Ɖ]6��'y5`&��-N�B�y$	����+u��Ñ�D'�z!6ٶ�sB���#X�E�ud%z/Pʇz|چ1����r2��B�g�8�BT�b�9����H�	o�Z�z��!���}P  �i_|n*/eF�-�>A�$.��4�d����W�
iV2y�&ڗ;XEY����C���D�W��$õ�Ƅf�C�'%�P�d�C�	�����	MT��4(=�^?P�u`�q�ʅvA���p�5�hv������i=�ϰ�5�@�.�)x�Eb�{�1;����+[���B%���Ӟ�U��Iq�� ���L���V`�����c�)�u�=�^L�����+�n�SA�'�1"����p��^hdCw@�p�u������Y�Y6�۫,�0s#�4�J�:���i�` ܸ�����RpJ��@�Ӈ�������� J�J4�eWx�V�O�_0k.�.i�w��Z$$"~�;�l"Õ�R�V_��Rdl���T��P��9�}X�ӏpll���f��1���E:�$Y'��9q�q~���g>������� з�Gݫ��~���i�? ��J�`�A�heЂI$C������.#YD ���E��Q�m�T��czc�[� (��W��sF�۾���ǡd�H�U�z���qq�	�'+�[���7�?��L�����
XߡwĘbN���31y��yf<qvE/m�.S9ޏ����&K����s���J
�{�y�|V:.?��(��@�eD_��F�{g�)ϳO{ͤq �����18��A�Uh��U�n�!�w�ULag�Py�~���z��97$U������'xI�&�L�/�۰�\E�ZmG�u��^S����<Q.�][U�/�w�4��k�k��Av�	�d	�8X><k�4�� ���A��T̖��,����	Lf�NЌ �5M�ZW�W�}�&�����
{(8[��c��n�
��6��K�N;wh.W5Wn���!�]���P>��32&�����FA�J^��+
�D�h�����O�������J��J��1�r�b\$j{��^��뮗÷�O���(�[�qb��2�'���Ij<6D�\����_<�5q�����C�LO�ӹ�K�\LS����I��;/�q�X���'�SK@���L��B�?\���%�z�f
0UXp�&}~�ꩩ<IM�G�1C�J�%�Fq�}z����������l�8��a'��p��Y��c��M@/�-$t���o%&��QB�
��l��1��]��*��n����W}�f�	��4����xj���q�*�~�� } ��y8fI0sKy��x��ʗ3�����a�.��<8�-Z�f��ם���.Ό&�?o�:��R�a)��t�u3����sU*R�`m_N��^�Jg�x`��w�8�3��,����J�t�7_���Ng�Lll6ȹU*��rI�A�����t��.����\��H��Π��/��PA\����4\D��E���;3�,Ƴ����[�e�=��(9���@h<s����2�mi��,�����6ԣ(�IMg�}�����%��(�c�M��])��nM�um�Ɣ�d�h)�Pe��(��;��'U3�o���A�����em
�"wP!ف%`c�K�
�jB�ܨ�\���n�MM��y6M��uK?�A1T�y��{����[�C������6��K���H)Qg�3� �1�M郴�>HWդf���;]�*s�����.�'��"ֶ	� f��KLY˫2�]>�"D�/�#.B7z�ո�w��3�-O��������?�'Dny�es7_��<I'׉�6����>x���\o.D�'�q���.���{����������OV|k;�bob%��m;�k��CT
��9M�f��ϢX��7�ęW_�e�up&;$=P�q��d Ÿ"��o�M$�S�o�z���BRߴs3����K�s�ǀ�����˟�� R۰R�������d�ɣ�ϒ�]�����)��p�����/�10���yU|W:�cO��WgQ�J>Fgtq�3ƃgv�y\�;��wK"�8��T�SFoT�Zw���Z\��7��(`�j   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          �  �  �    3$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���O����O~��G��Oq���v�	&���b@�9�(�*oR"T�dYH<y�/��V�,4���L� �H�M��Uv���i�>IR���򨛀*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   .    ލp�F˸��%�R(O5f��p"O��Q   �                                  �   �	  �  �  �  ;&  /  Z9  ;D  O  �Y  �d  �o  G{  C�  ,�  H�  Р  Ҩ  �  ��  �  K�  ��  ��  �  l�  ��  ��  ?�  ��  �  � 	 v � 6 �" �( +/ m5 �; �A 9H �N �U �[ 0b &l �r �x � ^� ێ � a� ��  x�y�C˸��%�RO5d��p
�'l$���By��@0�'�F �L��|�t���pd��46B���2�ZMۓ�U�(�^�ɗjW)�B�rrf��<�X5��½�u@ �jZ�͈�P��4�^.��� ��}&.�k���@J�+֣a$pJ��;U=H�H�+E*$�]�6z��Sڟ����6V��k�`�)>dK�/	0W��;�ͮ�?g�	Kl��'�L��v��7���'n�'���L&�Z�
��֬#3��J��A���'�b�'*b^� �')B�'{��W-���$��k41�#d�'2�'��'͆$K�O��3,9�l��#�:y�*|��O_2�B�I)C�6���NB�B�Tw�(� "O�O�IK$��~I�؋0d]�]t�v�%�̠lp���0O8���� �xA��Q�{bt�H��'�R�'�����T�'�b󩂤��xФe�0)S q��B'Q\���O��d�O�l��MxӦn�#������bm��#R�?�rE�/J8Ȳ�=�
�'c�ͣ���-�l�r���~�:��G�'
�@H`�X	�Q���+'#��0���hO?eЕ��'WʬȢK�w�}A�Fy"�'�
(��+_��U[Vh�7�$����<)����z��#	;V�� �a��?Y���S�x{�x�Ņ�-%�6mJ5l|��E{R�DŉA0��H�9��1�'O	[���
vlK)#��|b�'C��H�xWH�uD�Uǀ�تh�ȓ5�	�QNL/)FHБ��N0u by��g�\���i3Ԡ���g����
�J<+�dN7Z1\ԑQ�I6�,��	��?�n͚h�$�d�p����1�`�'}���I�`B�Y����9��t���9n���On��$�;�"ec��-KvU��˙q
!�$��P��X��۽A8�ۅ�R�i�!�$D�oi|h�c��Q��[�c7�!�ĕ/F�<���<ڬ|����4/�џ�{��)�6$�����'Y�~$���G�\���Վ�O��OH�$#?I6(2��Ђ��
�Ef��ӣ%Sn�<y3��/t-�Lk��צ`����WkD�<Ң\5X8�<
5��z�X�	AV�<	�
�	7�=A��TH�����O�<���?k֒�ߺ	h� �����I��HOQ>�Ѕ�Fy$����Y�	�^�pci�<i3��?y����Sܧg12�s�#p�X��v�C9V��N�d<�F��	5���7 �G��u��Xar��߄M�h0Δ�FW~�ȓH�Y`��U�����؀h�J���\��9h3(>{E.��1`�R�'�T�}B���yR������W+eP�Y��Y�WF���#��O\�O���~>���_�et��&�>�L��A�Er�ʋ�$�:0��O��Iqi�E���e�>��#�*c���R���B�<�3�e�k7'�O����O,��U�W�����Ô�,aD*��'��˓�?Q�����b��l;�O7=��$[��D�
���!�Oj�Cqd���P�b7D˞��)��'F�	�d����o��<ѝOf�0F��)f'b�����'?2�3��?�V�'<����=E���6S�p�[�Z,��������dE)?3�Y��{��iS#F�Bp�3�A9Z<z�c�@�&��Ƀs����O���~b>9�M�.�d����$�ȅ�?���O���D�j�0���J����Ez�џ49��)�*�:�v ��;W��,^��|��!�t�(���Or�'1��#��gϑ0��1��Cm�C䉳@Ȣ�XB�MŲUI'!�e��B�I76>l��('9�����Ƕ��B�I�dG��7��?:�j� ���:��B�	-f�L�[��* �v�@�ȃ͎�1U��"|���S�~Q���A�-z�������%��ϓ�?)���?iI>���4����.�<C5�3 w�I��b�7t*!�Đ �ʬ�`�n����l�c�OȨ7�ü��`�	�8-��9�]����'�B�'�)�<i@��Ac
d˶i��n� �:��;�y2��mF��:S�5La`#�N���c����'^�7XZ��Y���� L{���+�(��à�?AL>�����#�O� �Ԫ��Wv�>���ێq���'�| ����)d�F�R��'��@R�ǖagaxB◺�?	�y��V�g:Tsť�Z�CaE�P�B�	hp ]�7��>�c�F@+P������T0�Hv4��k	�.r��ss4�/���Gx�OD�az낽?y��3�m�d=�1p�'���'�i��Y[���F�^�W�#�'v���P�S3,JVm[&�̆����'T<�4+ݞׄH���H;����'ҤL��<M��SFʎ"{�f�I���WI�O�t�1G]?~�*8�Ù�k6FEI�e�*Dx�O���'��	-w��`)d!�C\b��1,O�C��8��٠� -�E��O�?cg�B�Ʉ��HH�ږ0@�q0F�}�B䉒)���7Ȏ�Y��)zDF��o!�B�ɖ"1R��W*�;7��)�g,�\�̑��|JG��c�p�32΁�-A��Z(�Dyr!�x�2�'ɧ�O%Z�9`��,�n�qTnY��B�'�,��P(��Ĩc�M�UJ��'�f`��.C)M�p�cA�>`$�:�'c��ز�#MB�ђD�-STA��'\\e9a,T�/��0e��"'`VL�O>ɒ�I�O�X���pߠ�D�"b�B\0�	(n�8�$�O��?�'����\�M��y�p�H#�Z x�':�X�$�C�d*�0�gեX�qZ�'�ұq����L%�"��Q����'kz�ʳ��6 ]�E𲊒5M���t������G�⹂�Q$c������6#RtF{"����^u	���}�8�Z杼7/,e�m�O ��!�O���ö�Xē%s����"O�xcelM�$����G� �P�"O��P!U'|Ob]p�A�?8����"O�<��R�MP�󁏞�� �a�ə�h�D��p�Q�s��:֎��Eު�v�'��#��4�����O��q�]���H9�rRHP�"��x�ȓQ�
���ğ"Bd8�wÖ,/Ōl��w"�́�mT8�����*¤9�Pu�����;��R*Z�x� bG�h7���a����(�i.�y`"Z�3��'�#=E��� ��m�&i��V��B���/��DEF�|��O��Oq� e�&��(!:q��Mw��C�"O$aZӄJ�Y�<�9�"כXB�Q��"O�)k�kڙd'4�u�Z�t7� ��"O�z��pCВa�?tHq�u"O
m�qH�<T/�B��T4 �E1��|"#+�
\��a$���˾	�(� u�^=\%���Ih�	��L��O��gc�������L �0X"O^t��W�Zx;raE�<�4X�f"Oj� THƣAܐ��o��1��	�g"OP�+�f
'v��ɰ�#��R����' ���֘�	b $�X�*ͪ�ў0H�I8�'��s��5G�Z��1��L�����?��"j���mG�E7��(���9y<݄ȓ}�>�&�ǀb��@���Ѻ%����:�N���N	i�X SM�t�Ņȓ{��z��T q2�˓��6<h2YEb.�'p�R�0V
 2;��,i�	޳��I�Z�#<ͧ�?Y����$ P�^�B�c��L7�i���I�"W!��ɒ\bF躐A0R��{P�&�!��qq"�JO:�$��69�!�C-���P��Ę��C>Q�!�� �6h�j�!�����_�u�I�HOQ>�j����p�2��!��A�F˼<4���?����S�'��Q`�3	lB�C]\y��S�? 4�34c�������|�����"O��:v�*R���Y��){�z] "O<�3��;!���a��[5C����"OvLb"�P�t,'��D�|�j �:]���~W�a!J��ox��f��s<� ��T�۟���Oԍ�#*0�hC�	S4U66�
q"O�����@P��͸R�ݍ+���:�"O|�9���gs���#cs�e�C"Of�0um��ij�Y��_^<9�'����S�M���2�A E��}���U�ў� �C?�'&s���#��$^���VO�du��3��?a�J��� �Q�v���ĉN݆��RE!uIC$M�0D;��́#�x��ȓ��8�t�ѓ��=C�I˷D�H(��{m�j�óM���*�5f ��G�D.�'LBJy{cǍ>&3i��DE1n���IH�"#<ͧ�?�����$F�-{n<�#&��=��"3�D!X2!�R.HN�E�%mS�@���H�mP�4%!��-u��L�g�
�;���	�ˍ�1>!��T-B]�c�z��D�6� k)!�$�Be���_#a�,A�G��ɯ�HOQ>��D�	O0�C���:���hA�<9��^�?!���Sܧ^�(	��,]8;׼�jR'�)�tA�ȓ3ƞ1{�Z��61k#��6
��ȓ#:�-�t�3�6H�"/�0��ȓ(쮅��Y�����U`ՖT�JQ��r�V���A�;�X ���w\@�$��B��d�Q_�D��BR��UG��(���9w!�?b"�|b�'k��?���{N�n�!�S�|T��@�rĹ�N�D�b��J8@)��Ds�0�LD��<Qp�P>oj�!�ȓ|u�m��Ë���q��B�"A�م�I"�?Yf��^X0�*D(�șU�'�h��i����A��E��T�Q��#�D�d�O~������R��"K�c	��+�j�n0!�D�4PJ�ľߞ���	S?!�_�F1T�3�]�z� ��k�9/!���͚��]�r���*�z{џ̉����-NN}��ヾaU�(������O�i�Oj��+?	�˖<t�0t�E��M�)
x�<1w�5��-�U'x�<�W-OH�<Iw)I�]H��"y�dI"�o�A�<y%� 1>`�����iX��Ł�U�<�CƟN�AQb�B��
Ek�"�iy�6�S�Om�U)G!.��j��c"Ι0-O�Ek��OL��6��IB�lW�9yRtb���C�!��۠#�����לWK����U�I�!��ـZ x��҃��+M��@q��[�!�$��I{��L�I��Qw!�Ĉv�t�S@߂ʦ$��k��q��'5X#?�-G?Ipʓ�l ��U�-iz���	H���%���Ia�g���H9��kRDр~���p�k��@m!�$��/P��2�i�(��h;�#%:4!�dX�l���0���V��eW�E�q�!��r@�,[t�7K@�j�gI�$����OJ� 2(�%�Zu(�c�KtLe30�	-�v#~D�d�xU��anP"$�
?�?A���0?If�E6�(u���f��A%){�<�� ��?��tQUo7ez���S��R�<�� �0�,3��]9l�4��R	M�<��� �&�"M]�kgpD�V�YI�'��}�7�)Q9
��ց��!����sGş`�bL?��|
��?��O�Lk'�U2j��g]ل)��"O�����	G��=�C�>�fT��"O� �e86� <��%ŵ��"O�ʓ�r�4L���}<M"O���	ٲ8J���93f�$�Y��0��哅{Iⰳ��E��6�X�`]@~�ʓi氝����?�K>�}*D��F_��)��8V�$P& S�<���E]���X�(M�k�N��[U�<���:��ْ��\�v\-Z�m�h�<�Z�O��U�1M	&�$U!�F�y�<�'o7pV��v拡�t�J2�A�I��O����OV��,ǩi��؈�L�n��i���'��'����>����Bn�u�m�x�X��d�|�<	6F�8P�p®�ٶ�Zр]�<��K��h=8��E��!C#�b�<��a�F)V@��.h��x���]��$
�v��Ũ3̄�h�����a��aE{rjB����`@!Ņ��M�	S4 N5"f$� ���Ox�$2�Of-�6m_�B�|��1DX0K PiY�"O���N�AsrI8�[�bm"h�f"OF!����qÜ�jD���|e���B"OرмP�q!Ԗb��K2ED�=џ�(��)F��W	)Fmn��GjY��\���j�mEx�O��')�	-�8�1�#�#̀ (&���M��C䉥{R ��?0�fh�%��+��C�	/@3Tj�&�.�V|8��)��C�I93������4TA��5o��+�C�I
d���EϦV����I�G��˓Bd���|�֧˒O��Ѓ�)��~'�8E��'��|��4ȇ�
f(�Db�eh��s��ާ�y�I��$��W�	�i������$�y���a$�kB�ٮYop9j�Eݢ�y��U>�tF&��:����SH��y�^�\SD���oK)v��v`���b������c��8�cA�V�{c���Ӝ���O6�O���<�3}����l��P�g�
0k��i��ʥ�y�I�,zܮT	䆊�[
n��&!Ƨ�yb� %H~��!�עb�P�#�a��y����XBRLH%�T����u��=��?y`�'�(}�<���z$(%X�����	�5 ?�p�.�-H݀t*@	^MUjW�L����I�����(�<x��A/S	u�V�0D���!Z�!�����A(�ĭ��#0D�Ȓ�� K��8��:+���+.D�L1Ѡ�>�>|ń��Y(b�: �*�]��>75
I�<�rh�No�С��̟�XgK2��|r��?!�Oz�Ϙ5Ut�H��� D����"OlT�)�9Ę��#�5[��M�g"O����Egz���"#,:i���1"O�A1kշqL̳U �Yc8�Z�"Oʡ��$�*V�����.XA��l��\��8���S�ْ�ȷ)�.@�� P�1��_+D���?�N>�}B��Ǻ'��ȋ�>=��cSLHm�<��
�&/)�娐�M���� Bl�<Y�b�7ST��A��	�2rbPd�<y�0%R�-(��,nx�y�.AG�<�q�J{9F��l���^�I���OH����O^��ʑ6`�I�-2)�lA�'��'(B��>ٷ惠'�Y��G�og8y`Sb�<��O�Q���`��:ۅ�Nr��ȓ (�h��%U5<���K���l�p]��g=�iȖ�B�I�� ��=�4$�����?��E(i��� ���R�<�C�Ks�'2�����)T";v%cBK�TQ �a��)\��d�O�����:�$�#r�E�	6��Ň̢)�!�d|ۮ��gO��2=٤�'�!�� 2D��߀<�z�9��O=W��)W"OF�kŅ�j��AF�8�r��7����h���"�+���{�@ђJ��I(P�'���J��4�����O(�U�*�X��	#��ĄV�h���ȓV��ja.@�S�(�ˀ���,���;UP�8O�
,׺u �D������cm2��R�q�x0c�o�Vt�ȓT n���AY'<�`��#�=�|��'b#=E�dʅ���v�K�U������P���*P�T��On�Oq��!��їp����I�m�g"Opk��
�Ez.��3�S:[�����"O*�a���+?����@
�S�LIq�"O����&�n��W��5��)��"O<pA���kҢ0��� �����|"'�7���y�~p@�����E���!e.��	C��`��O��j�!�6�~����
����u"OTɪ��S�܁��Q=w����E"O|ʵl����=��,�R�zs�"O~���lR�*c�����˷)�P�j��'���䌠:xR���n+�,�Ai��ўl��G1�<��L�0�C�(�t5Y��S�AϾ)���?	
����Y�o[ |�du� L��X>,܅ȓ�M�s��5"�|a��5L����~DP��ÈN��n�Sb�T2H��*�Y�2�o��]�T��6/z�G�J4ڧo6�`�莉4�S���5Y�ވ�ɉ #<ͧ�?1������3B\@�tCC��,�	 �
>!����j��¹�� ��!L�A!�$V�^��rfݪ��:��1�"O��T�R�!w����D��Y���#"O�);֌����'�F�i<E:�V��#����3
��bC��k+X�1�&41H)��P�D2}rN��2}"��m"A�Ч�� x(��K'C�'y�'�0p�D���I���}�
�4�^mB�Jƨv��s0F¾d��4!S��?z܂ui�,P+kF̹jJ�dj/hfd #���(5�(���B&�#>	�����	V�'M)�$���4ж4�S9aZb}�'�a~�`�s�~��RnM%*�$� G�K��>��X� 	w��^�6�S!釫l`9;�ʭ<�D�<�����yr�'l��Ic�{��Z"bK��Z��'ƺ\$��5M�A�21WH��ÒQ:e�ROEdy�e�0"~�	1d��Y�W�LJ�B'JN�O����!� �) �ˊ��Ĵ�'Ԑ��?Y�O�O:�I3aҲU�Iܗ)����DC�+�B��*�
�9P��*Np�QrB�E�[��=i@���-rEA����b�AZ�-�&�ǡ�d�����?�M>���P(@�0��C�<Ap��hF��y"�K$��D�E㚐'jP��N�<�yrG��5���["�Zor �j�� �y��Pi�ĺ$h�}y�u�w��y�I�_�la`uoK�uU֤(D���?��)�_��� ĈK)D�B����mX�����?sF	���?YN>E��@I�%�t�`$S�����=�y"L��.Q��U���sU��9�y"M��F��()f@[2d( E�Q��y����#p�9R�Z�Q�������yb��
I�"��擌 ���sD����d�'����H� 24�#p`���GȠx-<��s�>�d�O���<Ofhq"�2q�)96�[(Fe�q"O*=�P�ٲ:���M�'V |�"O��$A��T̂ÆQb��ٷ"Od��_!wͰ��G4���'��ʓ:�Pg�9r�E{5,��D��?��.Kw���$�'��e��сs"<���LG��VL[��' !�V�t��U��Ί�&�D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  8  �  )  )  4  ?  �I  U  W`  �j  �q  ~z  ��  ��  P�  ��  �  &�  ��  �  ��  �  j�  ��  �  I�  ��  ��  �  ��  ��  ��  � � � � '# �) n+  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9��CZ���1.*��5���#D�������=9js����]>+-B�I�L,����ơT� *S"0G��B�I�<w<̉@���R��Xrȕ(Uv�B�	�n�t�hՈ7Cn���ӳ;�B�	x�Ψ3�E�V�B�ʑ�ޕ-bB�	�K��� L0B��h�'��O�`B�I~����b��L�5��£~�B�	�0�dq�  -Nz����� 9�0C�0>a1%
�y�N���.M7@B剖+($�w������Ο&|`!򤂰V�dS�D�
��PZv�I!��"���㰁L5=�����	�!�ӄA��a Q�&�ʀp`�0#&!�$\(�
��.B*�Z1�f��+%��O���$+$�T�J6)M3i�j�+�R!�dI(�$-��G�!P�Ȁ��ѻ*�!����UaƏ�R�2@1�O܅M�!򄕑[>J�!2��+��Dk�N��t�!���-<��A��@�uy�q�A�4�!��wI���E�9��%�k��!�,���A�k�^��Q��$#�S�OT�A���Af�Q���3�ր�
�'ؘ	Xa� �2]t��O�*�Qi
�'�\�9����,����6�D>y9
�'��a KI�}?�!��K��{%�ł	�'�P���]�fDD$P&K tsX��������>�࢓!&\0 J��]�:F��A"O���D�%5��xZGKC�& �lP�"O��c�p�bd�SK8sI���"O�a��HabV�+�'O�}]�a�a"OT��fj*6���l�EB�LK�"O�в�,1	��0�&L1y>�y "O6p�bE�jE��C'�b&��B"O�6� 6m�>�*�Ř�&vP�3"O��p�C*R�TJP@�P�LM�1"O��C1�T y�4��-��X��"O
�jQ�	�1����#��0g*���4|O� ��v��C��af����`�R�"O�Xk���f�Q���X��< �"O��a�Y`&���!O+v���"O��``J8.D����� š"OҐkqOL�y��O3yҬ�8�R�L�o�n1��C�<4½ÖdWv�yD}��M	�i��h�����a�*(�DB�I�<���G�7Zʣ��@�"=ɉ�T?Q�-Z��|�)���!F́P�=D�@�'J� rl�Zg�RUZ��4�p<����v���� O�[1c!��fn�0$��&>-���	Qx��/C�Pnp�R�BP��y��Jo�$���E< bQY�R��~���ӟ��>���۱ ��V�_�nhK�Ig�<Qm��	j�X���ߺM���R3��xy"�i?�⟢|z�!p��烑S� Ӳ�X�<���{�&��'F�f�J���J��=q`�DHJ[tOǵt����LI���hO�'y��Mh�F�X��|�`�G=q�	��|�&���5^�,�
d�I!�������s����`�)�z�PTG���
�R�d�}h<)Ħ�d<�ؘ��Ss���o�o�,G{�k�:���f�S���(��ˍ�yRH�Z;�1���O�x	�����y"A͇Y�(�1׮��t�>e��8�y¬J�;�[4��~�*��֟�yr�ϲb��#�\'o��A�b8�Py�M�^<�a'V�H�����-b�<9SI�6���ش�[(���X`��b�<�v�R�A6PP�7�$^�4͐�`�I�<�7�7'3|\� j�j�ج�ѯN�<A�*�f�42B��Z�� E�I�<��d�#L��@�É5�t��B�{�<y�l����C��T�0���"@�v�<��!ٽx������;a�$��tfJ�<ya��������6N�&��e�E�<��
|L��)�샴���
fA�<�GDޠU�>52��X2{��тvk�R�<p��.[��@U�,C�ɢ��XO�<�
�)��m{O�V�`J��Ee�<)5��$��` 4f��&���r��G`�<I�DŴ^%Z�㧖�i�d�Ä�]�<AQ��O[�qre`W<n=D%R�(�p�<a4D�x���V��A��Q��FC�<�@J<(�Rł.�𢴣�c�<�1�Ð�ZDa���:!	 �zgjYU�<����`/��%l¹!�0ZrC�X�<9�EH�K.����`D�"sz�Q��Y�<9
ԃ,�4���%��3k�(H7��S�<�⩉�4F-��T�`���+!�E�<�'�.v~�I���K�)X����ƈz�<I�e�l�����g�
��P��w�<G���f7�t13��t�rXZ�`z�<!�	02���HU�<
��!���x�<���H��a'H�F���9w.�n�<���RC�M�E�a��!�Ke�<i�/V�R@��@�ßP��A5f�W�<qg!]�On�qɅ˗ca|h�n�<)Q�H
�@q�v��͐7*g�<Q`�)iub�;.-��!�m�<q�&qP�!pC��*є��j�<��	R�|�������8�fEx �^�<�n	T}�+��n��R��W�<�2kT�fZ@�V���6eR�T\�<� �A�f�#y�E��K���p��"O�pA ��T��Eӣ*DG�ԉ*2"O�h��4X�a"+�38�li"O�2��Z�b��4���5"���"OVMK%cޭM�t��b�ͬ�����'n��'O"�'���'���'�"�'`�|A"ʓ0H`��c1j�x���6�'���'���'���' R�'���'�D<��GٛY
F%H�HVW�4�2"�'@2�'�R�'�R�'<��'���'Nx�� �����Y��ӛ$[rظU�'��'���'�'�B�'Q��'��ԫ�i��
6�Ɩ4D��Q��?���?����?1���?���?9���?a�F�k�����
��(oܕ�M_��?����?���?���?9���?I���?���l/p	xa��;I�C��.�?��?����?����?����?i���?�)�+C��!GX
+��lj���)�?i���?���?���?���?����?� F
.K�t�9Q
65�T��M�?I��?����?I��?���?���?9C�D'P5U��'�*Ϡ���E��?����?y��?��?a��?����?��*��@��}�ǧX�*g�Țí���?����?q��?����?1���?����?���B�X�ka[6�
�;�D�?q��?���?����?���?i��?�LL�p8)XF��9��@���?���?����?i���?��\8���'"i�� v��`S.��2����h����?�,O1���>�MB��_S��Ô�W$]��y�H@�<�-O�qn�x�U�����x�3�A;;���A5�C.p�ah� �����3��nZl~B?�V���m���!	֦�� ��(]�g�J�{'1O*��<�����2w�E��� _���"��#<�<��'��I㟈��6��y���l�ܭS��E9T���Q� /Mz��'��D�>�|�e����M3�'T����t=����D;�򽹟'���_ꟴc��i>U�ɘOX�|�N�%�>Б�'�:.�r�GyR�|��1��ܟt�s��3����́�UT0�T� ���џ����<I�O
��"�
9ZRr��e�t��֙���	#:"9�,4��:,���[1G�K�ĥKE#��hcٱ��~y�^���)��<!��G ���×F��~L<��6�yt�"�>�/OD\���w��iK��6Ѷ̨��	�o�L*�'��'��L� ��V��ϧ���-ɾ4�zq9�E3��q��F�u�t�'�x�����'���'O��'��H��@SԈ��)�*V��tr4\��ѪOv��?�J~��I��a�,aCh�HS���j���؟$�?�|z@gK��,:�c��&NR�h�/�*T�fIP�έ���K�L)���:�L�OD��ƅ�R�V56�Z���W'�N���	��d�O<���H#��D�u�_k~�a)��O n�[�$��	ߟ\��ǟ�9H[�L2�X�ւ$F��������v-oZT~"J��p�'�䧲�/�NݙrT�sX�1���&/`q���?�Uh9$#����fZ��X�Q���?Q��?�Y����p$����+֚	��9��U3]ZH��4�IK�Iß��i>��D�]ǦI�u'.*Tsя?{rVI�IB23�4�R��'�x�&��'��O�H��ɱx�ne㕌8C��ٺ"�	:��D�Oh��O�˧voD9�GP�VY��""5�t��'���?i���S�T���"����۷Nc���B�Z�5���*b��6$�j�<�'�@��X�I�Q�]�叒a2Q�1�	@��B�	��M�V��# h=Q�@$*��9���_�<���?� �i��O�<�'��NƆ���RU�l$�L���*���' �K�i��	�ip��HUҟ��u������5�F��L:Z��1���$,|O ��%2Hn��s�j���9U%�l}2�'p��'��l�mzީ)�A�aJ�K*�
#s�q�������Iq�)�S�N�"Em��<�Q��{��� v��Ds*��+�<���h�&��u�	uyb]�@H��̇`9>� �*Ka��Ͱ��<O\��'�'��d��4�	�td ��c\1��O��'M��'f�'�� 	R��@�u���Q�f���.?	b�V�u#�݊�4&��O�D���?1fHZ�hӼ<���6k�zL�4bʆ�?���?����?����O ۧ�Ԑ]�D%�U�C��a�O$��'R�'֖7�2�i��%�فz��D�1 ۀ��S��d��I��,����`s����p�b�?��A'
����&��Yo�th���z�IKy�O��'��'�2
x����2��	a�T� A�-������O����O����YQ�n����Ӱ^�,���!P�1�'b�'�ɧ�O��������\�& kQ�	�9�|��Ћ��v!�V�����,B�n��d7�D�<1��B�S��t����grȬ"����?i��?����?�'��P}R�'��!Z2�1&�6=��ڥ�ESC�'��7-6�	���D�O���O
L�&C��Z�`���$W�d3�����L10}v7�3?����.R��|:�{�? ���jӽu��y�"(�$��15O4���O���OR��O��?a���D��saٶL2�$�ǟ������K�O0ʓY#���|2�U�h޲�Bp�P/]-P�����+��'��T�e�ߦ�'X}�F�	X�h��I�;h�����Z#h����j��'��i��'IR�'g��)sf͓7��)�gE�(>���'L�Z�<�O����O��d�|*����"��T�S�l(��I��f�{�I��?�O[�Qsl��Z"4p��I��2����0'$���CC@�i>����'|$$���F:6��� Qi:D�� �ٟD�I�l���b>��'G�6-N7 O������H��T��Jĺx,��O��D ֦��?!RU���I�O���:&
*O�R�ʕ��9-2��	쟴9�o���'�����Sbr-O��h�nE�v��
؀|�����'��I�L��ǟ����l�IB�EѮ��� uF��M�(B���0Z`t등?���?�J~���l���w�晊�lF�5� ƹp;���'O�O1���ؖ)i�J�	�v1䔳�f�@����B��xC�:O�������?T*&�$�<����?�©E�&��!fb['\��������?���?y���d�L}��'���'@��sfa��5t��%�����DT^}b�'l��|b��p��H��_�|���q������ݿJ�F�k� |Ә�&?�P��O��$ѣR�ʐb��4Ա��#,����O��$�O��D2ڧ�?��	�"�,l�"��7<<J���B��?��[���	ş���4���yG�0P%�T�T(J�O�paBGE<�yR�'R�'*��KV�i��i�	��?)uf�>T���0�Jy���a�� N.�'{��˟����(���x�I�n/�M��Ǉ�72��k�aF�Q��'������O^�?���9 ���$g�M�@�����O��b>��mB�q+!3���6f�>$ e����`y��Ud$��
\��'b�	5)�\I�qI�)LS�0��>w�A�	؟D�	�8�i>M�'����?i���o�*��g�Ƙzf�}�eL���?�ĺi��O���'���'���<Q��\��2�(���D�'Rp8ǸiK�I�I�Dqb�Oq����X�*-�3-��Z8@�Z��"���O2��On��O��$=��%OL��2����Z,�v��8��Q���(�����Ĳ<"�i:�'����@�;o`���#J�J�Asך|��'��O�}ôi#�ɪk��(zP� +S��(���Lm�x��LV'��L�gy�O(��'�"`ŒQ�l�R/�y���r�Y"r�'������O��D�O\ʧR�A�.ǽ>��v�/��'if��?����S�T�̂;��U8�"E�����Q�*e�ʔ��*� o_������~�|��0q0�2E�¡;&1����-��'S��'����Q�jش��C(��
�`#c�S9�<��?��?��čL}��'=��n?�2�y�o�<&�����'�B�� ���������?g���<I�	�Lt����sN� y0@�<�,O���O����Ob��OTʧ]�����t��ܸ�B�K���Q�[���I��t��l�s�@k����q�	�%
r�1��l� ̣֠�0�?Y�����ʹy��?O���H*`�x)K�G��8Ͷu4O���W�2�?��L2�Ķ<����?��E�=�\������imnQ�SGF�?��?Y����D�y}�X��	9�APm�PMpT( 	$��?R� ��ߟ\$��#��G�T��Fr�8���-?� ��z��ɔ���'r �����?y`�ݺi<�铰��H'h���K�'�?q���?i��?���)�Ol���cC�=�ijw��'?2���F�O^t�'5�	<�MS��w�2h��KQ=S�N���דz(ٚ'���':��).�期���!��JE�M�F7n0P�B�2z��+�F2p-xX$�����D�'_b�'���')Z�$�>���X��w ��1Q� �O���?����I�����$f���������?1����Ş= �i�Ȝ��  ���^
q`���Ab����'�*�Q�.���a�|�^�$�\�-�ܐ������Jj���?���?Y��|�-O8��'
�βa�
M�t&�E�\`�"��q���,*�O����O��d�)4F������T�<ݨ���'n:r@��o�(�g���cj-ʧ���,�d��A3�G���fI�<����?����?���?���$��4q��YB�I�a!�49R*� a���'����>ͧ�?15�i�'��t#G�/cj���.U60�����|��'��O."�i��	�6��]�iD	)41�Ǩ�=���� q���8�d�<!���?)��?1�%ˣU�c�E�Y5j(9�+���?�����Ēc}��'P��'��3�^��IM*���9,H�"���3Y�I��0��Z�)����-6���	ceöS�����T:������M;�O�	�/�~��|�m�'zj�0ipm�b���]�e�r�'�r�'����Q��[޴:� �H"o�:Zv��K�%k<A�����E�?��[���I�D��u��Չ'q�ҥ�C���I��D)㦉�'�0�@��I�?���� �!9C��$G���r�]|xFM�S?O�ʓ�?���?	��?I�����g�h7� � ��@���}�'��'�����'�6=�rl�N�jcL���-b��y�#�Od��%��)�bm�6-`�H�Qh�3;��ǉ�~� q;%�j��1�@=p�BPw�I}y�O���	`B���F_�Nb������'�"�'B�'C�ɀ����O��D�O~��E���IBoY&^�Z����7��:��D�O��$9��Z�a�`u *�&� �t, ��^R5+�! Fx&?�BE�'F\�I,V�����f�k��qaK[�s�X���ߟT��ԟ�	i�O��]�OP�=i�C�Ke��ɶ�]"�>���?�"�ia�O��B5K�+�о4�}��k��'��'��'Qc���4��AׁB����Xrct��s�*LHA�� n;.�O&��?����?����?����Ε�]|!5.�pe��/Fy↲>����?����䧌?���7��@!vH�*�o>6�	�p�I[�)�Ӝ)WI�l�<AR|���+#&Ybdޝ$�~�WF$�"D�O���O>�*O��fg|=Z�ӗO�M�B��OF�$�O����O�i�<9�U�@�Ƀ)q�H(���4��r5f�9�5���M3����>����� O�>�H�ρ/7��sKU�ĉ�Ԫuӄ�58�`��3J~��;�E"s,������V�z=:��o���	��L�I�$��՟$���e &́@S�Qk�|� �]��?1��?q7[�P�'.�7�<�D!Z����$%RZ4��I�'&��O��D�O�I�7#�7�-?�B���^�;�ሥ^U��*k���i���'�D�'���'���'_�pCA֫<��D�G�ƹNk꼹��'=�[�h)�O~��O0��|��ÚL�r�ZsjԷGp�M"�[@~�B�>!���?�L>�O.�i0�ʂA�Nm���GJ�T��"�#@����T���4�� 	��-��O���ƒ�VH�͐fmT-P-B(Ј�O^���O���O1��˓{t���P>&�VH��-A^P$ze���<A*O�Mm�j��D^��ӟTQq�ɊZ�	QЯ�9q�hKmy��Z'xқV�����O��� Ey��[q��y��
X�5	|�p����y�X� �	�� �	�h��ğ4�O��\:�d�F�k7%^)�zARc��S}"�'��'���y��s���+�"4���>#9Rq�͖;B�n�$�Ot�O1��� 
p�R�I�F��p� .,�$�gf�G$�I7Xp�*��'lv�%�������'c�\��
�x&JH�C,_��h�S�'��'��X�<èO���O����;$ց	6#Z9LEȥ��3[G⟤	�O��$�O��OX}��F�K��Ġ�C"y�z�����l�A$G�'c:)J��&��>'f"�F��G-A��c�� @fٲ�&��<�	�p����dG��w���̶t�	�u�W6�tK �'��ꓑ?���/��4�L�DꐐqheɃ	�@4���q0O���<�vJ���M��O���E#����DjBxQ����R [�^dۓ�r��OTʓ�?	��?	���?���?�ֱ�ĥ�eMҬ��)��R����*O���'���'����'Ǡ�H��+F@j��I9L\>0X��>1���?�J>�|�BJ/��ɘ[�w����/��I�����C~��_�K�����>2�'���6���BC��2{I(Tv�ѝȤ������ǟ�i>͗'.�듇?��_�N����tk�1�$��
3�?�F�i��O,%�'�"S�hR��J&E�IL<��,���#~�6�n�O~�`��&��0��$�O��cA�D�ac���&�h����	�y��'f��'&�'��	O?b��ڱeg=ة�vd�:u��d�O~��F}�W���ش��!��Ts�g� C��P�P|[�8J>Q��?ͧ8�(��4��$H=��tcBޒ$Mpb��Q�Ufґ����?�$'�d�<ͧ�?����?��i��/�\9S��W,|(J5��H�)�?����ĝo}"�'�2�'��S��<kn�m5&�C���0��$��	ߟ���q�)���?@�B��4
�A�6}�����A�.�Mc�O�)҇�~��|��L]�e���9�T�P��"�'���'_��t]�hs޴x ��HCnR�>��%eLt�l�Γ�?I��x_����T}�'�P�`��oc���-	�2�	u�'�B��Ƒ�֝�ow������	�u(9o��r��h2�a\�$>�ry��'i��'���'�RS>���I8.Z�aD���?����Q�����O����OP�?�������V;�\#�l�,���"�M�?����S�'*���۴�y��̃�:l��IB��U�ժC�yb�æu��������O���RT�V��S��R�  `��K6�j���O����O��g��	П��	��P���f�|�Y�ܪb��l��}�����៤�Ij�	7q)����IW $�
�UON�r�AH^��]'���L~�E�O����<bޡ��'̡D�2$�ナo������?Y��?����h���$�Dh���T���i$mZ @����$�S}�'rbiӈ���I��9�#��Z���"�(ߨ�p�	ß8����e!�1�'�Ȅ��ʀv� ��T�O�W*�q �T�P���0	,���<�'�?A���?q���?1R�֚΄͠�fF[��y���DV}�'w�'�Ou�����ȝ��N���XqW�W�5-���?I����S�'Z�\qD��s����b,ř	GRq�hN��M{�O$9ĭ_ �~r�|�_���pdӊ'����N��<"Θ1��ܟ8��̟H��՟�S^y2"�>)�w�XQ2Ќɫ/��<`��^�A��0K��%�����As}��'�'䄰'M2F�>y`���T� e�t,�f2���\�t���9"Q>q�%K�B�)G� ��y���N�H���	����	���������G�'���.�&��U8r��o������?9�>��i>��	�M�K>��#ʸ�.M���P��S���䓐?Q��|��II��Mc�O�n�8��95�V�T�Z|Җ� 9p\�l��A�Oz� O>�(O��d�O����Od�r�L�F�BF�ߏvd�yX�&�OV���<��R������	x��)��4�4<�Q���:�$|�A ���d|}Z�M����S�D�M��5{% �v�r��ʎu�@��Th$X)�����#���=��V<� ��޾��lHQB��R���O��$�O���ɫ<1T�i�� nܛ/�"�����^�*�'��ɖ�MS����>��{\�!S�F��A�f�߬NK�����?y2���M{�O����"�>��O?m;����{Ep�)mN3y��`a��'�"�'�R�'e��'��ӑ-��B��3%�%BrL��at�Y�O����O���)���OX8oz���k��\E7O:�ĀJtL�P��D�)擙	n�l��<��"N!�y��A��z{�1	���<�"�'S��$����$�O��d�
9G���D�k�~u`U�'K���$�O��d�O|���	����ޟ���BH9t�\es�J�,D���0CjJ��:k�Iџ���n�I�z�$Ec�m�%{����#kK3�K���S��E(��|�,�O<����?�p����I�R$�3)�<|.%��?!���?��h���Q����#�I��0Q��e�Շ�O�p�'_剻�M{��w
�y�N�d�>@)�ݤk_���'K�'��� !W@�6���Bw�d+������h�X$̞� MƘ��'�����$�'~�'t��'�V��A+� >�
y�5FO(B�d8p[���O����Op��6��@�^�2A	�#fv'�	�.�ic�Ox�$�OL�O1�F����_5}�d����(\�*}:�J!*�j7m�~yB�Ӊ@A�������$.|���d��kuD�!ܖ���OL���OF�4�˓��Iޟ��$	�(	D\1B�
-� �@�!���4��'���?���?A1㏘)�d�Ǐ;C�u+EA<2��ش���5$�x���O��O.�DkU� ���f�ѱF��,�yB�'��'���'��I�8J�����C�:�k<R�r�d�Oh���]}�OI�}�X�O�XI���`��!�h��/�d��)�d�O��4�>���q�b�"V�|�D��.�ޱh*�S����g$S�L�v������4����O��9["D�c�-W�Hp��B����O˓S,��֟$���|�O�8�x�[i����"_ dtZ�O���'�b��?9ѧ��$VD;��>� w�}<h��E��D����$�Rџ��|b@FQ��C3�y:�R@bQ))>����O8�$�O0��)�<�!�i[�}�%MT�'����j��Z�ZA�'���'�|6�3�ɪ��d�O�LH����\I1ϛ�a�Y�˶<���V��M��O>И`HJ�2& �<��$C�?����;t,�z�l�<�+O����O"���O�D�O�˧; ���-�Y|�CQ-�$Њ�2S����ʟ��	_�'3ݛ�w��`QO���16j)Ex�m�E�'p�O1���{�ja� �
=rh|"���\�� ��:!���'��tٵ�'���&�p�'���'w0�����4,�� �K�4u�-���'�"�'��U����OT�$�O���
XnYc���h�&�P��O�,������O.���O"�OJ�i�_9.�R��jA&P��۔���Z�&T�rt�#�B[��ss��ɟ�w΅�*�5��@��وXg*��'���'�S����d,�=�z5��Ѓ����p\ɟ|X�Oʓ7��V�4��e	Qn�� 0PT*������<OV��O����(�F7-;?�����;�j�iE9[*`K�"�ci�p
�-�1U��M>)O���O����O��O�3�#�<q�����*�����<�6T�(��ߟ��	{�ߟ�� .
�?kؕ
	���@������O���,��i(TF�Sѥ.�`�;�Q�4�1GMn���DA<��4���p%�T�'�r���] ?���ڋVq�my��'p2�'+�����V�h �Op���"cwЙ�G��o��P�j�9#�d���?)gZ� ��ԟp�I @|h�H7�ͯ��aZ¥� `�V%��E�'���`PA��?�is��4�w�Vq	��9�2u�N5���!�'�B�'���'��'��~8) �7zv��p#`�h��qk�<A�w,�)*5�i��'#�8�I3QZ�ig�C�.�
M��yb�'N�	%7V<lZt~"�
>߀ �C`�K$`ÎԔ[��-`RiA.�?�d+�ġ<����?����?	S+�$���0լ�<? ��3�@�?q����N}��'�"�''哱T<�A�ɖg�н �[����$��I����I[�)
�f[-ٖ��0�.Y�\��3)�1l�rC�#C�����Vǟ8#4�|Bd�&B����፻?	А� Y4&_��'��'3��Q��Y�4):�:1�X�+)8ȁ'oԳC1����?���^��F�d�|}"�'/�d�ˇ�^�萢�7.l�)��'�r��O�&����A�׭9q��i�f�X�|�Q��[,��d1O�˓�?����?Q���?�����ا#W@�����7?	03�C]�u���'��'�Ҝ���'�p6=�2��`%�H��d�P�F��Q(�OB�D!��IM^�6-w��(q"׮>>P���,�4A�(p��� U�z�I�Q�	Jy�O~bJ�/�Tq�$hJ�T��A1F��B�'��'d�I9��D�O��D�O����3Ŝ����K �&�,��3���O\��5�dT����"L�4
�M���ù*��	< 9����s_�c>���'U�i�	B�}��C56A�����X[���	͟���Ɵ$��Y�OHRL
=ͰQ�
"J�1eʗ\���>�(O}m�Ӽ붂;J٘A�ʍ�]-���'��<���?��]�xP)�4���Wn�H���'�Fh�%�� d�踶�*Hj��dO$���<�'�?��?���?��eˍh�X%I���F��놻��Cz}�S�h�IK��/"X��sК� �i��8��R���	韸$�b>��W��r���R���j�K�@ԅJղ�nZq~�.�	Q(Y������$C>N�	�p�[�F1���2g��?K
��O����O>�4��˓?��Iǟ����+0�z1ZF͉ou��c�g��k�4��'����?Y)O��[�f^>���hխU�~Ota�Y��耹i���.,�!Q��Oy��&?��*^I��5"�7<�f����2����	۟,��������O�(!ٗl^�qJpI�$�*
L����'��'%���|b���6�|B
�9c�(�C
W�L�bl(�C��v��'�����Ԭ���V���B���k�.T�gٯ_G%	R#I�=}�)���O|�O��|���?��?>�=
A�T�5���QtBZaĊ���?!*O
E�'=����O�*�ÎO ̆��͛!����O9�'�2�'�ɧ���k�uA�9RX�]0Q�O�@�Lm0$-ǒN^ܙsE���S
%�B��|���Bt�D�2����"����	����ǟ��)�SNy��g�llC7n�-���ѡ�ék�V�p�1O|�$�O��n�h����՟�F)�)G�P�+��uT��BL�ȟ������l�P~B�Q-T�H����$�z9��3$J3O��|��h����<I���?���?y���?�/������� =j�u��Gr.�ծA}�'2��'��O1�}��.�:a��% �?E��V���o�B���OēO1�Ę3�D{���	�jHu��65���Ù�v`�	�;�8[��O.�O���?���G��$DLݟ8���a�@��jB9���?i���?)O.��'�"�'���	�F<�;R�:|@�9�A(]��O:�'�R�$�)�Z��w柧V4R*�"Q�g���?O�hhRF통Z�6�&?IB�'�6��ɉr7�ybM�y�L|��I�@�����������O�O$"F�IN������X0@쒢sirG�>����?!q�i�O�NT�Gd<�A�J	����E*\����Odʓ|$VȻ�4��d�*d]H���'Edd�d��*;�~��Fυ%\r�*�i/��<����?���?����?�f.�	s��-��)�5J&"(Q�Q���DUk}��'���'��O�rh��,����\�H������>�l듿?1���Ş1�a3&D�\�t��㏪'*\�� �Q6cV��/O���s���?	Q7�D�<�boܡE]���GY�e��5�Uπ��?����?���?�'��D�{}��'k��*�h�^ݻ�B��8����'�h6M7�������O�ʓ��y�,ǣ^�lU"k�2_��5�Ԏ̥�M��O~-��,B����>�	��`a�"-�%SoĐ /g�D��2O`���O����O���O��?�y�Ï(lJxc�/�O}6%�!'Eݟ��I��x�O�i�O0�lZA�	R�PP�A$�0 �6�����*%����̟�ӧn�I~҄�((��Ę�lHHp�n�9D�t��@�IFy�Of�'H".^,_�xs���@�H�M�'��'��:��D�O���O�˧3Y4��1+T�s!rPW*�3q})�'�X��?9���S�ďU7��j�i��:�f�A{��!Q�
F.N�F���O�iW�?��2�_!�e�:/^�z�+h�2��O��$�O~��i�<	ķiD�u���6x:dAB��h�<Q��'��	��M���B�>!��Th��j�}hr����.#K�|J*O`���b��*�z�������r(O�
�/�k���C�'�5��h�9On��?���?���?q���מG�~%�A�
ܸh5�_	e-�'����&?��	.�M�;0ذ-4�ǸoF��3�%S�����?�N>�|��%�M˞�� �����-�f��0葵�&tr�3O�p��?iQH"���<ͧ�?eB��qD���@��"Y���פ�
�?A��?�����$]}��'�R�'Q��PB�O8@t�c�&�d�IA���o}B�'��O\�Y��W���&�5�f�jb��4�EO@�FH�Q+�D�Y�S�GM�D�˟P��"+\��,�=C��V�M����O����O���1ڧ�?�w�J�>�0�\2ܭ�G�����������<饴iL�O��0f��h`�X�rq�e��W�*O��OH���O(
Dm���gP���#Ꟍ-��C�$p��@GS�/`�q���䓬�4����O&���O.�䌘&������}_N�#t��	 N��sg�Iiy��'��OG⡘�,�Z�bN��.P�1��'��!X���?����ŞV�0r�~�ء�钗x�&%�gƃ"g�@�'�Jb�Ɵ�П|"_�@hდ4I����M�Q���r�'NΟD��՟�����SyRh�>���'q��r�����T��owF<q�"���D }��'���'���Q&�B*��k�/ǖu]<5�Ξ`��摟p��lF���'��@�8�2�&�"Fd��)R.	����Ǖ;=sj\�����?�zU2���BL$Isr$�(Z!�Z#*U �� ��Ő1+�<�2K�	A�L-�CE�$��a��0��~�$̢<#N�0aT*�(�#�7 ���H�aW/n�.�@�HŠ�::�����Q"+6EB񈖏^B�C�L� @ƕ#�%N3%b�C�Й�ԁ%m_�j��D�b�4~�X-�q�GB��HW+K91Z��vח�Dt��oZ	Y�h,R��>j|(X��۞:q`�%��6-���'�B�'0Bʥ>Q.Ob�䰟 `C�$%���I���	WonE�"��c�%�`�I۟X�I�w`iP����>�xy����9�ߴ�?�����d�O6���O��Ok,Q�&�$��6ђZ�bU�ӡ�'O��Ec���	^y��'s2�'y�'�l��$�Q5��P�[�Z�@�nZEy��'��'5�'��'N6�A�U7�P�C�T�DArț ��12��'q��'���4ן(}���S�M^� �4i�0:!��×�i���'B�|��'�l��D\9'*������YU��`'N��Y��	������*L|�-�l�d�
yP�	 1K+qސ�9���)1n�qm�ݟ(&����ݟ|�u�TS���I�ƙfZ�t���&g�5mɟ�ISy"�'��ꧤ?���?yR�C,z���T��$X�كs�S�NK�'H�'����'��'��	R"X>Tg� K="ȓg�Y)B�[�����P�I���ɟp��5�@�:o���B�L��pX�Ƀ��M[��?��@�����O��c@ F+���cl�4,o�I�ش�?���?����?Y���D�O��DBz��A�5Ō��Lh(lw֜��?E�D�'!X���Ã�Z���b���*Dl���M{�:�d�O���O,d�'��I۟��{�TX!��N6�Q7��(��qnK�I�lb��L|Z���?���V�[��+r  � �G=eR����i�B�'�����OV�Ok��"U ��C�Ѻ3<�:wnۧ8i�I- $��$�h�	�����y�� %x<yc���$~1l*�C�7ě&h�>�/O��$4���O��d�8s �t��X�T|pA#�4U�<��� �$�O����O쒟1̧<��`��N'ڈD�Db�a�˓�?�I>���?�A�B��~��ܴx�`�$6U#�&R��d�Or�$�O��&>�騟���Q�5%lm�q�Z�Y�@pp��1�8�m�͟�'�t��͟�z�o�Iܓ'�^�z�� 7��  R�S7G�2mm��4��Vy��'GV�>�d�Ok� _G�%�C/[�pqsW��.S�'���ן@��T�s���
F�zP��9�Jb��{Ml6m�<��f��&Ŧ~"��?!ᛟ��G�Z{ry�3��):l�*C�f����?���76�OP��M����8,e�4�oM'Zܬ���G�˦���)�M���?��?qҔx��*�)��9jX�i֝^��L`$�i���'Z|ʟ�I1H��5��N���*I�lȑߴ�?�*O��d�<�O��*h����Pv����[��h��cP��O���~����~r���h�����(8$�#�C��M���?Y+OFU�Oi�O�5����m��V���B&?�d�'�4 r�3�	����'��d
7rczġu��"\@�#�I�V^���	ޟ��?���~Ri�v�m��$�(w~���R���M� �\��?Y)OD˓���
1A�xiFw?HJw�ك�M���?���'!�	<MU�6��?�����֨�T��\.�')RR���'�ş�A �U�q9�cƨ�9��m��B���Mc�"�'��	�FfO��{0O	~
�T	��W/7��=9��i?"\���'������9��$�@���<�`E;�k.��O���<��Fx��u�өC�
(i�ޏ%��Ad�V��M3-Oz���mڮ�����ON��p�_�v6d<�[�|C��GXh�f�'7��'��	-�9OR��i@4΀�N�6Z�T	~r��7$�>A���?!��?����?�3�#T�v�x`���\�k��*���D��b>���T����ЂY-g�J<�a%�O�x�A�4�?����?A��Ik�����'���#� n�J3(��\���O>��!h��iD��'!�� ��9OD���O��� �F�9@������ *��5m蟰�	&���|j��?�-OD��!C΁C$����ݰe θ9Nͦ��'��T�,�����ISyZc"R��do�������3��\i�"e�.a�'��	ӟ�'�b�'MR͎6;�Ց�c��_DLk�k �z�\0�'1���<��ß��'�"Ih>��
�$9d4  5|w�HD�z�D˓�?!+OF��O��$F�#��$�o���0�M����ȵ�G6C���n��X�	��8�I_y�O-^ꧺ?�1"8�q� ��B��W�XSAbxnZߟ��'��'|���y�\��y���#DFm�&�ܳ�Ƙx�ʘ�M+��?q.O���Q�d�''��'Ǝp�D�^�"���Y�eV&�LL�5j�>a��?!��HJ �����/G�,i@���$QeH�VjK��M,OT����	� ���@�O�N���t�B�?8��m�L?���'s�� �y��~���OY�-�t�O�|���+)NL���4�?ib�i}B�'&"�'�J���d�q��)���M�bH>���J�Qt�lڋv=P�ǟ�'��z�䖲l���1F��#��hX�A3G��l�����Пh�������<����~b ;�f=�ᮏ6x��d�чE����<	wER~�O�b�'��s��� �̷.�ܥ Ɛ4V.<7M�OV�DF{}bR�(�IHyr�5F��*D{�{q�]�Z�^u�VBH��ď�/��D�<����?�����S�/���xE����H�2�]&7��V}�Y���	Sy��'b��'��4�c�U�0�bc  ��|��ю�yBU���џ��J�8���@5玔B<�1f�!J՞q� �i�����'�B�'���]����A���J^k"Q�i{�����	֟�K|��V?5���P"�|)�N]3��)�"�7f�ă�4�?q+O���O~�Z�L��|�Q`ȣpV}B0�̪T|�2tB�^�f�'8bS��I����O���O�MP��	�s�~ڥMg�U�R����Ov���OD�3Ol�'�?��O��P��oΞ�c�G�^��;ܴ���O��n������Ɵ��ɀ����2��ƾ#�d0��O?1�P��i�b�'����'R�]��}�qcƕz^��GSЋ���6M�O��lZ�`��ퟨ�ɡ���<Yp�3`�D���E�`��ʆ���Q,�)��yR�'���p���?هk�h���&�R��Wh�y�6�'�2�'��L�>�-O��D�� ���B��A	�Y�2��+�>*Op�ǚ���ޟ���埸�s�+E�R`cF�I�h�e�Mk��?�6S�\�'�b\�X�i��!�FŢ5˺a��)�
����>Q�.�W~"�'U��'��P�֝�4�����B�bj�0�w.	?"�~6m�S}"V���	Zy2�'�b�'@ E�Q���%+���׍�}
@� �j6�y��'��'���'/�i>��OA��CqD[�PJ&���*�R�z-Rٴ��$�ON��?!��?��o}��D�7�0��t�v�@�J��Mc���?���?�)O��C�D�5�g��f����PB�t�h%��� �M{�����O���O���5O�'S2���D�VH���D+!�ڴ�?9����$�O,��O��'��Ά�gl��y��9b��]��ɫa\�ꓘ?)���?�$(d~rZ�|��>+xؒ>M��Ty�D4��mZOy��'J�7��Ol�$�OV�Dt}Zw��	�ԉ��F�l\�e�ٴ�?������'r�Ix�'VB���N�KL� ��ܝ=�x�0���Ц-����H�	����O�˓L/
1;�O�
T�\��3�ȼ¸l3�ie���'vrS������)���$Q�Q@ŋ6.�$��i���'��'����O*�I*3h5	�/��Xɜ����Ƿ��c��D�+�	����I�L�UJ2/~��N��'�( � ���MK��?q�T�X�'��_�\�i��i��!w�,U�ǅ�^�2I�c�>9@c�p~��'@Zf��'��i݅����=��4*T��;*�B�By�D��'.�	ӟĔ'/��'M�6]�:�	\ QBq���6���(�O���O
�$�O6��|�B<��H���Y��V��:M��R���ɦ��'=�\���	ϟ��	Tx ��g�H���@���N�X7,W�#�P�O��OP���G��5����O����/JTx��kR8j�������e�INy2�'��'��q�'p��O��I�̌=,�խ�&�!��iO��'���'8�y�����O���O2<S3������T�ѩp�v�)b�ͦ9�IHy��'	����O �X��s��=��]�9�씪��<i�$*��i��	��PS�4�?���?a�i�i݉��脵d��
�Ε�0��]B�i����O
�0�2Oj9��y��I�8r8�\�pͅf�z(�����=֛��'��7��O��D�Oz���u}"W�p�a���X�q1��?gt��&���M�Wύ�<����"������U�J�en]���Q5����Á$�M��?)��?Q��x�'���O��9�+U�.T�1��úvx`��iD�')�H�!6��Ob�D�O���Չ�>�(+P �@����S)����Iڟ$Z�}��'�ɧ5�oTSa���#�ܨ/VP�AF�C����Y�1OH���Oj�$-�dg��j��÷*&b(ъ��M�d�$�O�Oj��O0�� py�u@5F�@��!�O�}���XG@�<Y,O��$�OF�D1�i��|"A���+�D�K2��$+��Q/�E}r�'N|b�'O�i� �ybA&@��]�2H�L؉�d�'�,��?���?Qg��Dj!�)ؿ��ũ�"j:���W1O��$l�Ο�'�"�':ҍԎ���>!6�_�$�3�Z�^kP���ɦ��I̟X�'�rA)�)�O4��]EZ���S�И�rש5_��$���I�Ċ ��x&�D��ESL��D��54�`���^�Z	o�iyR�'�f6m�p���'U&?9�%*4J�cwƕJ�-�ĠT���	�d���W㟘&���}���׿Tl��1t��?�0���G���I�M���?����?�7�x��'��¢�	����1Ǉ(*�ac�s�.�0a�O�O>�I%'Ƕ, ���6�+�ȟ�2}��J�4�?����?��#��'���'W�dӒ7D��ANĹ?+���̇
k�֖|B��yʟ��D�OP��_�J��O|�@xrb�5N>-m��|�	���'>��|Zc �=��
�&bJ�$�?j�t責O�0@fN�O�˓�?���?�O?�Ha��&P�Z���� �hav��#	r����>������?���u�N�h��W�O���ٓ̀v�v`���?�,O��D�O��$3�I��|r  ]1F�� n9xm����B���'�������Y�㟰�j�R@�(q'G�?q0h�k�����O���ON$>��K|RPʖ7)Y�T�E֯M�^ �თ�6�'�';"�'̼@��d�F�,�c�U�O���ySɂ�ab���'O�Y���I��'�?���#��&jn	����# p��i�Y쓽��O(�֝�C�!��0oLm�)*�@��񄘓U�XIk�E҃j���rюcЉ9���|d\�H+	 �0pPp���|��X��8+�r�Wn�9I���)�W�Ow�8�a��z��s$i��HM$��5�.�"PK�l�3]��h��P���9�!d�A���� 6�����)$*Y��)ʚ"xP! �فP�Da1!��]���9a�M�E�ւ=��S����oϬ	r�|���̇7��Dإ-6��|��eʊg;�����J�G�J\blȢJ�ܘv�ɍ#�z<�P�_� 6�YxfϷH0��V�q8�g+jx��4�?���?A/O&���O���!	�"�J�qӃ��]�4���O����, �˰mⶇ�w8��k椃( ��!�p:�yڡɃ#'L��7@a�|��
߆k����	*�`����Q*T�D��Ĥ�BlP�I$F���Ot�=�)O��jg��K�lE����.i�X��R"Oj�������Q����<�+MI@���)�<i2��-Z~���H�v۠��a�ƍ�>e�4JT�c��'C�^���I�̧g��)kv�%�J���A�=~�P��$ �$��0���ir�@����i�Ӈ@�ZR�3������9`"��gD�S�* �ϓ�������i'��IB.Ş1.���l�q�'�џ�1����w��qԢC;��)��3D�h� '>("t"�� ��P��q���Op�G��3P���	H�$��n?���T��}�X�z&۲�y��'�r�'q�*�-��~@@t�Fo�F}*���!�9o��5 ��xcƤړ�I>
=�)�"-� �4�)��t�5����7H�v��M;%ɚ��(O�%� �'��IS0X�(C׏�py���3 "f�$/�OV���G�+�b��!gީ="yk��'�O�h�u��.��4Z0EG�_��E ?O^%@��NC}r�'g�O*��'0�EB8�o_	/��p��p ���ƫ1�:��$DV}*��c>�����s�X4[��H�z�#��M�N�VeBD���6���X�"~��!�t5�BGA&b�X�xWM�"M{ܼ)�O�����	G~J~BI>��5�Z0�T Q�І�a�<i�d��j�4�QGϐ�\;t����Q[�'kH#=�O�<�TCY2�^��8"2�@B�O8�D��O�p�nZ4�I՟(�'��'?h�b9�`�-��X� ���'��	tÞ�[����1Ov$�F@��[˚#w��9��D��O`�E���S(LL!�8�4��-^-|��C`P�a�pd��,������O���%ړ��� L\�9�)/t ĺ�aG�!�,f�L��)˼T��Q����@�~=Ezʟ�ʓ[��i�5�a�U�"�蠳m�)�>�qW�'���'��IƟ|���D��d��9D^��ܴP�`d�F�Kd�ܡ��]� H`|���NR^Ȩ�O�(�v=J�+ r�1 �%�{-���r��+$�H���ý��'=t9�3&X�,�l�`Aj 4�b�w����<�����2�ӧ(L�{��Р[@�X�l x�C�I5xt޵�C&ٌ/T�J���=� ��঍B�4�򄈦,��n���It��B�VFm� !E*Hz��9�ş-�y�'��'LreC��'1O�&a�=�$Γ�WcЕ�'C�(Ӏ�<�����O�9�A
z�l[��UjP	��䕱"��dLȐ��hi��a��)��"O� ��;��^�o|(t�I�����'�F�O�W�ؤq��)�$�K<G�@Pz�'"���֏��$�Ot�����O*�d�4tE��P�!R������GO�Q���$�ʧ���?!��$0F�8�.ȴ�bI!r�1r�� C�ɧ����;1݊�J@ע_�6�iYhԼ��'d��'����OH�+e�W%;~�d`���>F0�H�9OX��+�O�E�ՀW��H8�h�b��j��ɯ�HO�S��Ѫ/�ҝ�u�p�
��I��$!�M�9�M����?�������O��0$�>p��ᚠm���h%��J���Q9���3׋*lO�T�p�_�)�M�#$�w�%Z'�O��1�� ���D�,��,Д�A�h��uH�M}f�L�Mi���O��ԟ�ϟ �'p�����Q���Oü;� �'�Bt����*5N
��HH�]�Ṉ"�;�S�T��O�VT�P�E�u��ܫ� ��KC!�$��]��y���Q�nq` oUo�!�Ĕ Y�2�a 	�7:E�wn^�&�!�A��Urۓ���]3�p��F]�<�G�^=��0G/8(�"`\�<�f�Xò	���7!�pc�f@�<Yt�`�5�QD�7Gȭ;0TP�<���.J��cg,^���D�G�<�M��)���F�=
r�tk�B�l�<�2�Kz��L��j�~���'M�}�<�Q��(0����B�?	�����u�<�L�$=�&�St`��wJt�p`�Zy�<I�e��Kt�I$␗[=X�(uCM�<1C`X�B�0i��
�"�P0G�_�<��`��C\�d�C��v����v�<���37�����O�'��5Q��J�<Y�c��ܡ&�SUvLQ�I�H�<AFK��2L�7'��?�DU;��j�<)�#
	:cL��(��`��B�<� �<BZp��,��]@�J}�<9�.&	��ib� RI�H����{�<��(F
��(���@{"E@a�y�<!��X�8��q�C"�^iz#ŀv�<�̝ 8��(�buc�Dz��L�<�0O"p�v���K�"[�0%j��[E�<��'_�EB�xAꎪ�칱�g�E�<9ʋj�pv*ՠ��=y�k|�<a6�@g�4X׫ GJmz��x�<a�;d�2tآ�ٙI�$Y�&��M�<9t�����k��Z�m�8�9"���<�2nFC8Hȃ����N�� �e�<���`�썚�c�t���ۦ�Of�<1�g_�G�04"�"W�{G�6�"T�H����"yBy��iM�.�Aj'&D�@� ˈQrHM���8a�Q��"D�t2k �qr�ݛ$�zBi� �?D�����bD���AK1W���"D����"S)@��Jqa�}�@d҆m?D�����Eh�ܝ� M�8@*`�>D���f�v��9�O3f�0��@�&D�P�G��)5��S�K߶5�Pe�D*D��ir�c���1�5Zph���'D���⦊2h�M�B�\#JmV�Ke+D�Ȫq�ɗ.�v`ñMY�3�2x�2�)D���D��*ЀK`�U��$�`��'D�`� �>M ���"*U���$D��s ���əd`I�V5�dB8D�d��͗�L��M$J��LU:@A9D�4Y�㛩ed2�!&,��O~rd�$}�L�Ȓ]�S�'0'`ax�jT�hN y �$��r+݅ȓZTD�g��X	D04h�l��=Y��2v��� ��H�EK�n��e ��xK�aj�
Oj���#����GH/���񫜖oȞ�q
�'�©�"c4"�J	�B.J>��Ǔaؘ�j�`*扐o"22�4Iޞ0a1�� c�xC�	�3���a���8϶��f�$�nO�Mۗ(�|�S�'R�D勱��3(�5���;-�,��C�,2#e�m]R�	�m�TU�ȓ,��Ҁ�V|p��%U$j�Q���B=	!���7�!J���Y��I�� �fkХ{5P�� zn�U#�'�A`���@��@PD��c�T���'S(�0�ذ �bt� �ڿ?�ݓ�']��зD֗	'��s�n�+��<J�'{��A�:MG<��H�F
tQ�'���� ��qL�i����'I�����'���!�ǀ-;���
ŢڔK-ؕ��'��H���[���"EJ>���'�p '�x^�u"" ]
Ut����'7E��(N�O��UZ�-ƺI`�l��'�0� 6��5	�Ļ�����)h�'�\�	�<���20�$� ��'�Z�*B�E�BikT��6z�~<�M>i����j�6��@��$m�A2�� �!��D���C��Qclx3P�H6��O�;��'���b"x�� aaCU�4 �'RR ����|H�+�hF�{�cu�xh!�d%6�}� �)צq`����DyZw��Sf��
�@!�����!4WHx��D7�nm`��2�y�]c�)C��W�Y �:Ui�99�D3�c�Do~��AH?E��'���:�R!�(d�জ.�9K�'Q��C���e�Z�C��A,vW��I�'��AR�� -�`s���0<�ʏ!��Vmzi�4�Uk��h�C��}$Jp[��@�wSt��fX�*���ɒ��dy3M'�Hæ�L�/6<���,�υ͞&�O�X�XT�%��Iy��|���&a1�`�b)��6���CL*Upu��"O��ذ�E���10B���H[B�]�McJ��u/�>C�T0�h��e��n��C'�:�@!�60$��xi��􍓶Xp4qB�n�7?jp��+�_8h��O`eF}���J<�?�a���S�
�T��S"f����^QX�b%���o&D�p�퓝b����Ζ?c�H��v�� ��+סP9hl�1�$�O��q��9  �P�hҽE��dc��|�`M�ea��=M~�@/�?%>�[�'Ԉ\H�z�L�|�^-��O-D�ܣ��·O!dU��AA�E�$�QBF�Zk�}�JF��X�O���H򧌜�<��]Q�
�4Y���RH<ahY��jG@�	��)�d�S<d�D�6� e����V<�A�闗(��Z��M�S�N�J3�M=L}^�Q�2<ON�H7�]�^�S���Oة�Fٚ^�"	˴��[�d3a�.Đ��a&�Px�14�A�9`x����&Ii�Aꖧ$���	��@蒯�0�e���/���|r�2/1.�E�Г:��ѫ���D�<	�B�' ��[R��� 3SV�0��]sJ��e5Z1˥�P}��d���y�U���Z�
j��@�����yr$Вn��Z���  $)	Q��-��$�l,(%AY�2�n�9`Y(䑞��\0J@���K�0M����+\O��q	\�<;b��V��/0U�$O1v��/B�a��q�Q-  ra3�>�O�`���S	CV}���'�,�Z ��K-�r�-N>�$[�-G\��ԟ�u����vY6A�&S�9�d� �A�?�pC���(�z�HADզ.s��;�9q��X���G�T�Tl�6��C\`�C���,O�����W�׿[ᄥ�G��/F�~�Sa�<q��ѩ+�j-j�EH
,���� 7��lZ��˓h���5�yZm�&�]�L���#O�J��o��Qޤ	�i-�O\��"eX��U�&�!#�!)%D�.=�X�X�Dͫ*9�6���$�̓�Խ��+,����9ǧ�0�@4 gP�Fx�*�4�w�_�q�`�['�*�M�矤Ia��u��	�K@<eN�y�\�T&L�S��'���g*�O�μ��f�* Qp� �O�:&rA���܋��� *�M�g���� R�ZƤZQ�9�!d�>�j0�"Od�����:4be�G�o���HVMF�y�0BT�SC�i>�	�j}!�T��y��@�O?��EҲYo܄@���x��P��:�r��D�k�>����t8@����0iq�4�@'��g�$I�<�l:몴�nN�=�L�O���f>?yF)�
4��T+��̾�~rțKb�%�"��>2�TM[�O��� �Ll���'(3,O��;Q� Z3���$��Qeհ]�0D)OH���W��f͂�A����.O��؁)b�U��g �8��%�j]'V�xu�<������%)��:lg�T�$��m���*��"n�����]��]�BA)?Q��ܹ��GO�pqd=�̸q�g���f��Fj^t� L�eY�̺1��sqO��̹s�o�r�hѬN�x��H8��4��'���� J�E�G_9� X7`��
��O�h���9>�U�&ݶ#h@P���x�!\�-�Ё�'8��c0�z݅��
j��}�RmU0q�����U����Q�'��c(�(^4�ԣ�@8�D1�w� ����5;�;�I������V��
 �!8J�ط�[;��a:�n=�韔8 �-\�k�IA�Q/�����	�/a"]�4����袓� $~<�4��E�M]2��^B��׀K�Wy6t� Mםc�R���?;�V�J�F4��O����h ��O��i�IS�@R��JD'�D����=%'��#�&��;�N��N��B�����(�⟄���5 �t�ɱ62h��5CJ(!�.qY�]7��>�e�#^���{#D��H9n\B���$��8�1��w�$��Ǔ_�.#^3����L�[��=SaXo����YF�h%�"zN�g�
*.^����$U�hY�qF k�Pp�F��֏@�?�L�ZpBº(��ib��C��0<�b�ǢS��D��G;]��l�C�����Y�S���ߖ�z�N:VZ1�'̤<��$�7���ւɦ@��+��ĝ�P�3���B��0J�;(̙q��3x^ *�@)c̨5�ʍ;CP�=y�¦x�xH�	D�f�8)���7p,m�Ç�+a}�P�w.�R�݃�8A#q�F�%
�����o����$ϲHB̨PA�J��� � �*��խx�� y��B��nU)�R%!t�*�E��<5������#e.���IlzL�E�G<(q���8s6݀��*�I%jX��`�\n1OX���`�Xf�,���R�PФ�'�fQ���ঙɄ+�c�BԱRH������>���jT#>9�d�.8Q���I�xmt��N��T����x��WN�Y`��S�E\a�܍�iݵ��o7�U�R fFـ1�@ !���K^��&���'ސ�Pa%�a�gy�@	7�Ay��Wk-BT! �O��~��C=������9zZ�-A�E�"m@�uaB�H�`X�1#uT.6���vf9�S�\i ���&	�x�Ж`��pm#?I�O0g�4�?�2���\� ��D�5o����4��YP���H�tX��A��>�[��r�,�2N��PѠ��S�L��'��p����f�S�OB$���V�>�;����.�����4�0��$K§>'�z�#<O�]�7�E-G4��e�P�FN�1 �x�ց��>�O�H��s��%�VH��'Z��D�R2��v�l����-1�Ь�4�I�H��Z��]��52bdϜ��d_%B�Ι���#��4b�A�pџ�8c"SD�O*\��M�.�Ll�]���U��'�� �i�)]k�d0�ޒ�0��'+.
橐'+\؋DHQ~e(P��'�R�26�`X䫞+pOdu��'��BS��"`�)ಅЄnr���'����Fԓp��U!�C �i��<Z�'o���S0{l�E�ma ���'��<���!W��� ��a*�I��'j	���?&oT����X�l5r�'�`�a"JW����@曹Km����'F��:�C�#��y�$#�0<5���'~�æMȅ\'.��3lB&7o��y� ֟/8]x�H�=R�����9�y�N���ܻ���#kΊ`MX��y�++>z=��&��g�X�R�Z��y�L�?[L�H�D��<d�tl��N�yr̀��4��$ˡ��X�����y2mJ�"�X@QM $>��j�lʎ�y2%G�_P�˅��f�P��Ҏ� �y�("{�l:6n�)?�	IN��y�$���2�N$~@����y
� ܌��G9I1C4�U�,��"O��QV�յm@��(C3��	c"O*qQ�2Ȋ�� hN�s|j9�"OA�D�0���H���҆"O��x�۩l^H0¡5k��P�"OX��FB�&|����߂m��t�5"O@��Iτs#�9S��
&	��'k	����	�`�8��U'aT�	�'�F�(�K�VRw+�#�Tu��'�� �*���Ћ�ˀ6!tx��'�*y�K�8M��	f@S��\��'/Z�#�cÁ}̸�p�R���̉�'��ܐ��D&w�"5C��`�=a�'�� w��$Zm2�G�3Q0		�'5��c���3
����A��l��'B��h��N���B,M�P��A
�'� ���
c��1���X���	�')�	�#H�*YA��Y�{����	�'�n�"2��L��R7c�(�0��'�T��%�j.��Uf�t���K�'�xkċ��"�v�"V.��Z
�'������Ў�zgh��6�����'mN�k���?V6����L��"��`��'�����#Ƣc�^lY����H�R�'���h借�Lʜ����J #�p��'���j�j�'�T�(�(U�x3p��'�dI��8|{f��>�H|��'Rn��gOܚz� ��R�5�`��'l��X��ڌމ��W�5��yB�'���2WZ���J�Z�.,[�'�8qÊ� ��� z�I!�`�<�q��R��<�%�*~ ���\�<�a��3.� ��㊋C�yǹu�<)�#���rC�w攑!M�<��J<����eOq��Ã�Iq�<iG�B=]xQ:*Z�p���Մm�<�e��3�,�Cu@ϱ9�<\sBM�d�<U��+a��K�D�za��G1D��37 �9S�0̑�5�D�J�.D�T*��ˣ?:)b�Kʣdp�I��>D���`Y*l���r����\�*>D�88���%AVxP� �ߔ:����&�=D�|�Eʄ4r����dߐ�3�'!D�4@��ND@���cH���^���?D�@@�H )�
�E�/�HxȦ,<D�8I�	H[�$�`��J�$�kUb:D��S�fXC��4�p��4��i5�"D�<"��K�b�1�BI�:o��X�/ D��!��Mx�B3'ۆRr��3$�!D�l��X4>�
Uɓ��*Zz��em:D��O�0;aD�F�D|��Q-.D��bP)�%�L�ZF"�Kƪ�h�(D���B�U�\����_��FS�:D����~�Z�P���ug3D��(a���r���%h�
��QN3D�֠� ���Z��g4+u /D���!S�< �{�)ׯ �V(�. D�4b�nG�K ���@G�L�f)"D����ϙl��B5D�2I�����!D��kDK�C2�t�"�0K���a��?D����@�� ,��.d;��Ԡ>D�p{7%��u���"5G�I�d�=D��QSe�b��Ф�sWz���:D�t�� �w�V�pƄ��v�:��"D�� �����Q��0�"�>5��t�"O���C���L�s �D�*@�$�O&�=E��+~*�#�23a��x��W��y�\�&���P���%���h���(OT����H5��#&iE� ����� ��!�d�%G��e:2'@<lrp���3u!�d&#riRoڿʜ��GB$0\!��>���2`��O�����*i[!�D@�_Ø�kY" .����d0!�DkZ^����0�@�1�E�<#!���q��]�͋9`��p�$M>u	!��8m�����
���#�@��!�D�	��Q�d

�2�f0��a�!��[�,�|��UĊ���)�t@(�!�dͅ_�Z|[�K�a��Y; �Х
�!��
�(������
-����&>�!�d��'�z�(�]e�T� O���!��'��S���.",���aV�/2�C�I@i�s�J�4ev��T�ֳ�6m-� )Ȁ�z"	qa�"^,v�a�4D��3F��h���I
9�V�K�J=D�D(����EHZ\�4}��d'D�r��tA
��7W'�,izJ&D����M�C�q$,�f��9��%D��*��S
��\ �	ʩ
h�����$D��@���U1xM�rg[#6h�ѱ�!��oZ\bԀF��B�t0°j�d�B�ɞ9��})BQ�vn�
��X4?u
B䉚x��_>�� X�m��C�	�;�>�ڦ`G91�I��!Ԫ"<�C�ɜQ��pi� �$s�� J4 R�Xs4B�I82A���[,`W��[E`��gH�C��N�f�K���#�|�x�02�'�F����P�X��އ����'��5�F�]������Yr^���	�'(h����!5ָ�'�F%8�� �b�fA3�k��D�N`;�'��D�ua�3je��h�CB�0�	�'�t0'�r��� ���MHp��	�'��M��F1A���B@C>.P���'hx �O]&1��ͱ������r�'n !��D��@�
肥�'&R�Q�']�|Ch��G1~�z�#�'���Zc�-�ɚ���!o��)��'^< �ïH���ЁiT�w�P܈�'�P�c�d�50oBd���s"	�
�'-*����H0EF(m�� �FQ

�'���eO�8s��`�6o�6��	�'=� ��,E.)(ٰ4�Nn��X	�'��ͩ#��&B2p��m��z�͙�'�\�!�ķ'�:�r"B�zn2Tش�Px� �)h�*=Zv	&�6��'����y�G���%Zc7$֠�k����y��F3:�� C���j�(i����y�5Dn�qTy�r�[fm\�y��J�,0�)R��d�r��`<�y2��d<(�,]�%�<�Ł��y�n�5"� �b�N��v�c�o��yK4"� �N��daq���<�yRD��V��<�rc�(BK �Bc�5�y��g�r�Q��٘O������.�y"�ym�P�E��{����sH�yboE�xqysA()��|sI
��y�j>vF������.Q:"J�;�y
� J1�vl�F������1%^�l�"OR����A�U��L�1R"O��;��z;~�)��Ė+�T)��"OF�ST�ʈqd�Q�.P�hҞ]�e"O�X��	>1�,]��J=mĸ`"P"O�e�DNQ&3JL�*Y�I�jT��"O��WA	!@|���G�1l�r��e"O�1j I^)]��R(��1��q�g"O���o��,�ƹ��ĉ)����"Op}�Gn�*(Dx��`ŭCo��W"O��fFǾp;���&��pQH��"O�����N�t�����J�	8>���"Oia*1n��M(���J��h¤"O�$�bɉ�V�x��jW8ḧzC"O�� ��:1,��Y�C�zXr8�&"O��P�#5Y�� 0Ç�fh�2"O����-W2:89�� jL"Ը "O8�PVk��r�I���A"l-Ј+"Op��@	�<V�갓�F	�v�y"O��@�Cm$��vc�+��I#�"O�P���I���8c@۾`��'nqO�ţ /U�X²U�DH��{+�a�"OJ$BL�}0���eI�"�=��O���	�'X�.�r���>:>(�E�C9C�!��=,�8�0nZ�;Y��AC�'	�!���B#4$f�y��N�iNL�"Ob�
p`=�(��`�y���@"O2i�cl��M�D���(��vRhA�Id�OGB%!D �8����_�~��91�',8\`��G�w��2�m�2le��C�'��x*��8F- |"#�׾d�B���'�8�� �F
:T.T�uEǣ+"�!P��(O תR����QKɯf,�#�"O�U.����5�4�rMC���:�!�<"T��A5�H�ȅ�Q�|�!�dN�5�R� A፯�$�HA[�k\!���x�@Q���M	\f� Ӽj@!�d�	kW<���a����A@\�D,!�D�&���qh�9�	/��X!���+xl�˕�F�
:ҎҺ!�!��Gx��2f �~1J�-G?4�!��8%�\�⤂+o0�Q���P�n�!�S�}D�	Gb9�HM�K��!�Q6UL��;�hA��`�IF�Eh!�$�1��Y��,��ՅΉ�&x�6"Ox9*P
 z�3�䎌V}�Q��"Oа��̜�q�@�QiN�	���"O�
g�U�k�0�mf��ehU"O,T��vT�eJ�*�d�r(a�"O^��D�\�b��=����X��M��"Opi@��I�4$�ے�&twtSV"O���R*N�:4������@q.�!�"O"}z�)S�|�2	�ȸp� (�"O�q���'+Ȳ@
N�:�Y�"O��b#/5p���҈Ѿ60F��S"O!S��B�� �e(1|,@�"O8X�C�A�޵%(�I���"O8�㔮�!D�B-�&G�\�̡�"O|�c�U3C76<����[�4Qb"O��1��OGCh�1�&�&��(�w"O8��um�#m�$���D?X�TKV"Ovh�qc׎~ �U"��L��� "Oљ@�ʪk �2��5�JD��"O`|IpCJ dj����!C���1"O� �� �L;Z��1e�!�☁�"Oz��3�2y�1�Bǟ����"O8����A�����H�/l����"OX�� Jא1�N4���gdtU�6"Ovx��R�@��d�&�)S���"OJ ���9�Ҵ��f�21V��`"O�m
0!��u�� ��D(�	�"O��9���*V�Lb���%&�yu"O�p������R�n��Hr�"OPm1��U{5�A�pM�7c,�RU"O��C �
�!�,U���!e(���"OL��kV����4L�ZF"O��X�\1Ć��M�hs�I��"O�ő�&��?�e���$�3"Ob� ��V
�jŢ�ΰk�!Pr"O�Y���Ӆ^��3H�2P�L R"O���
PF�R�h������"O��c �J2�A�!�9-��+r"O�!�MLm:	�ao˭q����"O����J�q6~�SC.��\%�`0"O�M1W�*}y� rM�	����"On����y��q���߄2 ���"O�|��R5�n�QM�
Iy�Y�"Of]�b��m�&՘PM��q�ʑx�"O��2��;����N�u�5�E"OhPy�hް �mD))����"OT("d(��b�1ɛ�Z�2QS�"O� �r��<�,��)�t�U:�"OjMCVʆ+D����1��SE@�[R"O�Hs��˶*��X�AN6-;vqi�"OJ�"��9J�+��$�d��"O,�s��ē>�$�@��>䉈�"O$�@AO�c"��Zbi�6Nd�g"O6\�6锿_�ѵ�1 (8b�"OP�BG�1�4�Q��߭]�����"O��aH�	�8-��2��ȱ"O��ʴl�'a��� %��
��7"O�9�o�6`Ű����чwMp$�g"O���4i� 3�:�Ic!��xKpH
�"O�0:��F�tDi���Z6�1`"O�c#ه.s��˅M�f'L�;B"OH����|�aB��,km��)W"O<��%n�LM�M߆$^R0�#"O*	x@�٨�Ĩ��L�>y\N� �"O�P�-[�2����]�gW�!kd"O�%M��|�px{��A� j�ՊB"O�E�g��%(�<�"eF>	,nl[�"O��"�N�T��H��i�b��1��"OU��G�1a2����ڬH���P'"O���7+�(I�Xe��t\�9b"Ot,��צ�y�"X�!ǔI1�"Ot��ë��8���;�g��Y�HEI�"O�0R5ˁQ���Cv��7g��	�"O��82
]�mD�` �N����9�"O `�&��P2��RT�D�E`��w"O�\fe_����k�O��/�Z}�"O�\�C�ޘc/�$��+S�V���#b"O���.�p�O%�hIx�"O�H!�LS)TIE�WB
@��q�@"Oҵ�&t�إ�@N~U��"O�����ݻV�����HZ29�\Q*g"O� H�M�00�ǇH� �N�A�"OR$#M��$�1�B;x*�-	�"O*����4^uP���
 K�"O� YH��VqQ@�`�l����"O*�CŧQ�<i�Ub�2�(8y�"OB́�oTTߔ���G��jX
�"Olz�Ē����2g�+�� 1"O>@ �GO/�$s�5B�=�v"O4�w�[�7�ػ�b�E�HH��"O�Æ(�nT��;�a�QJ���"O�����\3 �3�J��34�I "O`H{��L�E��43 T9 �"O�ē!��D�l`2%L��u#�"O�9kG�~&4*�-��(�"S"O�P�C�]_�E��"8�N���"O0�X�	�~����L6O �-�&"Oz��쟞 ^`A*�4[����"O�<�b��p�.ءI� *W0qc�"O��rE(��=d$鲓���Bl�4(E"OX�C�/�B��(1�A�����"O\̻4��% ����� � yzL��"O�,��nV�Xc�[�w�n!�`"OP�ae
��b���P���u�ba�"OFx@���9p�UzR�U�JM.M�"O��)�C����! H4^�h<��"O�ܱ$j�X�^�b!)ޔ�Q8�"OРP)��/V�� ��_���"O��ʣ$��TMp$C�\��4"O�dZ��N0'��h�i�9b��"O��Хd�<w�L�#�T�X��;�"O� SG�ػ(6h�#�@Q|��"O,��A	άVH�$+3��0FN�-��"Ot�K���A�4���I<\5*t�"O��SFI	N�P�ǩմ$'
3"OxQ��	�#5Ь{���� �K�"Ob%DOњT��E�0p��l��"O�ԄJ�!������5�n)�"O� ��	>�� �V�=	(�%��"O��A�UBz��'$�Ql9�r"OB���6>-��ɗ�ڨj7"O
!�TĤL�J�A��!�d|�"O"��i�=���>��p��"O�11KA0V��a�OZ�7�xe��"O�T���)�D�"�M=��,�"Or�᳃H~�P֍��k�
�J�"O�-�Re�Z�T<kЌ�>��]7"OJDk�;4`j	xd,� Kt��"O"�;�7CY�|�P��<v���"O>��e��o{�HX�Z�T/x��D"O�`�"M�"����T@[+H \�3�"O�$�1)˗y�s��շF㨠yA"O]�ahL�Ѩ���.ćU�Ь%"O*y+7�_�	����P8��) "O��Є0�N��Eh�U�����"O��c����3��J�f�-V*�00"O,̢����4��,y�σ9ɀ�"O�A���F�2�ع��EԔI߀��t"O�h�K�]���N��Hbj�"O
hȱME�F9�%��`P��@�"O�`ՒM��]Y����V�ܕ��"O���Ehĭ:�����A'2�ȡ�"O�e5�	�`��<�v �n�h�bW"Ot<5"��q^h�	��H���ɓ"Ozy���=��E�2(H�.���f"O�	���h���ض&P�U	V�"O�$�2OZ8	���F
<L��"OX��&a��Th�����U�5� ��"O� �d!��-��a��ܑ�T��r"O�ʠ��oK֑��Ę��8D"O� ��Hک<|���L ���6"O��+2@'+*!;5K�`�6IK�"Old2 �w"P�s���>llɂw"Ob��͗7����7i�`/H��R"O�X��7|�JyB�匞l8��g"O|1��LF�d���z�Z�M�d� "O��`7h�=DkZ!�O�O���s�"O��Y6���|���"%�z��lʥ"O�U ���Y�~���D�##�hQs1"Oa"���Q��\��
^EA�"O$M��l!����� �ru��"O���'���]fN�����l��["O������ ��$�'�ު;Y��YU"Oh`�@�X$v��DАFO�OE�S""O�Q�qb�8o��z�EY�U(��0"OZ��A�Z�,*E�BF	��"O�L���U�*����㐍`�NM�"ObX��c��~,p��~bL�"O����.5i�,I���AV��A�"O����H��.� )�A�A PLYq"O����N����G�rk��!r�|��'�ԩ�r�Y	��I
#��#&�N1��'�z0� Q�{8"" �7����'H,��mS�rBvAz�'��,��-B�!�4O�63��	�'��t��m��=}F�@�R>�]�'D�XC֡E�)���g�ݗB+0��'P�z��O�:i��f�ˊ4@(���'� <
��͚F`R9{W�\�%��U������5Ax��c�=�Z���Cv�!�W�~������L�4���
�!�Ē�i<�l!�J�"I��pG�B�!��[�>�I�6�7>~a�V'S0�џ�D�ԁ�9��		��ȡx���)6�y�\+*�<�&������W��+�y�2�*P�a�OwU8'����yr��d�B�	cb	�Đ[v/�y�٠K�P F@��U[�mӥY5�yr�����[DgA�N�&��R �$�yr%=r �|SA��;N	,���T�yŧ�V����oڙئY7��xb��v�t)cN�s����u�F
ZV!�d������P/�z	.�*M�'�ў�>��Ɗ�1"$� �֟4o�e�%�#D���&+Ԗ,0�b�-.h�Bq�"D�(�"CїE�(�C R."g�T1��!D��Vfܭ_��lp*�"n
��$�>D��3 �:#�|�SJK�|���s�9ړ�0|����+�� �&`�p�7�o�<���C$`4�d�!mz�:���� m�<YrL,,�1��r^f ���h�<�T���l��Lu��Xc�� O�<1FiO�^<a��\6��%bI�<Q���("���1�A	K��#cI�<I��H�{�2 It�V
	S�aB��@�'=�	Z�Oe���T�)B��e�P�o��T9��x�iG��D����-�Ȍ:W̞���x��X�=��������y��r�
��p�!��X1!�f|XaaY-1��s�(Ɲ1�!�DR�R��*�M�G�����:!�߶@�t�y@�8`*"쒐늑c:!��|�MB�� ��YB��Ζ(+�'���5�)� j�S��Of��8�	ч1����6"Oz@çm�9+P�qF��HE�2�'���	}Q�h�2���\�sn�<B�8C�I�+Z���[X���"e�	�C�I9L����d}7PH��`)<+C��?F��!�f�-��l��V�B��,(ҰI�����,4i�0I��B�ɤh}<p�ԧٟ�9
���}��C�	�~������J��g�Q-r�v�HG{J?�K�CW2�,�e�+T!� �C˷<��_`��#��]�~�L$#6�JI��ȓy��sT���tE��_1|�p�ȓ)@��)���P�v��ti�*�ZɆȓ/l%9�KT(,`����h<p��	���d̓m��dY����Ro6|�sA��bN�����	���O<�b��>��ȓ$��Bd�%p����6�Μ
RE�ȓWў0���G]=��icb5-ά��j�n(���30�$�)�b���W��0�D�e�Zq�C!Q/��݇�NR���&j¥~�B	�e�Tf
���7�����	Q��8YE$XiG u��i�p;���U��IX�I�	bI�݇ȓ��Y	U��3~�|��Gib\�?I�Z��0se��7H�b��׿,O:��ȓ��B��́LF�Z�D:;�>���#� �IMV�gR��2󋙲%�rq�ȓ�b�
#�\�b쑐h�?~0E�?y�Y�dŘe�5�^�9Qi&h����	�<��NF{(���BX^A�%�Cl�<Y�1K�J�,ߗC����TaL��<��~��j��~�?��q�q�Ņ#�b���*�yRL[S��]!�$e��C�3�y��c��B�.�8n怼�ă�y��/>*�L �A`� A�b�F��y�πj�: �3U,RX� R���%�?Q/Op�O?Q��H_U2H��e
.6Hiw�h�<9���M�����N�x�c�b�<�ABP )G,��	�%�b�P�jCu�<Q��? t�Ҳ@�9j�X���Bs�<�����(��&��=JwAům�<�cI%o��[U� ��0���ZOy��)ʧh�T��Gꅤ^�0����)!@xɄ�Ix�'��y�S��): ��+4�Y�,ٸ(O��=E���!q��xJT'�6 
}�G"D�h���z��4.K>'iH�hB�5D�H`GLT`IҗJ	�*&HAs�5D�̓ᧉ�g;�9�a(����)��2D�d25A��Y����Do�8�9ʰ<y���ӯu}���
j�F(�1�֔F�.C�	#F�Z�saL�b"��+��N�C�ɷF�I"$
T8���.�'��B�f-�qR���&_�8��v�.�xB䉉GƦ)�%GDx,�1���TB䉍s6�2�(��ww,m�e�E�R=B�I�İ f���0|�vl�r�@C�ɢS�D,��#�>hy�:C�B�I&+�����@� Y����旐n\⟈�I[��~�4L�b�c�����ѭ'2Ѕ�*���QaJ��Lq��2�*]����ȓ.'\̨c�?NΌ�6Û1�|�ȓy��� w�V����$�01y��ȓf�~t��Yn���&��R,���Ɠ>Ќ��v��U����ȮU{����� ��I1�ͅ7s4%�'d��D5HW�	|�'���	��a�)�nI�Z�#ۈx�'*a|b��%�J �Mߢ���B�_��y"N�����;�&�� ̛�ْ�yr��*��T����.0�� CD"�y�&U:�ȱ�&�*-� �a��_��yB��5�����B��#0�&�y"�.��JcB��"�Ǖ#�y""�9*��$�0�f|s�a@?�y��N�>�Y3�ވ!:v�z�ꖂ�yr��������: W�U;�k���y%�/��-�ņ�-e��;4��y$yf��pk�I���hE���O�㟢|�N�j�l����Z�l�XiIE�<���U��(�[�.b�@F�B�<!�M 2�޽A�!��(��k�z�<A�Ŋ8{"d���=a$�(ÊJu�<��i2�C�ܻb��b��U�<� �/% pr�Ahzd�"P|�'?}00N).����t	(~�x���=D�LPp͋�d"b�SL��|�p|���-D��s�A׼3��Pf��VD���*��0|�Q��6��U�T�K����TkQN�<�'��(a�u҅ ��v��`'�Eb�<Iu&��2��@�!Y!�$���M�`�<YA�P�zX(%��)`�}е��Y����<���3NTUs���5A��Saf�S�<Q��,C�>1 l�Yl���e�<���O�+%H���? ����'Dߟ$��	n~bC\�4��ID'�r=J<Y�*�>�y"W<Q���k�>!+�)К�yB��'($�Kp�Xu�"��i�4�y���N\�̴֣r�Z!��QG�<9��W]8�ݲDB�[ZH���Wy��'h
�R��5B���ۢ��5&�M�
�'�^y�R��>!��I�I�K���
�'�f����MH�cG�Ld�X��'���:�IE�Er��ã!�Q4p��'���z��ɺ/�֡����)�~1A�'��0n�)wS��pԎWf�x��'k�8�H	
*h�Sϙ�Vy��[N>y�����O.���eۀW�M"g��w?� �'�tU�-ԃh��2S7��@���8�� �S�5�T����V��y�h��^1��O"�=�}ZTB�+[�xH��_�mb�&]D�<����-*�8�/<_6�Q��[�<Qw��N �E9��2F�k�k
ş�G{��I��k(C�Ḅw����h�v$ʓ�?	���߶������ʼ��㘿2�!򄋝����؝��iQ���{B�$G�����УNV{r�F��3�!�DZ�i��`�H�"U�A�NO��!��Y�2�x�`���sP Q��:�!��?#��`���N��̋�b�!�W0Ly���B׶��RK�O�!�ЋQ�d�y��%�\=C�/�
+�!���c��`�l��2���;�U�W�!�Ęr6�Ia�"������f�]&u�!�$�6�|���`7��D�g���'�����.^A�Ǉ[�C�ֹ��'�Q���" _��`���B h��'&f����ޟp�%Y!&�/���M>9���i�4_,,(u��A7v�xen��O�!򤖓�z�I��$8T��B�!�� ��Ha��%[B�9�XG2��"O���Fۏo��T����7;��if"O�Bt��	�`8��_OV�
R"O^x�sk�?H���Q 2B��p"OV-�Ca�G�>�!�i�#AC�8��Z����}�S�Of�}�W���LU�D�a\�K0�I��'����̐�U��l'ѥG�����'?�Tq����3o�A�D�c���'��ĸkY��Qs���4@��'�`u!�D�oFx�҂��FR�m��'�Ti�S��2��1(�#�?�)�'f���'R4A6���������'���B�T�85����u^н*�'��X��D0)�*��$l��' �J5�=+�hXq$��q5����'��k'�Г��ѵ 't����'qp��w`�j�#�g!e�|�+�'��y#�!�z* ��ۈ[T�("�'Jt ��9
��'�+��QB�"Or�#��zg����L7�\�5"Oґ��Ƥi+�q˱�<7v���"O����
a���D�O�Ҍ.�yrM�ր�:�GU���\�%^2�y�*�TQ�����c6t�F��?�y�a�{\(���8Zl��p�Ί��D%�O.iK�`�(�"=x�JxP1�S����I�,e�vH�V+y�D��-LB䉊y4�ѥHڿ,������� �4�=	
çK�l��n� 9\ɹc�I<]4�ĕ'ua~������r���*$@�mK��y�ļ0�-�s��Bi^v��,s�'�N\1ā�)x �`�
ͅf40yK���'!<��`�aXp��LUp��:
�'��ch�	hV%pl;��x	�'%Jh�q�+)��8b��X�Z�8	�'V�:���&3�U	ECzA�j��y�-Ү^�
��`F\*9��%��y�'։H��*PX4,��4{�)D��y�k�#Y(�u����U�4��� ��y"�(!Ib-��P4=����'É��y��V��f{K�5S�]��bC�yҦ��Q
�牾A%N]���D-�O�@�"Զx�Eᅎ�6;�T�A�"O`*f��y�@B4��v�lS�"O(�06EZ(W�~Q��_�@j��A�"O�)� �5�@�
6C۠S�P��"O�XV� �p�P�p���&,��9��"O��
��ɨW!�4�A�U(c*H�d"O(���H��T��,Y��D�F:�AG�'�ў"~zj��?:�E���O a\}�׃�����0>I��I+
��xW�Ĥ/P�uK��XA�<��Ê�R̢!�� [�Q�^{�f_U�<�ů�5HU���� �V���"�c Q�<�&M�J�ְ3囋�L�2�M�<�D�4�dE1v
tp�EBV�Do�<��G�4e��ik��W���)AF[d���hO�'�n��i �?zJ�i��œ���"O(Ab0O�D�����d��a1ڽ�U"OL�Qɓ�R���ew.Z�ٖ"O���"힆RʌJ7�S�> 2�%�S���9���gi�.�� ��!v�!�, @^\��a��G���񀍮M;!�[5p��C'�]�'�V���OùzB!�'&t���TSo��)�и!!�� �|�b�K(5�Q��/XW��xҔ"O�I8ӯ�AҐ�ⴎ�6Z���"O��X5�^�;��q�%�+57�eJ�"O䄫��.PWN���.t%Dq"O��jD&�"�&R��$�"O��H���Y�HYW�ץ5:|Ò�'V��2=��`Sv)6W �	k�	��H�$B�I�D�ɠ#Jf��Ί+S�B�	�!���s���h҂$�B�V�r��C�ɿm�:Y̍ ޘ�c��Q� Lʣ?1���V2Y�%!$BY��4��0Ŋ�`�!��9��I�F,�m��JVC]�]!��͠4��HHsO1P]�|���J��	^��The��<t�q*J5�����'#D�0�嚉͒�`e��"HT�Qrj!D�y�dX�`��DHDf��*�+'�=D�0��◸)P0����61H�iG*?D��7eF&C{�@�:i���"D�0ر�^��3���//��D�#D�,��صJ�J𤤆�]%����"!�d$�O �0�%@������&Hc�d>LOF�#w��J��y(f�2i�N��"OR�f�����*D���"O(���jP��NP�.��k&�� �S�	K�����㝏���r�2C!�dێ`�6,�B�Q\�r��Ĩ��0!�$� �p���D>z(h�Ʃ�/j!� &\���E数Cg���Ǌ.d!��YF���は��do��C�gL�P!�֊�$�f���eq�E&%G!�DF�,�k��B �I;V�:wFb�	o�'��@äU�j�>�����(l���
�'��4+��)[����fJW�#�jD�ʓ$��=�	W�+���#U�Q�	�'�ў�|bCjG��: �K<Il��@v�D�<ywn�b�J�K�%N4r�|�%��H�<y$W�H,���{z(�-yGB�	�UOj�`�}:��Q�H�e��?I����.�΄rx^�8�Q��!�d��^$E�+؜k�ś�AL��!�D��uO�,��&/�5g���[�!�d�*�1@Zl.�A�v����O2@H�j�U�ZD ���%j�l͹"O����ǔwC؈���/�N�"O<e��-C�=������3r���"O�uJV)L
<b��$f }}.�x�"O�}ѧ瓧B��<9��c`��b7"OT3#K�u2�;��]�(^2��b"O��I��V�iQ,�s" �3�����"OVli5��tL�F��&y�V�Q"O���-V77Ѻ�3O��[ q "O`���`�~�
}P����D��y��'��,�RdR'���pPΉd�R�j-D��K�m��tL�Պd%�2=�"�%.D��P�
�:�L�d�͚9���K/D���);��yD�� $阦�2D����$֬]	���`�W�y���0D�L&K¹sH<!҇��>o�䓑�*D�챵��l�Dj�'Ѕe�FE�fn)D��0vn�53H��Q��;YDDY���(D��e�N�<�(i���Qb\R��1D��jf�Ʒ'�|���m�A���/D�K�$�!l�s%��/|��h*B�.D����Ǫq�����N�LՌ�P��!D�� DhC�"1x�Y��/q۬]!�"On퀂�عBׂ���D�>�� 6�|�V�h��S�~<����#IY�4��a��A5�C�ɜd1�7�O��詢$�%�C��LE"�1��$�x�i�iީU�B��(�U�V�\�a�����(���B�	�*I���HםQ���P��{��B�	=u(da��[[��(`����B�	
V�~����˔
}�`A�J�DڔB�	4�r���l����z1MA	h�����	�Q>��uC��A}j�x��P~��B�I%rf<`���5$5Q�?q��C�I5�r��c
>h�
	ؕ&_ �xC䉭)�F�qLX3uc�0����5ybC��+!�����W[��PO�1C�		zb� ��lB"��6(�	B|
C�I"��
s�	
�f�@��XJ�B�	u�ع��
RI��M�IQ�5xC�	�nY�+3�A8t�^	"BE�{�C�	ɩ5�9a��4��.H�S�.C��7r�����͙M��GO�U��B�I�M�b���@+.0P"1'_�B�I/J�NlHBц^Ϯli�.M9��|F{J?��
�R|��`�.
�ÈP�f�>D�����[��`�"B����"��&�;D�pУ(C�Q����Nŀ7��S��8D��Q��@���Q�*��k���b�+D�4AFƐ?a�p��s�c�!$D��"��*��RR
_�5��%))"4�Haw'�VW�b0���������DD{��)p�`B`���e"w��,x�ڹ��'D�d�vo�_��bE�:d}��J��$D�P���<0*SF�}C�rDI#D�h!	R�*ֈA���� ���5c;D���"NL��jK(	<�I��/:D���#j�Ot�U�'H�/S��U1p�6D���r�²tXk�n9��M�T�(D��S�'��Qi�K'���iG8��d'D���nC�7sVA�b�H2�T9D����\+U�M��D��c 8D��c"Ԇ1���4�Q0��X2�!D��B����+8�i91h��wȆİa.>D��8�G�kW&���,�i*'�;D���qk�#�|8��Ԩ{2�c@�7D���3# �Q��"�֬x�E2D��B�F�RW���V�Lx���0(4D�ȨBI9@������&0:֐��4D����`ו'ð�P��M%����.D����/4A ��X 	�,��K'D��ڇ���,i�h�s
W�_��PB�%D�X;�`y�j�S���A�l|�@�=D�����f�Y�7�k� ���7D�`�AI�p��1g�W8ZT��;q�'D�غ�)�(F(�,Sӆս*�(8ƅ/D��[�'C>Mx��r%M�<��T1�b#D�ȋ����⨉��8�� �bL?D�;"��W�&y�2+�\y�i�c<D�h�!�ɴ{3�]jw��Xi��#ï;D�r��9`�(��\m��H��9D�l����`�c�.P�BQN�M6D�p��fݔI�H�U�Ln���b�4D�D�S�BR�q����o�x��4�/D�FH_(��	8�
�Q�z��8D� Xfj*Q�����0��!E�5D�� $ū����Nz���"C��&�T"Oļ ��"5q��� J��~�"OPeq̒yd����RZ�N]y�"O���f�*�J�%͋�k$PmB�"O@���*�V� �K�'A���t"O)��\�@�޼Y�IZ�m<�DJ�"O��B&�[}*��ǿt8�y�"O,��V!ǅp���@Wn4�6"O��
��?�J� �o�j�e"O��5���T�$M�Bn�?
(5��"O�`��2z��Ԡ�M[��[�"OrY� �Y�:��㔁��a��"O�jW����u�dkJ�#^*|H2"O����En��c�o�x�S"O)�S��H8; $R2�&�;�"O�}�"͇�Y����6cݜY7N���"Oh��eK;#�z���"�-yF�:"Oވ91C�7cP.��D����@� "O6U��`�,"b�l	")� M��l�"O�� &�E��AP��6,�> �"OF� �_4Z�4x�� � ��c�"O��:#I�Mײ����"���e"O��#�R�G��%@b��?||�Aj�"OԬc��F�n��g[�L��HB�"O�X���.��{�G�s���f"Ol���ǡo+�E��  c�x�"OȘ�C�tE���&ѴU���c"Of�ȁ��+UX�2% %�	w"OT���ș�`��de��4�4"O܅B�d��7gX����	�B��"O<MIv����ċsE�0l ْb"OB�� ���4^�Y`p�)U�>��g"O~ (G���X{����ă��d%r&"O�d#�j��-�]����)��|ɣ"ODY;�2d������;��E�"O��Tϥ<�xP1� ���HT"O��� �V�>�#"��M����a"O��"�n!!$ô���#��p@�"Op�
�A���h @�i�4X�6-�o�<�a, %�0\��+��${�)BE�<�1�8Z���e�B�1^D�ʠE�<�� �, �t���$�&���j�nD�<y`	 >��	u戮R}d1�M�J�<I��Ԡv��
,�n!K �`�<��)]�:�x��3!�: ъE�F�<1�W6Ph#��8����m�N�<i¢�Q h���@�C�r�h�H^L�<���&��i�.S��иA	AJ�<Y�`� � �ѐg��@C�(Q�N�^�<	"�G�A�c�&��S��a'[W�<Ad�[�Ba6H��ȵ�� ��DM�<���S�N9X�y�� .��e�v&�H�<qd�ͷ<�Ö�&�k�N�<�sG لqQ$l&+��ʰ��F�<�A�P�b��Ea^IY�p����/B!�D \���d�9@��3"��!��ޣ%�6p�f�>*>�)�fօB!����`�6.(�Zg�D�a�!�$\�<�帠o��j����Hf!��P�-J��(�Sx�D�d��;UW!�� 
�@��ِ	��Pb��P�\�!�^�; �u��D��,ٲ���Oz!�* ��)�C������4Ӛ�!򄔭��Q�O�,-@��ۄr#�C�)� $�KAڻ/��Q�<(��$"O�]20W��bU`N�)�	�"O$I�녜&�Ѣ�G,JE��"Oly{ �ħx�& "V��k�tx#"O����U�>��"�?w9Z��""O�M{�j0a���ǇǠ}4� ��"O^QI`OE�5@� ��k�-r�"O.86A�1>=0�ɣ%"�ؠ�"OX<J�I���F$��.� IS�"O*�`b�ɸf �H%Dح,�4;w"O^j�'�%���1���3}n� �"O���`Y'Ak������teb�8�"O���0l�*����j %bLA�a"O�`-�<x"��7I�h%��"O@�Q�X�eq�a�Ɖ'=�AS"O���!��¡�wϑ�s΅��"O�tR68}ȝ��#�;l�T�5"O�:Nr�T�N�B���J��y�)�_bj���K���rσ'�y2�/����jR�}&�	�0�Q�yR�Q671Y����K��`&?�y�m�MxΔA'A��E�~=q�5�y2b~��=��&�=CR��N��y�,!$c����m
+��PZ��	
�yB���̙&�^uG`�	��?�yl�T���iP�W�ZX�2���y��¦�$�����}��1
ѧ��y��I�,�R�@QF��q ����Z��y���
DS�����J�k�V��Gf��y���!%�ɩ�h�f=&l;� ��yr�H�
�=�7��>^�t���H��y�j�,ˮ�zb��^Tzf��6�yr��:f�ŠVD�V6@@�/���y�$	t�. ���8LP��"F���yƖ4^	@�إ��ѪIGpD��'�h�:UFR8�I��`FI.f�p	�'�n�*���6��	���	)H0��'r�!ۆ�H:g�V諱D� r�p�Y	�'dF�2UϞ:d�ޑ1`��b��Q
�'�<�B`J�Y���bT�m����
�'yT��U�ɘ	*�E�a%�/;���3
�'�h�nR�T���F�@a�`�	�'��Iv��>q�$�q�'61?�D��'�BH�w�U�-�Р��ΰ. D��':-�F��n�V�k�τ1(�"��'�.t�#D۾����K������'�> :Ņ�uƴAu�IX����'�r��f�C/�ĩu&B�VnF1	�'fn���1f��l"q-��I^VL��'^Xrk��.]��\0Pc4�'�����hg�qb��F��Ia�'����d+�2J�h��W�\�M>j�'��8�HY��@%Q���6����'�8�W꒝0B� 0-��1�:�'p^�3A�Ց0��ɲ�_�%��	�'������ɖE�RqүH.,$����'*n,	g�е@�V�a����r�pP��'���H7��1s⌝����$�����'�$���0E��03"l�#X<q�'�8M;w��V��Hv"��(��1��' F�4cs��ē��B��	�'���ˆ�N4%�5ڱ,��\�	�'�.�!B��� M��ƛ� �]�	�'/n�� ��-<j ��ҸK��D8
��� ��1k�L���ʕxw ��%"O�����?y�h�J���nEh��"Ol|Zf��,��!��Hb�W"O���$���/��jœ�w���d"O�\�"N	�R���cU�W��V!b�"Oi�/ؼl��lQ6F����"O��C����FB���fKZ�Yc�"O��� ��;s��X1c*˛Pd��"O�Mz�c�>Z�.��JF  ��{�"OfM �ϙ��N=���SN�2U"O&�DڪY�z�Ѕh� +�0�B"O�@
U��x����*\����t"O���&�^�+^x�A!�*�ِ"O �	��سb���Iv��&pz��z"O*(@��_�_�)f�W`o�A�Q"O8 ���}Y ��E��(��Y�"O\0�Ӭ�k���Ҕ�M��[�"OP�xD/�N<<�t"�`O�@P�"O�8 E�-�Ȉh���%�&��"OH�Ц�dm���v� 1�P��$"O>� ��Q3ܸ�u�M� �h���"O��!��Fd��	
�5�f�[U"Oh�[w���
�J�FK7V��i+U"Ov��� ��ơ��G�J��S"O`}@�k\2*5+�E�=Z�ɣ�"O�9�A�*$�r�� .�4qPR"O$rAE�2,"4(�'����p"O^`yǎ�C:����٦SR��P"O vg�/'��1�ŏ/����"O�U��R*^rR�0 ��	S"O�Q��:�1�V�/!�N��"O�p��2���хB�ppS3"O����A�j������Z�cTa��"O�Ъu��6r!�r�A�MN�#�"Oĕ���ŏg߂�0֡C�e�X}c�"Ob0�#,)0~�����a�ڜ�"Oj�x'<��ʂF°xp�i�`"Ox�&�݈
�ĵ�+�gf����"O�j�JH!r�D�	i�4<c8�P�"OH���J�O^�{MP�9^���"O
��я#��5����=芕"O��J��W�f5\m��+��L�ܹB"O�1�O��&Gt]�P!E7x���"O�U#C�O�z�ȂU��(�T�C"O�2u�
W�R���}��ܢE"O2��bLL��
��‏��R�ha"O:IA�EP="����i�60e��2s"O�����4bp���]_��2�"O� C=n�P� ��AO5<q�&"Ox��G�#vzl`�k
2%� �""O�Ⱥg�!{�\�8�ꘞ2P���"O��3�ޝ0*�\�����\��"OJ��R�W�7�)TIP��@�j�"O��bu�߰|���z�X��"O�}�%�X�-��<��
�C��%�E"O
���!!��a��bH8q^�� "OJ�``lќm|�s$�F�Y�	y�"O�PGl���F�3� ý �:�#@"O*�zc��x����E�BG�80"Oj��Q�9�.�7�ЌD�B"O($Sf��� #���8�0q�Q"O=��BǕ)�<O�t��}Pe"Oh�3D�#8Tp���%?|m�%"O틆#�6���	��3�"O� �|�a�B(l.����	�" ��"O �q#ڱG�pYBG��S� �)$"O�H��?WV��t$ݔ@�|X�"O&ݙF���*]`3��eE���"O�pha���9yX� f^7X�l10"O�5R��Ј5���0EN?�$�1�"O�P#R���n� ���6��)"O�CS �>`�fK3�ɷ)��x�`"O0�Q���H�6��G��W�q%"O������G��r}�|���B��yb��2,T0kpc�D�QA�lY�y�?~YN��3��&hY��KX��yP�QT^�I���uL�t��J�4�y���7^�z̍fT��K�y���-��"V`	c��h�m��y"kD\���9����b稱�eB�y���B�$'�XEHL�E�S��y�B;dđx0lN�J*HA����y�ˑXh�+A$Ï?�jT���y�#�9I�Z��#��&B\
��H��'" F�"ov}�V��3g�X��'�D�+��6r��(��[�a����'�&)9@+^y�е{�GLf�]��'6|���
,vt�z�#�����
�'���(ׅ�P����9�� !�'�Y;��Kj���Ӓ�F�+���K�'����b/~�H1#�)�5 a��s�'� ��`NZ'^�!a���,.`x
�'tVQ�`��*��]�8tHl�*
�'PD���߷?�Rh��
�zWN���'�ly����b��C����@K	�'�����O����Kv�I�x�nEx�'�Ha��C'Ө���X"rblQ�
�'���*�/�UDР,B�x���
�'����Q�0M�,@.�|�� I�'���p#ŅE�D��G�J#t���0�'PHⳋ�8&�&a�W��b�����'�
0��b��,x���I��h	�'�}Y��ͪ&��d��s�L�)
�'������6 @r@c�qG���	�'�R����=
d�-��
�>!��'�1p��;�ll �R%�H��'���。y��ܛ��� n�\��'���@D��E����iM�x����'��F�݈L�hkwm�m�@�x	�'ބ��VK_�CY��yv�>q�B�C	�'������4LB,�DU��X"Ox*¬?#�`H��A�bb"Ot�{�/�҈��'��UZq"O�a��A�*�HǦɱI����$"Ol<��� s[���bOɣv���B"O����`�5!�0�%N�9<!��"OX=*PNGN���띧W�L��U"O�!�aLG�N�lp��@�l�Q�'"O,TP��_�Y
�����)�J�*$"O�H��.Μ7o 9JaA^�����"O��jF6$r�;�ϟ6	��y��"O�8�FI5h� �[Ce�%t|��p�"O���%������0Ik��"O�Ak�I�WB�<(�IL+Wرcf"Ol���͗0l��ay�bӧVP�"�"O`AD������	!��D���"O�+[�@�K�%o���W"O6q�ѱ"n���ʘ=g�l���"O� �ҡ�T���F�Y�Mj��"Oz$*�@A� ��q�$$��"O��i ���Ur��ʜ)>�2�"O����-G����[���"Ob�c4!I3F�lkE:GN�xr"O�dYR����|�cP��|;�I g"O�L)Q�Ԕb�Z*Uf��-�`"O��HPa��,�h����#`51�"O0ݫ-�5]l�p ��J G���"ON�ҖEֻkJ��b[� q��G��y��X
&+�,Rn�R���h��yB�ڪ!��@�X/R�"��c���y2#����τL��mA����y��Y�P��Q�΄@	��t���y��+*�>]Y��%K*B���_��y2%��k��x��"��R�L(r#����yR��6v��qĀ\.4R��E�M��y��Q�
*!�蝎|�Dp�c�1�yҫ��1�j%��ȯp>�t�S�Y1�yr'��m����%���a��+�>�yr�ƹL�"��NT�Z�����=�y�F4"zX�x�C�2W4�l�@m�y" ��kR����JCHբ6���y"�L�)���� �)E�
i��k�y�!/h�(�a��@�J ��ش�+�y�	Ԝx�?;�|�d���y"H�(GLU�Ö0�bx�T*���y��^��5��N�+N`c#&Pn�<AïW&o��8`T�>�Ti ��M�<�3ڍy_��GF�Q�r�1�*J�<	�`��Pu������H��Iq$�}�<��lFSʼ�V �t<�q�D�m�<ْ��+ �VQ��/�Խ Ņ�^�<Q�@_X��հ�ê_�e��l�]�<a�蜕/n9�O��]��0��[�<�,��Y�|�R ���>�ْo�<eaN&�(�!�
>�̫q�@c�<A���E4�]1�ڃ><�xC$T�<i�ߧ0�}J�N��j`�ea�d�<Q�K>\#�S��3qn�I�X�<��=kR�uKS%B�,�z%�MQ�<��,�3$��mF���h2b�
M�<Q1,̴c�����
�q*B6��S�<1R�ѝW��2�e[��$ήWܤC�I�.�\�iDx�:��@���C�I2Nz����A��6dv�Zco�,HZB��8M­p&)� �P`��q8B�	��eK1�ZY1�)��#]�q;B�I�k\Z0/@��b`{5%�'�C�ɴCs�f��}�U��lݯG<�B�I�A2�9�g�(�*hRS��=u��B�Ix����̜D,$@�Da�E�B��3sb |�c�[ u�M�T(؍r�C�	��gE�j��I����&�C��.M�8��0�N�@�D����F�hB�80qh�	4&ƚ}b����=%G�C��.[�� �/C���F�5��C�ɕqU�y�Le ���cE� � B�=u��i`����B�<�#c&�:*��C䉠t�ʨ@W�בV����+I�|B�	r��+��C��J}�ui#`B�I& �D���ɼj:z! F c*B�� �^����$Kݲ����
;n~dC�I�?��=
&�=j2�4�V/<)�HC�)� T9�	����T#�l$�s"O$B7c�2}t0��BC�#xW����"Ov 8$M���#c��JI�50d"O�Qi�
z�6А� ��gH�ę!"O�m�"�35��Z�A!G�#"Ohã߇0Y�Q�%f �);���"O
��p�Ȫ/'x��Ve�w�,�QD�'��d6d�=��W- ?�d"��L�SF!�J�Fh|��c�^�^:" 0�!4On�=E�aҸ!���Qk]�}�Xٲp ��yb��,zrD�$�(wc�dr.:���>�O��"7h�!z�lĊ��_���0�'T���&N8�n�9<��5joD?I!�D�+S����ŬT��.�mY:,!�d��d���d�J{n�[��C��hO� )I�m�:��#�?d�eK�"Onx%8�ȡ�5�م.��9��$,lO�xQ ��	�L��5�>$"O4�H�
K+@��(�D�j��݃4"O�+K�6p ��&cE=��J��'�\�dQ��T�5-t�z���2lO����V9a���S�A=����h+���S����d�%l�\Ls�)�"(ZjY	��!0�O�=��j!�D�D�=e��'�J�!&< riXZh<q�`��F�|yFG�[x�#�Gmx� �'���{�4#Q�F�C@��dݚ^�C䉛�E���ۑ#�:H*�BW�Z��C�I2���s�Z�~y���B�L� �����X�t��h%����r@�*Z>!��"]p���I��ZKP�w�K �'=ў�>=ZDM��z�\��愺VB̄�5ʔt�<����t���V����5bTg���'���p!c��VҔ�C ���7�D��e�<D�$���K�3���)�զ|l"�zH-D���2��>\��T��"G�F-�$"*��1�y��i�"��Z!m7��-���K�'l!�dɷ#�zڡ`K55�Y�tn(�!�	��RS�$]��a5.�?M!��Z�<��PN
��$�n�/{/!��A�+f��@Gc�~u����͝�/!��T��A�F�W�$̠��R�!��X�2(>+��P�Q�<��f�ȿ~��yb�;6���Qc#��8�d��@�12��C�	�(.t��'Z(��2@��kª�O�=�}ZWD�G�:y��6`ڔɳT�]i�<	#�
<8T��pO��C_�0pF�j���=�B"�B)sq��	9/���C�c�<��� ��,��E�	V\9�%Ǔܟ,���$QyV.�;IX�s0�,8 a��?��a`�5f��A��qE~���`��1 $��*�{eGTm�����Y�F����	Z�E�
��WN�)�����Mc�.�^�d�@��/~lH�J�`�I;0Q��>��(]�8��iABW����ۃH!ONb��ɹQ�L�a�h"�~�+��B��9r���Gy+G<�J����� ��c��׶���HO���< �	��[q��1gn��f�t:�A)D��g!�d,�E�Y�k�H��',O\m�~�>D��Xs��=_ ��P�,�=[�L��<9
ߓ[SzDJaK�/r��B�\4X^J�$��A��4�,1��C4(�Q�T�V Z�0B䉣[���p�,=����G�$���?1�Ig~�`��8��&�3.R ��F���?��n����k�&z?��#�ʀ9 � "O� .	��#T�69��C�GPk���1�	�P��>��wh�9
p�	1 ��	�`�k0D�t�a)µ.�؊��	����6A�<����Ӹ+��a飄�% j�q���یUSlC��#4s��+��ѩ;�����a�P7�#�S��Mk�H�I�>���гM0Nܺ��Of��'�S�'90�F�e̩��U)zҸ���4���ʕ�E�֤���(-� ���u̓[$�=�R@ÆDӼ}��ܤQ��L��*jڵ"�g_D*x���8(^�&�|E{���oK�D� ��䞾c� 0i��yr���:h���d�׋Ym���F�̲��'�az"��a=ƍb��A�:�q��С�y� �n�4� ��}}�d:�B5�ybI0�>,�G�Rrs��H�#��HOޣ=�O}4-�Qf�+������3�R���'H���0䒞E��)\&,M�=	�'�<�¡Ɨ��=���_x�8;�'%��˓�Z�*��Fn�<��ы�O���d��7�Ј�6��'��I)�C��Ug!�Dٱ	%��zG�V���l"a!�dJ�m�8'"C\��1�֋D?S!�>?�ne8e�œ�H5�p�[�!F!�$A-P	��&��w� P�BN ~�!���eS���a�7q7��a�.'!�]rv  s��M/�J}	���1�O ���/z�����6[_���e�!�d��KN����#P��85�R�!�$�3GgF1K�̈�eL�XJ��z�!�ԅf�P�����v>-�b���"!�$ól75�낻w������=ma}r�>��)&����բ�K����t�W�<�Ɂ�~QP��.:x1it�T�'��F{��n���4���o��XOF�zu"O�YIV$ڜ%�f1[� *LZEh"O�U�&ܯyt�r��s,�z�"O �� �Z��-�0��M!��"O�3`ܙ;�1B�O*l�%"O�jqDŶ,����e�ܝ}�P�J�"O�`s�L�>xbm)�F
�E��Ò�@���	�U��A¥OuR�x�LχC!��,y���Br	��6l[�L��=E��'@$i*@�{��u��@I
Q��}��'a�}�D�Q�^h�ipr�3n���'�p�C�k zDűA��;#�5#�'ɨYFa��;�U��/R�:�a��'/�!�QF�*�	�$&�83.b�!�b�>qI<a���'�uPSHW$Wk�u�� ��l��y��'�O1��4��d��
dq@�'�<���=|ON���CX����/ʰ%ZF+�S��|��'���M���HbWd�~����'�
��q��5o��qBw�L���	y�O�$#<��+��h$�l�����%YC�<�4.�!J^t�x�@أ <�K��@�<�fm(sK����
�4�P�C��y�<�g�ҎKR��5��0;d	P6�l�<p����aáE�l(�!J�`8��$�P�
o͂��PM�7T�$a�W,-$�p��%t-@'�X�'���`m��(OT�=�O���� �
.M״Pņͽ5�9�
�'E�#��Q�8�X��Q}�m�
�'Bb�MW�y��؋�FąLU �8
�'�\U�Ҩ�4:RT�a��M������'�H]���[�p������a��� �uQs��0Y����
ʟe�s�"O�[��H�r�.Q��韊V�t�2"O*�8W#�*u���ʄ�7q̭��"Oƕ���d�"]x������u�s"O�-��U50fD�x K[�n��"O�]H��9_�B����9`6��*OP���ρ��pP%!4��
�'ȰP�e����G�՜��LH	�'v0��I�
�4$1�n	53K�,P�'TX<�B�!�8�ԓs��3
�'Ǝd"�a�
��i#m�$:r�9H	�'D�Sq�(X��ybrh\�+��p�'���Z�@O/$jH�K�#V�'n���'�v��O���h�ۃ���8�'��0nF�^�R6cU,����'x���dȊ6[�8��E�ڤ`�'�̙E�P
&��|���9q�$(�'w�x��� 2k�@�.���	�'���Z�̀+z� ՛��4 �1�'���e�G�<�����˸bX%"	�'Ofi%�=Ԕ�	A }y�]C�'������o$0���ؾE�X�
�'��Q��ם����T'؁u6.�Y�'�H��b�'.�t�r�`ŖKb��'�^m�f׼dC��y���Aˢ�J�'���{���:�����8E���b�'U~(#���f�1d閺?ߞA	�'g|�!@	�8X4`�0��I-/$��'Ora�箍��蕘���1'����'冔S�N�`���D��vyS�' �5��ة�f�Z"�?��8��'� �F
Й5Q�-���/� P��'�E�7�7�D-�q�Q,�b�B�'�X���bC����wG�� �>��'�r��Ad�4Z��w
��$B�'��@��D$ත�yb���'b�������k�l�rh�~MnpA�'/D�� �P��qS�(/v��%��'�v�q]'U�Z�` ES�f�^t�	�']
إ�:0R�����]��9	�'s`8d�� (�� A\�P-4Պ��ty��#��5Ǵ(�tO�u��d�*�u�lu�ȓa�N�q&�A=]s&��K�2�ȓ�t|� -�.����� 豇ȓ1rAa�CB�� ��D��v�"���`wҹ�஘ ��l�2U<m�؄�r�pcX�`K8��H9.L���_� tc��НFB�5��١=��ІȓH6�8�!��:VTi7�4uP����!�t<�d�JܬI�k�l�Bl�ȓm���"�A�l^\���Ð�9g�����m�F �7j6.�M) ����t�q2�<<j���
����ȓ,�\�I��4�F����Ue�2 ��Vg�+�6*�J��&���Jm�ȓO&����M[(&y�l9#�]�Y��фȓ8�Ҩ(�C&;��)�2��d����ȓ{�f\Z���D���ռ~22��ȓKD�&��390鋗�Z;}B���h�řq��\aE��D�ȓs�� ��-_���K> ���ȓ�T�JfO�{����d5&��<��c��8���U36��K�/�,'�C�	�;�x�ju(E�d��p`U�x�DB�)� d�k�ɜ��|�Sg	� M~d&"OV�P���8Hu�䀖%r2I	W"O�����v��X%��o9�(�"OPp���H�lđ��� w�%�"O�����-[� ¡�34��XQ�"O��Ad(�SSd협�؝9�XY�r"O�d�tE�#�
	ڔ��=.�X�""O<�@����F���j`�ˋWyF0Y%"Oΐɢ'�7��h��~T$e/$!�dF�b�z�x�W7Y��Y�R���P�!�$U�"�^A����%�b��!K�a�!�H)I*"��uN92�ഹ��^c!�Ě$zʲ)�Tk����cV�9r!��+�X�*5�'G�`�Ҵ��fz!�I	߸ ��$vi��B&��;f!�@� X�l��qa��k0�.*Y!�$���mN�3��1m�%4!�$�%�R�Y��̜v?F]�Ṙ� !򄀡lM�щ�
ΌA��0�@@��O.!�$S�U��FGO�wc���ӯ	4z!�D-8�p "a�F���(���54�!���q�8���!�;Zk��Y҅N1Y�!�$�|���PS�)X%X�]!�Ć10���&�ĻL����2,!�d��Q�ْ�@�b���hÔ:�B�	$B�m�sH�ø�J�O1#�B��(7�M�C�Z�I�r}�#��ZC�D�4�wC�
+�t��1,;J��C創|�)��M�e�~q)�:�!��k���)�b
:"�lA#��A8!��ع^������ĵIc6�Y�W�k!���1����!�(x�d��'�0�!�$�t�.�³�P���a�Хj�!�F��a���J�'���3��K��!�۫=�M(4ꙏ]�`-��"ȓ�!��G� �h(���9-���aB+ńC�!��1+;�\ [7D���6��\�!�ރ^|�]s�!�v=vij�!��
1R�V���č�PJN9��S�au!�$I�*���j(��ev�C
�!��<e3���R���H�E�9�!���&r,<���ĺz$���Q}�!�D���P�Ё	�bs��*!���<4�ܨ��M�$6��CZ!��"_� )�lCT�Q�[*20�	�e���r�'by�6��}E0��U
�Q�	�`�VL�E�ڎ��A�T��M���ZFC��T�8��J�<Y�"�y�z,ׁ��>�l���H�;��b�4uS������2P��8;z�L�ܺ���aW"O6�Kb
�3o�x!B6k��HT�$�9&�)۶/�e����I1O�Q>7^�pKHM)� ��XBV�W�+<`*�$K��x���Zz>=+aDLd!���Q�=Z�0��GS�A�X�!�yi�I�aw�L9s�|Zw���*�$�3e!������X&,�
����h���=(�h!&'Vay8=ㅍΣB=~q�w���
u��
��S3_��(�׆~�<�O�#}� hƝ#��)��oߙ��ՙ�%�d̓�����%��
�r�ybݓX���9Q�:������(�4>ɚ�A$����Ѯkz�y#ɹ.axr ��5��I��ǧ\�`�Q��$	 2�	C�ɓa%l`��6�r]���)פ	:�9��
��9�T�6{����u�T��2hl�Q-Y�Z����g�L�����Æ�݀�AaE�xw���,L�_5lX�q�\�ّ/Ozŀ�%�bu�)6L��(��QTfR� �V��dC�*��qA����NmH�'ܧ�� ��I%�`��$JzU
Q(�pd��1B��L�T˓?ιi��4 ���PÂ�	����O�b��'��;���?g�|�8��	�
98(�@�ؾ�wfYP��&I��-�+=4��ʓ�*M�G Ǯu����Ó ��� ��m�t�CC�1**K)�<T`�v��81��$���!�q��9H��Y�K �� ���#Ĵ/Wr�`�T=�Nl��	�81��A9�J�+�(��ET��[ĨP���#q)�?�H8�E��@�m�K���N�;a(��d��p!$	7��-�8�"�F6�&���+<O�0�r@�2�2��s���t�0�%�tTi`G'�}aA�F1]�v�1�A�r|x�H���3BC�)��$?�����b$����˗�V�.�q`��N̓W�&�A��	u��i6YZ�vQ(u������'y���+�X��X�o����'�
1 �*�9/!�y����Lz,�Sh�<����9L��t��?�ZȠ@��.|�3Dʟ͘OȊD���
LH<��a�q�pUI�\�en�0+�'](������9���7�.)Is%�+>.�1`�_23�fl�Ш�7]*�����Oh�W�V3U22���l�59���@��')�  �N�t0�9�E,�"�<���ǟ�fuʕ��M��K��0�iS�Kq�i9&�i��	DlQ�Y����e�R�4��!sd6�	� ����G�`=�7� I=��SRG̐��4�؆H&�,BF�]�M��⚃�yR-<jM�U�ٜr�������g���ړ�Z���m52}>!C�lX?[y>��9��i�@%.�qj�KF/�NC�	>7gz�`5�Bz�j��lM�<�[#�V�" ���VQ?��9�l�����_�TJ������7,�~>�{R�J�L�ٷ�K�����H'c}��F�&r���an�O�|"����>�������c6b�ʽX�� k̓b�ȱx�΁)KV>e��>qɟ 8��M�p�Jdhħ[�s	
��R
OQȷ�	�m
�QCF�ɭ)X^�����,cϒ�f ��gq��'Ĕ#}�ep�����J?"�S4.l�6u��/I� ���B
QU
�  4���<�h��A0Ra{ү�� r6eRXQV����bC�[����d!.$�em��M��̇�G�`PS��/�jp��Q�<!j�o�ȹ2$�*P�4�;ņYv�{����n�$ �2#}
w�܁Y9r�)&I!H�h`�C�XH<1g@�z*��D ��HIt�ӞQR���"�IM �I�E&eEj��~r��0��0��*9� P�C�;�yr�Y!N�^p�C)u`5���	�'���l�:ԀBGV�zY��ir�		Z�=�E��n�գ�`+�����V�l�TH
bbaN�ժ��H3f1yf��:Z����D=R�����V=-��9w�_��APDF��j�G}��w]D���(_�S<(�hT�p�[+m�(�C�f��X����d;�ɫ7A X)E�(�0�EG��˓I]-�@CA�pҧ(���!��<I�L"��G�tl�B��4�S�~V4�����xB\i�G��*���O���@��}@8'?�p�3���@-B�2-\�f=��c�d6���Obe�
�"tsX��L��F����F�B�"���4��?Qg`���||���|��i�f*���)F|�,�>��殟`��r�v�x�L` A���.b ���$$�ɛ�t��1��5�4\�B�Ʋ�{���� �H�ҧ(���A�c�*���A����y
0"O��3W喭&�:]��ɕb����Ti:��I�`����t��*;&h�U�[�j.%j�K

M���dݺQ�g �B^۲*�8:r���훅�x�^��(0�I�!���`!���S���O@l��)�~[���aɏ�lft��'�� �l�UₐKФ:O��0A�t���I��1@��''v���L�xˤ�R�-,w�aӌ�$�OH�����mڦ��Ν;4o򨪱EȦ_��+ab�	B�!�ϋD�p�G	U��mHsA�	��������q.�B��y�,��:�l)x��Lw�.IB'�:�yRNJ^�ݺ4
ޑru~Јaσ��M�«���'���%��3�G)��2��\2��dw���'q|Mdc^Y�LA�� �2�4�?�	�sb �	�@�zU��ˠ����=D}2��x�}�桛��r�*Q�C:I!�d���x�<1a�a7\���bң:p"q;�(U{?�����&��e���ٱbwD���"�B�ɩ^���Ke�1O�$�ӆ>
j�B��,�,�Qm(5lM����\�*B�Ip����F�"��%B�Z �C�ɿ�@��V�^�.��jKA��C�)� da�q��=�D��Sh�(&"O�E�!\�,��,R�00nF"O|A!$��ռ]󵯀�A3��P�"O�G�#��l�2kL�X,���g"O�PI���U�a���W�d$��`"O���2��}L�<A�AI���D"O8�G�Q��H2� 9n�9��"O|�jT�� nV~�#�ǩy_�L��"O��J$�ڧ1����d�p�]�"O^�����4��ae"�o!� Y�"O ���Ć�͂L�҂^�k���{"Oܕ���	�y����%`A.B��X7"Oօ2(D'h�1�7��>��훗"O�3G
�7��[�/�=a#��&"O*�0�g��:,)I� �"OhB��Q��`��B#��h�"OP�1�Xt��]S�C�*�1p"O,�cE�]?���c?�Y�F"OpUP��ޞ-'��ّ!�9�5�'"O�0��G���u��.H�i�"O<Ћ��N@�#��cx��"O�٠�^�A���BA��<N����@"O<dS��Y6�:$�� �6<���z�"O�QH"�_�,�y�o�J|Vp5"O&����<�Ps�� �L(�d"O�,�0�y�N�"��A:��5�"O�6/�8��x&�ݘo�X�M:D�xAWgEQn�2w���5E� [��-D��`P�Xx���M�������$D�����,�����l���lps�f"D�D�B%�5�\q�t�P3r_�TP��?D��ȆT%[j��]?�h�Rf�=D����E��p���+��7?@$óI8D�8���'��a�CP7����cF;T�􈦤�=�(�^�/"�a��"O��0�L�77���M�7<,ly�u"O�i�CF>|��1�B�I��e"Or0�q��[��+��ƈ,e *�"O0i�E	u>���E3��]�U"O���4-]`[Z1�6͏ fH�""OR\he�VH��}�w��eD����"O�؈��C@���7&�>����7"O�h�A��ڰɧF��<��]�"OR�	#)Q"E�j��`�Nc��D�"OtD��HRvؽ�֭�)䨚�"O< �T��K�� 2�ö?�}b"O� ;sɔ!:�3D�ƍR��v"O
����ލE�
ԹkE�g�>��1"O0��#�2�y�e�ܖJ��d�Q"O����O�*0�6�a�̸�0�"OZE��HFwh  @�k��܀C"Od�`�U�h�R�!uΟ	�.h�p"OtCF-h���L������"O��h#gSN�P�!e�%Py��p"OR��R�*iC���.�5I�ލ��"O0	��j�)#l�ܣ�n	��͋"OvH�s��4����@ʘ�M�.���"OlIc\�d�P����JU��)C"O `��&ߕ<e�M"���(�{�"O���P' �>?��QF�En�̼��"O�}3�e�6Qx�ͩt�)q��<�$"O�M)���/B
�(6b��0�,0'"O��xΛ�_%z�� �n?p{"O�M�݇#f�a�&[�eK@�d"O� ����HϾr)���5b��"Oĝ
�Bn��	��#ڨU1�8y "O``��B0a�v��6c�!{[����"O��Y��1�`��<�|��"O\uX��}�,)��C�X�*�I�"O�rue�w������R��}�""O&� �cQ����d@ߪ{�B�r"O��)��!W���T�WB�h@"O��{��By���B����`��"O2����Y31�L��!�>`�"O��P6ꕷ4�DX����K�*T0�"Old0��J�%�z��q
�z�|C!"O���e�T�2�բ�Y�!���9�"O恰2i31�"�*P���u,���"O�!��ETU��53$c�"yzpQ`"O,�q�R�2��A$6�ô"O�1(��R�;q��GG^Y"O޸pr��)?0�H��m�B��l�<�C�E�8DDk��^�\�BjYj�< ��'�<bb����Pw�N^�<���7�p�6�NK�I8��U�<���%*��K�۷��k c_�<��¥\��a�d��&&i�e�D`�<$J�YbS��Pj��'@�<�c�"�NMj�hB��ۀNKy�<��݂.�<Y�`�.H�Gc�m�<a� } ��Q�J	k���d�j�<�QВ;���0� �bMR���x�<�g*�>_��z�Z�l�61���Q�<YO�Ts~�8�e'_� �+���D�<��C� x��M�f��[��G�<�c�V�[�u�@�F�t D��ERC�<iUn�9�LثW�܉�N����t�<9��ɳ#�X�c��H�f�E���w�<!0�]I�����0p��J�<��.�#f�l �m�o�L��fA�<�s�B,Q�0���
�1G ��4�YW�<C)�%Y�p�NR3~�xҁj�h�<Y�(P��p�H�-{$)�*NL�<���X*�$q1	E�*,��!FS�<���R(�f<h��'��q�t��k�<�1K^�F8`P`�,x���#��<D��h�C�\��:Ti�7Ӓm9��=D��0��O,_����'T>SLi:T@:D��e�F�F%J��S)ķa������;D�Dy%	��:��بT��Q�ԅ=D����K4d�8Xr˖8q�"���i$D���tbP�1���(�dS�g�z4#D���Dj�(v)XE��d����!�#D� �"i���pA8A�բ@k"D���lS)
RnE�WM�
�P�;q�'D�(2T��+ϲ=㲅��0$�"D����m�� �.����ǖ(=6İ�#D��P$�77w<\��V^�>����5�O\�pd�`���F�1F=��Q¯�9`���a�'��A`�N�W��uo�p���Y��d�IpP��ӈ-�Ӗa���H�AR������3����DN�`��� &�@$p�e�΋^И���)�c�
LWڗ�P�%�9}�SLW`4� E vtP\�`H�D5�#?�"#�)-
���b���&Ŝ�[���o�-X�)�(u H�kք��U�H����.=�=��![#|�U�@��-{<�Ɇ���m��|����B�/}2Ā�(g`P0��T�F��c��+]�T�Z!F&��(���gg΄cEk	�঑h��a���+XM��P��"E|�P��04k֥��T��;2�V4Y�ǟ�q�8�JT�A�I�F����:#܈;� �%��M	$`�
����L.l��E��A[nӊ@z�,����vX�Dr�q��h�!�a/��I��!�D*G㜱j���X3�Z��4lt@��b̟(QrP�	r�ƥSC���!�m�]��2��q:� ;�a�t�jV(��P��*D�s�h�5M��$����S-]�[ղ�ns�'"�je3�(�#k�L���dΚ�ʄh�a�7q� )�hԿ�x��1	�҄���<���С�)A�	�Po��q��A޿F* ����g��I�a����k��I%�ׯ-m>��%gӡ?p����+�O0��b�U\�؈C���3@���# �10d���iM9��9S��; r�'��C�4s�O�����C�EN��]�@a��	��8"0
X�#�z��"�
"��4�ӡX����(�M��g�M�����F��!��,<O
�R͈!\���1�9?��"5\��J�ԜB��$��ճ`�\�}�e*؁2B���E�D�d�DlaSh�PΰQʳ�6T���5�������G� ̠2��K*X?�Qy0�>Q55�gy,-/(D�&K�0��=j��^/�yb��u���� �ë�,���KիD�$�b����2�*�j��e��%�Y�(A7"2`��	;Z-p�ɇ���#g����
E���1,�*~�!�ݭ!̀z� �#ka���1���
1���	�$�Z�.�q�NV�(��N�3�"H�N̆}����$���y���y�P(���"Xa�-)��:+�ٹ`JP��=��O�QͧQ �<�dj�zB�YI+x�x�	���L����WHGSb��t�i��h�m�!������3y�0+�<ӢBq=�O8�;P�U�b6�� ��&Tp�[�DΡCX��`Z��H�^��☡s��q"V'+8u���"O(��oq�B݊aI�Jq�!R)d���A׊Tm�D#�g?Y��A�<;z5�e�Z�z leK�g�A�<�n�
��Q䇂a>��I��8��m�Ij4P0�'.1��M	��`�7���\$:A�x q��"B�w*7Y�a�¤�9��� w�ɡd�!�$M4X�N��W�0!��H

h��OYq�m�$��x�����<�@ܑ�d_#bN��F�E�!�>Ss:=�a�Y�sd�ZgF��;�l�EG��*g&��tg���p��ؓB��th$��`R�ȿ�!�d�Z��hAu���x1�T8O�T�DV���N�J�Ӕl%��gR\8���X�ab�4���;}���	8��ؗ��I�]c�!8@:T���:�΍�]�@S�aOx؟HB *N)�	HE�N?;�p�Y�2�!�4� �`�9���`���/�t`���`��_���"O$�3!.�D[­	�MB�"A�ܙ6T�d!�f�5%�9S�>E����\��H�0����녹�y�)���9RT$D�b����D���F�'�@�S�E�H �ϸ'o6颥�ֆ	��q��[,�r����>j8��u(�����o��K�d�� �)z��!� �+�O
`���6 hћ�N��{��1G�	�8��o�;��O���"�@>?F�ţƭV
����'�65�B)��P'L)vly�!+O@�`PE0nv^�J��|Z��[#�X�2�m�2&Q��P�@QW�<q�"N�iF.5Q�ϫ5�d��'�����5�l��w!K�g̓e��pz�Dý@���0���z1���Yy<m[R/	���X�*�"�Q��I�$��B�I"�l�	w�r?��Zpo�_�pB�	�^���@��T7jfp��\��tB䉀��D_�L�}�����.B�	&I�bC�!�c��V*[�pB�	�L층�2�[l�DS2 �'[�C��5Q`�����СH�Kr��C�Ɍt]��DO�t��
Ө?��C�� *#<�{�'Ĭq`��cȝ�N�B�_~m�҈A���S��X�,*B��pZ�&ݧ<���'��(�,B�	�G;�l�a�X�(QщN�2�C䉼.�yA����98%�6 C�C�IcA�%�d��69Fy�t��
�C��v���'�=�,��S�N�B�)� ]a7���$%h`�fg��WP����"Od�SAŉZD`�藇�kS��f"O�tK�)WR,��LM1!H�\K "ON8�Ѐ��l`���j�{��E�"O�U��l��oF�<����h����"O�!���.R���qt�@��ۇ"O�0If�*qA>��F�M�_��yg"O�l{Q�Ҥ)tA���B~kF�ѳ"OfL+��L��R&!�@�G[��y�&��/� �)��aIb��!��y���PX{#��*QԎ�3��^0�yb�q�n�F�šO�<�`�^��y�B�X*�ٖ��6ikb�����y¦� 	�I�7�ֳ?^�"g� ,�yr�_�����SA�^�̜���L��y�	9~���p�^G&�jE�ѵ�y�����5���"�0 �k\��y��I7逩 W���^m��R��y�B�y0����	<�<������y�aƸl���{U)�1-�5�y�HN�_@8@Q�<kZ,xҦ��y�e����ف��]r�̫�HG�yb'ֽk�T2�H��V��~�n\��'8,u��$��,L�`��qX$���')�5;EB/_6$�3/�l���	�'lJ��b�:I*ĩp�ڥY~]p	�'��9
vhR�}{�i�a�j�03�'�M��  `��]AW%W/o���J�'Z*)�l��? ~�)�&g�n���'��9��V6f>���&AߑT� �C�'2vd(U��
8���[��J��'�6`
e̝��ƹѰ#�9<�,�3
�']�=Y�	�`�q+ЂV�<�x��'0l ��ɏuu�͉w�D#0i�I��'3 ��9?��v���0oz��'_���0ѹz�:��d�T ��'��03u!_�C]PPE�ߨJ>�A��'�����+/\�H�T�B�NhS�'�L��'mO�6�����Ak�&m��'�����	{�v<bQ
d�f��'�X�bF��Pwv��3Gd�����'���c��!a3�\�'�\K��a�'��`��&��R��2�.U7C^�|��'
\h��#BJ	Z4�OjW�q��'�$s5&�
%ټ(�fcӮ��'C�H��{���ŋ8�� ��'��mZ�&{@�Fœ9'��i�'���k�#*�&}a�,p�'��tBFF.��v��u�$��	L����Fұ4@�F�G����L�7LI���ȓQs�\��E"0`Xv�| �M�ȓ*8BC��F*��t�!�]|\���qb��Y l�K���A�ȓlR<}!&Ţ{���H�|��Նȓ|�jIA�Ϫ��ɗH��|��\����~_� �b��?_��X�ȓ6�Р򧏕eO�yiGȍ=e��8F��S9���H�Һ�U��bB�#���}�c�5��O�R\�ON��Q3Ո������"|!^u�*OV��JN<���XM��|J��W����G��|IT�[2�AΟ�Pe�y,��ה>%?���4a*4IP
Ox��ç@G��@�)��@����g]=~�II>�꓇�(�P���ߺڞ����B�<}i�R� dy�ޒ�0|ca]����6/�9�r��� 2�K@���o�:����+���|�H~v.����a�ٟn2�����S8b�j1p ��)ۓ͆�l*/����� \���a���i�ǃ5��J�O�!mE�|0v��$~�I����ʧ;�zH{$�7I��%	�H�0p��+g�l���'T���Ԋf>	CoωH\|�%�)T�Γ0v���I-k���M��?��BӃM�bM`'+�,2F>��P�1��&W�-�ᓼ>0�M`R�C5M���{���g���O��[��-�)�+8F�Q�3�Ly�\$�TR��I�c`�؃���S.u+�q(�%�j�e{��	�/���r�b�0]�ɺ?Jh}a��7�g}�T9&fP�Z7��8B���q���s��#<�zV�λ��<���BR�5�`�C�e⬫��v
� �&���&Q�a	(��[�X � @�?