MPQ    X    h�  h                                                                                 slI=:�	��_X�D��l����Zm���,3h��D��/�|Ib�+N��
v�I�c�?.bӡX9@be9�J]3Q��un� �w�م�BJ�܂qw��n�O�t1�m����F�ײ��=��S9&�Yݱ�]]�����R�uTbÁ�Sfǧ�9��㎧�t~���h�^�j��
aA;����ȟ��F2����\q �o�1 >�p�|�,��:�VO�`�!L�o��4+c"2+t�J6SA��e��%g[?C��s�h�� @r�nBtI���\���8�@��N��x�w��|�G�6*`VT�衬+b.[S�a��~}��N��
c�"i-�dG��WX3�~T��[�@z�~g
�$�nlyie�x��F��٪��g@P����|x�B�,:Z��$�o�97��U;�n�l|1⢵����{<��m/lh���Z��;<�=�c5�O��AS?#P�2p�e. f�T@(�ěW�,�gQ��-�+�&\%�#ފr�̐-����ȷ��v:���{������?2�C"�d��h>��;��}��I�(3���1BM>�/ -ϥs��4�_�Þ ��ͻ4.�(�� ��l?'P���]�:��1�c� �M�%�ٻ�

�s�ג�uG����U?'`�F2\ ��~�AZ���V>`K=�_x�v���#�e?�[�ڭL�r�ݨלl��j�2A��ޡ��ZW�������뽠�
x���z��q-�}�L3+ج�vV���<���~1#�X6g��N"]�W�9f������2��DP��B�\�Z�T���1��5:kx��C`x�c�P�/yRK����ZY��u�K.��F�:^��'���(YWwku&)�d��xʆ>J��qyw�ĉ��cZ�f2B|tB�gx�C�6Œ�QP}5�(�>�*��WN�yp<��F�:���v76`�v�w&/����;h�<UҔ��O��I8zJe^���x���Bk
��LWF?�@�>��j��:(o# ���*J��dQ�t�`�ޤ�,v���8NΫ��e���VI��Kl�r���x�!���= `@��h1�A.��P($������B�{ i���-�ڢ����9�)��j8 ٢����N\�������(�ֺ8�y5�H�bD��-Im��w���Q��2i��4��&z���8�d"ˍ	fD�jq�j�&�z�e��J�C���l����&����ƹ[�Ƿ����0���LsH����Ѥ���[�|�n�zI�ԉ�ǫ�F�As�<䰰tW��_t�Zz=�5��m��v�f����a��[e�3��>t=^�ќ\K{��v��z�������T���R���j���oH5�L_�{�k�s�Ȉ�.q`�X�bB$vv��U����z�>Ā����V����`�cg~��6F�t����NY�s�jH���x�,��s*q�pB;�Ƅ]uw�)�S��p��g`�N�8Q|V:2���`k��P�l�ನ��h�p7%���y?ƙ�U�L���>}a&��
YY�9u��o��D=f�8h\S��O���+�j�z���8�(�ad*Cj�S��a��tp����,��& H�vz��U�1`�\K$6�@|�|��H��1PN�Ms;%ܣ��ڸ�q�xc�4Q~�'_Q�a�.RH���	h����)o��N]�9?*H�z��/��^�c% 3�K�~���m뿾�a���KxT"����	O��%M>洸��h�~�#��W����f�<�9*�uW������1�uQ��j� �$�cSG6|l���hkC�\��`�M��ԙ�,y�X`��Ut��." ��p	� 7���t"�d����0� q���g�W	����A�KM\	��X��&a�v�13��NQpC�O�5)7n�X�W�򾳆�H��do#��d�j}b�u�z��}�z����ᒋ<��dƒ��>upqkWrY��%o9d�p���O�N㶾���Ϩ�6G�w��]Fz��iW�r�~^�`Ց{zV�
�<'��:�'RTv۔��Ç��c �޲ӆ�p��H��JyL��Ţ����*&/{��:Z��=���WON��\�/��M6,?ii�-f�#\�hx�*ͺl��_s�&;����Jw�H5� ��"�(լE�qd2���Z��C��@�X4�a˦�v'�dC��4�;�����|�A� �]\(���OD��'�D�Ѡ7\� G�b�/� ��G��|��n���Q1I�RX����� �n^��0�٣����$i�΋����d%�拱"��M5���79�/����`"��M1g�~D:PH����kд&�xb�
��!x�M0C��B2qF=����{�״�����䄆t<ư?�Gu��&'s"/Ϝ*��Mg��I��_+n�E����Xr�Z G�Y�e�H܏]En`�Ze������3$���a��S��[�L��~�]p�r�o���`n�ej�;��t*Tr&c��@̥�ÿF��;�/�u����V��k��3Z5��uѫ�"�� \^"�e�hY�+ +��ׇ��VD�#�hS%�
n�	ǡ�M}�]&L���J�Qb����󸘗O��s_����F�`X��Z�M��ĩQXW�Mk'6����	�Z@�� _�Y0.� lfݼ���F�
iy�h_���C$A%�"�x�:��|I��o`�K�0���J�X�Mr0x`�28<�%������{�"�����h��۫7D���v�Dl��������KQRT�m����A��#9�ݗT�:Gy��#�ʳrj+0RD�=(D
��B��WsY�j�h'�g歺�~j|@�W���W��s%�D��z0btb���jq�)��rE����"�{�����,3���c��s�J!���+K�	����ĕ��71s�)@��M�An�V�}�?���<���d�����)�L3�J�V�P5�g���<�.p\¨�${p8��>ă"�T��}���ޅ��o�mmN� 	9Q!�{��Pu.5�Y�8cTh���i��S�̭w�$�k�JT^ن���~ڱ�$3҂NC���%���?�����S����
�.K��n1E�T4���]n���T�Ȏ��;O5�S@f�U%�ӲY��f�~F�����d�\�MZv�wr�1��n�,q��޹��u� ��x�h��SjgK<����˨�:P�F-�zµ�����x�o+�:>`[u|s���,3VJs�|�5�*��4F�2�:HJ鉌��@m�,[:���L�h{�@��$B�Z>���ޑ���ӼV������x�y��еG��;��T7P��ư�.Vu�a)�}�lj��
ގ�"D��d���W�z3�k��+�@5�L����I��i���xt�����8���P�������KT���,u⦄���j��9�d�U���a��>��~[S<w8/c
�Zс��E�~�3�s(���A��~P�?�`G�f�(���r~��o��u����\�R�ޅVd)0�-hXA�4nQ�e���F_���`*��}��2�D���hȃϺʶk�}w�0�}E(�6ڦ,��>f�< �Is�9U�ږ��zK��D4ɠ��e}��#��ڔ�������[�S�������
���Ȓ�����?�^w�Ul� �k�~ ����^�ĴK4O"��Xcv�|��^Ǭ����S��n�:�c�l��j^x�_y��	Q�){Ɠ}���{�l��x�͚z.n-��ɇ4�G��V�B���аC�i#�Vs�M�N�d��p��.�f	���y��i�Dk�?Bmi�Z��朿�>��4�k	�'��T
xN��P��R�'x)���{ݰ�q.��:�jvň}����W��&�d"! ��^>E-�q�����8u����2ft}K�g��C�i��#P8"(�Ӟ*����2�'y���}&������`�:Ӓ��/
16�[�<�i��<���H�I�bte������D^
��ZLC�&?���9j#	(*�� �`ND����rQ���`��Dޟ�mv@h8	�	*O��1=��lm���ԢS!Z�=��4�锸ʼ�T���*$z�&�܋�BB� $���H�+�����!)�I8�R��dN�Q�[4ǃ�Ȃ�Q ӮT�)�D��c�(�S�(b�e���Ţ<��uƅ��@��f�ˈ_9iYJ�%2���?����e�4��7�6����&6`{�a[9rX���]�u��	�V�Kk��tN�����*|�nz�_����a�Ĝ�F>�<*Y�zc�/y\���%�ս^=n��R�r�t%�f�������R�3֝=��{�^��ܜ��/*v��ޡ;�� �T�#lRTEzj�I���% ����{��-��ÈA1�`��b���Q���o#�mjv>�c��K5�����{�g�un6�="t-��̀�NTby�ŵz����,�̿*�CB%߄�s=w���S�֢�{`[�y8l��:�0��;Oz��Y��n�����+bp�S!�'� ?Ac30ԄL����&�� Y���u\;%����Qq���\�OA�C+�D�zT��8}Tm�=R���. ]a$)�pwV^��в��JGHlF��������zV$q��|:Y,�C,11��+M.��ܾd��3���S�4��r'���\ۉR�O���}�->v꤯��)��9zu�H�-��*��^() ��\��@���v��\����T�?h����	���%:N�Ӄ������?�����f8�7a<*�����[���0O¬�u,�a�֖ ��V�^��6�_��w�k^�D�H�ז(���,dL�S�R��y�龭��J���(����=׃���nY:$�15�����DM7[��=�����=v��y����	�C+�s��v�n�UP�����^����ڹ�a�Ӽnd`+b[!zl3}��L��T����ڿ㈘T/p�KJr�h%J����8x��VdN��x�L5Ϩ��/ ��w �F�wЄX"i���^�T:���Y��ˎ<BMM:#��R/ϔӰ,�-ԗc�|��.%�p�v�H��J����d3�!i���&*��W�E2��܃�O�"4i~�\&�ִ�5�6'�pi�!X���Sw��>S*�v�l�_J�;�����nH�� �Nh"��Շ�:q���T��}�⊭X������'U��� f4�ȯ�'B��2�A�@]�|J�����ҶD'�
7��:�ǎb$�L J�p�2��K������I%�X����lUn�a=0�Dc�����:��f� �/�d������K�5�NI��0Xª��ڧ�!]���?C�`�:�i���J����M҃߆���7!�*0�7R�=�"F� �[�V{���/k������<a�c�B�O�"ݑm�E���J)������s����(�>:����t*
��$�] ���H�/_M����_�� S�g���~�~�`���
9}��b����t���r�܊u���h�ፐ�6m������b��! �]�5c���T����^9��m����/�+�5��g�V�֔��8캀�n�C���t��L�6�Jz�sbhJ&�.Ci��fsZ4�of����X�9Z[ ��4����觢6�P��d�吸���_��.�l�}��s��F���yVc7�B�$\"^"z�:c�i|��o���K��՚pmX��0�H�2�f� ���:�o�Q�Mϖ�c�h�D����#7���m|[D��T�4�%��WQ��+mt��������f��T�CG�x#���r��$0�HXљ
�M�[��Y�A�hR�L-~j;@tT�����w�����t���e��)��E�H�=g�ґ�T�p�.,H }52�����J|#�>�$l��z����4�1��i@;<a�Vy�z^�P��A�6�j��Ů��,L�q�Q�sx��B���|�����u�~��]^d�9M�";���8P����#��{m)X	tjO��!�ؤ�.����Ow_c5j#��Ӈ��\g���$�r��Esr����9�I�?4c��gS�����+��ώ��=����ڂ%��7�bސE����AJ��D�}n|����J�I�#;jp�μhfh_e�����S4~Ap8�X�͋ς\���Z�r��T��jk��ȭ��^�Ш��nh���j�[W��'��UF(��՗ޠK>+�ho�Ha>;fo|<���pZ�VET���埥�Ó4aI�2!!�J�b�/(07
[5;H���4h6�S@�kBj����"���,�n���yƶ�xU�K���G�	�Trמ�a�.Q��a^��}Gj�J�
YVe"{Jd��WQ�Y3�x����B@���H3��$�i�7%x<���ib�;��Pgi��8��n�O���),���Z:e1�9�fWU�g;�f�����Y{<S*W/�}U8Zm�'�w����f�AoAɛNP��[�tfz�>(�@���Y�]�T�����I\[C�ހZ����-#G��O4��iҜ�������xh�2\�'�{7�Ȟ��1@�}RO)�\J(i�z�'Vd>�t) ���s����U���։k�Cpf4d�n�����"(��O�L��0x�����얀m�[���J=
S���M�ˠ�{��,VU���� "s)~���<L��iMKO�ϧUY�vь,���Gu|�����\��l�E�j����:4K�Dg+��Xm�x��Q,�'bVx� ]z��v-�^$��U���wVמ��fӑ���E#�t�]/�N�#���I7��Zf�0�x�!��;VD��B��Z�������5S�k�3�X��x	��P���RA�aS�j�н����.�A����,�8�@�0�0Wm�@&��?d]nƼ���>@�q/fF�:O
S?9P��2��t���g�#^C���gX6P��(�'*U����y���|H����,җ`z�ӭ;Y/��w��mW<��Δ�*��1�I�je����'o%��\
cQ7L~)�?/b�4�xj~:w(�5� /L)�}̵�?1Q]P`UAޚ|�v�i�8�H��2j��^�QArl@����q!���=v����7�-�խ$LM����נPB��I ��c��ژ����f)*�;86R���DMN10�������e�/(+��DAk��#���l�   ��,颷u��P���!���H��˃��Ď�������@�p��en�X�DĿ���A&����o~�[TU��"�Z�\�D�w�D�����Z�����w|��Yz?� ��ry��x!��%�7���0ְ��%���P��=I�Wٍ�L���f�!q�����^?3�A �4��^�ٜ����cav��9��ŋ�zT˲�RϷ�j^$��"����{���)C݈�S`2-4b83,ox��w}�z>�f�֦�Q�;8��H�gt~�6�Uth���a5NO0[� C��M�U,��*gaB��g�ӑ�w+ՅS��7�h]`��8�Җ:(������H�	�=�Z��=kp��F�B�?�L��L:��t��&�3Y�iu���f����\�]O�+�>=z��88���9� ")�	o"a_sgp�:���!�ܮ�H'6޻�z���Up�$�&�|�Ub�>�&1M�M�4��6�ڮ���.�=4�q'� jW6�R�	�b���H�����9���H# =�%�f^�w ��ғ����c"��w��Y�T>}���	�%�U:��j�^�6��E�l_�U"�2[*Ụ�������'1qu_lc� <���YAd62�&�28ykyGu��Y������,��q�N�'�w���{������������E��ֳ�������x��*��7�M���x�3�\�v��q�m����oCF�?�+�-nfrϬ�jG(o��̹t3Վ�d0u�b��YzG�̼���}��!ߘ�Lp�K%rOlH%%�*���Ѕ�N�(/槝N�^����w�YFѕ2���ܨ�(^~h��1����ʤ<]##:�:R
�r��I��?Qc�[p���`pY H,e!Jo���?���\X���ll&%���n�3� G+��/iOR�D�5\a�r�1w6"	�iP6J�z#���qn�.*�@@l4�_���;��͊ �pH�A ���"��k�b�q���u�x��=��X�H���f�'�e��� �47�������Aw+T]|����u��E����Db��7����h�b�a L�M&�ƛ���hI`�bX0G�����nMN0\������,��A�l^d[Hf������5�0T�J��%82ڂ�����nw�b\:���f�������f��O�!�j�0y�,�8�PF��+{��{ת=���7�� �<���=����5��0�`��h��eþ����{_�r$��������v�>��]�=u�� �9}����L��ד�S�w�B2Q~_�\��v�Q��2��{c��t�@�r�a�P����|> �11�+`�B��<�����5>���!�9�"T^�`��$���i�+��ԇ�`V��Y��q �Uin͝�b`L�ӏ�L��J��bC��i�-����sU7���*8��/�X��Z�JQ��O�Ǣ<���6�@ ο�B�s��%_�$�.��Fl�=��S�F�`�y�}O��V6$w?�"��7:>rm|�e�o�&K��q�;X><0�P�2.|��`Ӂu�6��� l��|*hM�����@7:RRH��D�?���l}�QkWm/�;��ݞ��EA_�T�,G�_�#�x�r ��0�Gts�7
����6/Y+9�h]g����~�,�@/qų��H��S��)��`t���`K�)g��Ei�e�X	�}��Kx],�-��� ���4J�j�Zq�?����i.����1��@���7t�V�T��<�#��=�����P�Li�o�L�������P��$��^U6�z��S��4�F"��
��#��˺e*�m�?	��&W"���n.�k�
�VcP��y�юx���#��$B>!�@���<��􍥄ZU<�D�P�y���f	,�)?���G��\@ϸ��@��C���m\Ew2��|����<nw�g
m���Y;�f�I�fC���I]��"`6~<|�� ��FZ.\��Zl�=r��2����b@T��o��+s&�?�~h�e�j]�/�`��R���p��F#O��0�g�����o!t>��|w_���{V@Uj�2�����4|��2�'J�tˌj�����[0���zh�ac@��	B����t��05_�	�*��_�mxݗ��hG�p�4kT�~[���.L5a�K�}�M��
�=o"�Q�d�<5W��3����`@�(����u:�����i��x��J��a(���nP"L��S�d�&����,�Rl��	1`��9H�Ul�佋���b�4��<���/=�� �Z�K.mp�����z����BAz�PS���V�(f�]~(<�Û�T��3ƾ�y1t9\�S��{~f�V-�Um�j��[*�wئ,���C�sW�2�N��6ѝȹQ�ʬ4V}-���[#(�s�"z>n� ^�=s���������{�~z|4�#F��O��}L�X�C�󨒫Q�±��ѕ���X��E
����'�Ɲ^�T�U�U��2# ��n~���k�y؇/*Kj)E��y�v������6Q�����$b��i�lܭ�j��H��÷_V�sE���;��=Ex�S'z{�-{�������}V�����R�#ײe�0N�T^�2���(�?f�&�����c-�D��Bc�SZp�
�5BՏБRk����x�ycP�R�6(.� ~�F*'.��� O���ޗ�K�hW�x&�td�ۀ�I��>;]%q�����^n) ��2ӵ�t�zgI��C�/ޒ�*�P�.8(^x*|���腌y!f�3��A֞���`5ll����/ ���̠=<f{�r�":�II�He�R�B{�:h
>/�L�£?�"�/�jٍ�(��� J�D�ϵ�ȟQ?�`�1uޕ�v��8�Y�M�` xu��	|��l��w��V�!9L=1~��M�ʲ�rⰌ $�΋S�����&B��� �cC�~0��쩍vw�)e�B8Ѿx��DNm0��鼃�,/�G��
]n����D�Bs�JU�ޖ�ە=�Zբ2F
�+f��\׳����~kt��؛M���)���eI*�����q]��T�&�@z�*
<[oX��w�Ԇ5�J��,]��z��ѵDI��h|��mz�����SA�:u��|%i�2���M	����� �a�˖=$yt������7f���r������3+���^hIŜ"��e�6v�����_�FPRT�a�RJJ7j9�Z� @2�MO{�0ʄ�����`M�ab�\�t�����d>����/������g�6��Lt��g̶��NJ�{��#G,�*�ԫB��`���w��BS�V���5%`љU8�-C:��"��JI�L�i��^�����ph�]G�?7V��%�LA����&�]�Yj�u����c��kg�!\��Owf+~Xz
q�8�=��Uf�������a���p�����z�73�H�E����,�0��$盢|pr0�9l�1a��M�����(�)��	��4��'0��R�tRY��v�c�sꚐh�߬O9�k<H��� �^�0 d;��ϰ����������XT�ڨֽ�=	`"�%~���	��ٶ�ʴ�u����#�-��*�':�N���L\¢�_u��&N� �c�T�L6�L$��'k����>����d�J^�,J��IVY�f(Y�_Xu�&m���<�g���a׹�j�ȿӝ����EKX��_�M�^�_���^pv��Du���%Ca���q+nA�~�C������az�u���I�dK��bQ�^z"�l�+󂯊a����y�u~�����p�k�rʏo% �6�!��� ��Nԑ��&N���6��w�fF��$���H�C�^y�X��4A�;�^<x!:��R��ƔI��c�Bc�Z�����p��HGF�J���!ę�g?�Qc& yǾ�����{����O��Dܽ\���؞6��i�j<�5���R��S�*�*�lo,z_DÔ;�N$�[5�Hf�� �r/"y��=�[qOǀ�:��s7疘Xe����'� ��`�4r��]g����A���]7������V���D�D;7-�x�)�b�p� �7N�h�O�Ab��h��I�CIX˿V��d�noX�0d��]���=���Pȳd�+g�|V�/f5A2#�.�n ���]��y?����r:a��!D3�"��y���j!)ݾ0��3��FN���{��w�%0i��=t�5��<��s�8=e�7��S��{�Қ����@� �d�������ЋIh��ԫ���]��w���ie4���l�5Z���L�S��௽�~:�z�#9]@�>��J��v�M�lE�t��Hrx!�+�p�V���ț,���Ȩ��j�W9��5��\_��S$^w8�#���\�1+�7?�]VV�*��1���n������t~L-2Jp��b줤�� ��sP|��%Հw� X�NZQ��dH-�x͸�a6�P����.�0�Y#_��.x"l�ĩ:�F�;ky����ܕ$�|6"p��:b�|�Pgo1y&K|���jX�70�xU2�=~�����q��T��=�*h\����e7��#�7D���j��xN�Qc&#m����F�w�PgTX��GJ��#��r{~�0��c��
	�G��YfP!h�e0���~ >�@ꭼ�t'm��p�+7�t3v��[��)���E$���sś҇��&j�,�Z�k����KRJ2Ҁ�$�Z���pWe�tN�1$@�@qM3�2�&V/�5�xl�>���,G۶�5)�@��LUF�G��)ӳf[%��е�����9Hg,����i��/��"���_�/g|����m��	���򢶖ά.F����T�ck����G�S�)�^D�$�)Ц;OٗA���ńu�]����T�ܡx`�ĕD�{q������P�@�p��X�ER���~�z�&nry�e�ȿٓ;��đ^f����Y����~7�[����\��Z��rw�@�kЧ�ײ���҆]����>h�RPj�\�� 5��=���8F��ދ�P����ݠ�o��r>�۳|��ԦV;v��F��[;t4���2N�J�jČ�j�>�[+�]aah�8@ާ8B`O��OD��k�E��'��Ǘ���x�>��!!�G|h ̀T�E쬗\�.G�a}}��43�
OE�"�H�d3KW���3��<M�@f������8��3iQ��xE%|��y���P�N�n3�d�J�Y�,&;����[�W9��'U'c���	⎗���<��/�����Z#��(������;�mg�A?xJP�~�QR�f0�=(�gv��o�S�ƙ��l}�\����v�:-����� ���|�R�Rg�&1���nf�2=-��^��Bj�'I,}w�5{�(��Ħ��>w�� "�s n'�KU��|ܹ��4��������ؐ��~�:�=�&�~�������ߑ5l��
�
	q��=���O����U��A�2sx X�k~��q�P��BKK�Ƃ�K��v��Iz�����0��ݔڵl�5Vj~����	�ĺ�Ϸ�s��n	����9�x���zQ�-V��8�s��VͶb���t��#�SRtN���m��é\f��k�.V��?�D�+aB�NZK�T�p�^�k�
k� `�IIx�P@�R7�Z	���F�<���.���{������f�(Wc�<&�j�d�hO���v>6%�q��%�����3�FP2��Ct.�3g�BC��^�Pil)(8S�*�e5��-�y\	���=���˞��y`�41���,/{{����<A���Xzc�I���eJsE�]���<
-�L�{@?e%*��j44([�= e�2�P���q�QzŃ`�}�ސښvQ�08:���h���<��������l>�W����!k�=�rk�:پ�-�#⋋�$¨���h��*yBS�� U�~ؙ��ڎFčQ!")�n]8lK�d�N�O*������������4��Dw:�5p�9�K�+������6H�f����/�~.��y!�zYE�V4z����f��e$ըΜ�U?���&G���o[�{;�����ĺ�u��d�u�p�e�G5�|�z5tp��T��u�]���-u����`^���F��=�$a��|�E��f��f���y�G�-3'꽏*Rr^C���HT_� 7�v���&��(.T1�R��gj[}Y��1^{���r�r�=`h�7b.Z�⨡�A���>�o>����\�L���]�r�gj�6~��t�@��Q��NE,��ֽ�Û�,�*]hBB��ɄI.}wa �S�/�.�`���8���:lf�����5�?��̂Ү�5]p#�}�x�?���~(L|¤��<&��KY�l�u�(�C��N[B��\?<jO͆+y�Wze�.8������ſ�}a�g*pHk\��s���H�uR�-2v�3��$"1�|���4<�1�˂M_f��;%ڤHV��Y4=?
'�/'MLR��r�`X�~՞�1�\.9+�HY��\�^99I �� �Y�
�^K��d6TtX=ָb	�ry%9ힴ$�a�T�ʏ�6Cώ���=�(��*�p�	���
�zu����ۼ rU=�O�q6�������k�y�ǹ�t��2�ԅ5,�?ŮD�������U��A���B�=�P�q�Tw�%Qj�Z�Ch>�`�E�-�xM�f��L����v�6��2�:��C|lП!�n^�C;�^�
��T���C�6�df��b̗/z��\�f�s�%�ǋ�s�������!�pݫ�rEӂ%�D��\�лwN���]�ͨ�EQ	�w�V�F�1��	��(3^t���%��'�<�/G:�ͶR��ʔ�����vlc�y�?�&p�s�HbG�Je�s���ęҖV��y&cg�$ ��v���-�O	o�:6\�E��gZ�6Soi�.�����)�d�*�4l�qF_߯�;������H!� �4"�~o�Y4qP���%�o�n���)�X ���L'����t��4�z{��)%�DA-��]�	��"�;��^��Dت7��
�b5q {C�����H�Ci�Iִ�XfX���nʃP0Ҩڣ���o���Y(�D�d�/��w�\��5�S��I�e���8�G��+�����:��b���=� f6���|�v��!dow0�dJ�.� F��o�&�{� �נBs�����p;^<2`�3����z!���5�x����K�籞���%K���F����٨�4�=]�����f Oe��ژ����M%9S��2�8��~)	�^���<��������'��t�֪r�_����̑d濲���'��FG��ι�r�-�|�g5��/ї3!�X�,^FL�~a�=u+����*&V��ДTl�t(nñ���IyLH�%J�db�7�ߡ�����sK�pr�2/>X'o>Z���?�=mr���6����u�\��t��_�o�.Sh-lRd�DB"F�6�yg@�s�9$��N"뺳:�qe|5\�o��Kw�'��X�P�0���2$�l呶ҁ� �"2"�t��h�[��70_��M~DX�ќ>Cs�$Q��m�\f������`�T�+G妗#���rք�0>���K
��6���Y���h��#��~{o@�
��4hn�2ް�ify.t��7�V��)Y�EߟԎ�����|�,����>���J�Yk�6`�uj���dH�O*1_�b@���-�yV����v��YQ�租E�k���{�;L���B���?!�,�q��>�[gi��.��*��"L�4�i+U�J�4�[�Lm�۾	%v��C���`�.������1c�lE�o �.7̙�$x5��6�����j�����Ƃ:�/�/�\��i�__�v�7�3�A$�'����7E-�
��S��nm�5��!�z�;�Q�?�+f�<������X�~2�ױi��ͼ��\�Zb�rR�~�Zѧ��Ƀʥ���g,��Ch`�jSE������*ȦoF���י�|�N���o�]>�F�|��P�A��V6����ޥ��4���2�� J}�M��;w��3[&������hg/o@�u�B����*ɑ���?��͞Z���x��|�<��G�D��T#-Q�2+�.B=Pao�,}x��O��
�l�"�_�dnUW"8�3�_��Y�@!8�k�͵�pi�φx��E�����L<�P�qzÉ��߁J��,aC�+	�Vڟ9�-pU�m��5��	�����<�/s��^*Z~F[��M��W@�ťH*:Az�vP�n.�L�f��}(�+��ު'��)�tl~���\,���q&����-T�)��FI�Q���-����X��i�X2mKP�d���S�ʢ}N}�:�p�Q(:n��>��0 Ԇ�s;j�����gvl���45']���{�3��ξ��U�Z��w8�xŁ�G 4�,2���*
d c�~�L��!�J\U����m� �I!~�3�!����K������vb|x�J�F����+O�ڬ	�Ok6l��j�K���$���iP���2�i��b�e�XU�xZ�z�G�-1P��sy�س��V�r��w%��/��#��ΓNe�����^��f�c������p�Dה�BY�Z&�n��P��ok�r��i�sx:�xP.��R������D�|ݼ.�8��֧c�iNR��$qW�׌&p�d2�1�>1q@�ōkgt�]���;2���til!g$C�u��x/�P$�^(Shr*r9ݞ�1y��g�MhF���=*{`�Z���r/�~���fZ<|�0����u��I�Ce��x�>�0��
�J.L/Uq? q%��j���(�^ �ns:�Z�a:�Q��+`&�ދ��v�D�8��ૃM�!�֝LP��l�c�����!��{=����U��ʨ�@�f��$����o�ȟGB��  ��ش>��	�j�,�)�s�8������N#��GC�|�=V���&��o��DRc�@G��KQᄤ:�(GR�����������t����u��p���:�e��	�#�,���v0&��y蠁'[���m�{������RS��pd_�k� ��7|'z�eZ�du�԰͉ǲ���(F����@�6������=���>/���f��k�(�E{3B���^n�������Ivԏ��J��żT �R@�$j����ڔ�S6{�#��:��-|`�[�b�w��u��|P���h3>�/*ַ~��lt�7�g�W�6Y]�t�,���N@Z)�1�)�~4V,�*��B�𢄄�zw�E�S�(E�yF�`G�A8�C�:�j���X�¾h�ڟe�F��NyFp�N��3N?-���iL��2�Eǿ&�[2Y �RuHb��6x���\z��O�SM+t��z���8i�k5��`�Ś{azp�\���V��eHXŒ�Hy�}����}�$]�|���/,�1��MA��*m���=��/4x��'f�HPR�5��~����I��,]9f��H�7��^�~� ����������9�M�
;�T��ֳc�	�%�h�?���C��j�~��&�o�#`*f>G�Ķ���	��u�q���1 �O�J��6C�_�c��k�B��4�����S��,S,��?������q͌\�`����\䋆u��`���^������{i���D�M���)Z��-�v�Y�����C������*n��m�~S����g
�+k,տ�d�t�bG��z�������V���Q��+�"�@j�p�'r�6�%����1X�VmCN��:渖ͨ��lTwTFb���DGy�y��^od�B������<�e�:��R���ه�B�c縍���)p�]�H}hJ�#<�Ш���A���c&mc�i�1E��H�O��չ�\����-6(gia3!���>� ���	*f^�l��&_z��;�n��T8H܁� 
�"����-=q�ڀ�	�i�N�cX�)\�-n�'W{�O@�4�������J�A���]�?��>)궭�9�jD1<7c\��zb��� 6o<����7O�?sIF�X ��܋n%�A0�_��Zv���8���5��zd,S�rd���65���dU�����II��T�$��'�:/����,�;���o�Q�Qt^!�!$0J^��)��F�WG~�{P�u	�]!��J<�g�.���!�\P���@�~����t�ԋ�Ln��[@��0�Ө��m����]�em�4:����hX�ԟ�S�l��~���Նv⛖�ܑ�,����,�t�rn�8�����Ma�M`�"=Y�<�e�sݬ��傂�BY5ϪV��'#��*m^	5���/]���|+��S{V�Ĕ���&[n�k�s����Lcg�Jf�7b�Er��4�V8�sFf}��7���XB�ZG����x�+�Tڀ6��%��:��@�^_�D..�hl�>��iRF�Qy�.H!$�V/"fۣ:ϡY|p�og~�Krnt��E�Xo�Y0�(�2��F�l���&�C��/�	�Ԧύ�h~�T�2l�7����TD��x����n&�Q��m`���48�m�ґ�T�w#G�zg#��Mr1��0���ĵ�
�r��b�Y���h.�n���~��%@`�W�O|c)�ދ^.�ۃti�9�Q��)x��E��ԩ�Y�}��ܭJ,4��1��{aJ� v�ɿ��T��f�ו*�1�s@�,��(m�V�k�J���t&��"|�F%���y�L:
|�=�v߭+܌��&1������������8�%�N"��	�$_ϸe�����"m��V	`%(���4�.�&��;�c����y��	����l�$a֦1/�Mw�%R��xx��9�
�r��E���ѫq%��m܆���B(��N�GEo�-s��nh�V�i�5y;֨x���f����Li��E�~-��ľ��w�	\8&Z�rr-�촕��3g���p��<��p��h'�6j�݁�������A]}F���A-C�7�"�Go��4>�Ѹ|(�\��P-V1Q�C'I��2e4͕�2��JX�f�-�t�q[!+���h"Fk@dBV�T�滑��/��ȕY�p��xAb�W��GrAd�x�T^4���.=��a��}3Rj�x
E�"��d�SW���3��ӂ�6@��	E�摋͐��i��$x{����	#����PS�
äG6Z_��dS�,�k��8�Q��9Y��U���������2;<?7/(W�L3Z���J����}t:�#^A��P$t��G�.f�=(mh��?�I��O����\�E��l��� '-B�������Ϧ�#��/�g4��d�2�y3�g^,�
���Ҽ}�,��(�Wo���>-� ��sV��At9�BM�/Yw4�؜�����y��� �p���b~�S��삕���NF��J
����9S����B�Ua�S�S� �ю~��|�ظ@YK�`V�A�v=2��?��ߎ�qJ�5�m�
l-�cjtb��_��0 E�0��d��-;��*x,�zu^-63ɮ��Ny�V�NR�Ҁְ�F #(-�I��N@����:]���>f𻖙�BC��¢D��BԇmZ�X���k����ċ~x���PIJR-��kq�����;.�uB�1�ˈ$�����AWYi&KnqdI�(��>,�q�Å�&Z5���<K2d�t�DCg�C�H���aP�G�(n�*���y��yү���j��J����`f&����/q���]��<��9�CA�p�IZ��e�z���۬���
ψKLjN6?�$� �pj�Gq(��# �d����<#Q�`�tbކ�:v#�8�/ʫ�.��%��x�-��ltZ�T�!!��=b�Y�pQv�#+��A�I$8� $m���4�B	ֽ �B����ڄ[���)��8�ħ��*N~�j��+�߸;쮛�X���D��o�k��������U�J��w(���q�)$�S~�o�?0�"��� ��U�\��eڊ�D	�:��7x&����[mc[�!���|a��"v�0'��f��k�i��}�|Bc�z+wp�?����)j�Mp��#�	�^J"��A��Q�׊<LL=�ܪ�y���{n�f�����u���Ѭ3]� ��^��*��
�6��v�|��w7�T7/R��mj�R`��W��ZD{���ʕ`����`�U�b$���b������t��>���aH�'/�ig`��64��tTG̇��N;�{���ŝ9�s,4��*S�3B]3섿J�w��JS�A���~d`~8��x:�킴8��gF�up��*�����p�E�ٽ?�2pw�[L�JW��{&�
UY{i�u�/9E���+\��#OH�k+of�z=8$�%Pj`��uj�aKܽp~n^��鵆H��H5׻c�������$���|A�+�*<1rʲM�;�E�OښS�� 64��s'��C�WRj39NL��/M��l�p�9��VH����P^�� ��� ɨ�O��#��E1NT��N֮Ԟ	qsN%��Z�y�J�7�E]i������M�*������!��w3usbw��Z �\��E�o6����?�k�+ǯ��oJ���Cv,y�:l�w�����όw���d���=l�ƨm׊���?� (������(��#�WM~�)�d�[��|�v��jUK�аa C����,n�%������\��Κ칆�T�z��d�	Kb��5z�Z-��\R�[s��O�چV���ҭp��r;�m%�
���2��gNŌ��M�Jw��-w���F=M\��o�
�^j�ؑ�ͭlf<ɻ:��RvK��eƇ4.hc�e���pEgH���J[�P���6�HU�"&�����h�����c mO�O�X�\Ml���)6�i���f��7�Z�*A�l \_�[;�.Њl�H�,� %�"��#��"vqƟ1�[�J�dx(���qX�_'�H[�'���*�,4#�R�.���:A��c]h ��:�1��	pDN��7���,kb�ѵ ����rk��uS��4�IL�tX�����ȟn�:�0H6��5�2έ{���dǖ��m��?5r�(��,�jT���o�h����:r�w�R���VN/��Ē�,k�!���0�wH�$ �F_~?��{*��ז�+�8É���K<h� �)%��H�q�_���X���	��6g������]��>�м���C��*o�]g]`�o-c6䭆��FB���6SS'��.@i~�Nv�����>��U�ɇ�Чt!�r�<3��Wp��@P��Oꗭ$�.D�����rw5��-�<�����^D(�4k���H+,�/��3Vf����.��aHn�EΡ�l����L~CEJ�^wb����U�ɗ��sA�6|�����X]ݵZ�4���&�������6�@�+���_�f9_v:�.	��l�~��z�:F��
y'1��-M$���"�`:��|���o1eKmt��
6X*�0��2��G���a8ېXM'���*~)h9���M�7&��y�D�[��;/zi�9QtGmJ!�O�/�����gT	��Gno#�TTr���0�����
z����^�YV�h�!��~12@$��j�4����f��]�ts��L�)�q�EU������Ʀ���,o�s<����CSJCȠF|C�^������C1ը�@B̑�# UV@^/Ҕ��睰~�!�9���L���8[�:�w�Uh�AX�������ݥp�djZ� ڞ"'_�߲͸�h��Q$mp�~	��L��ʖ�(�.W�����c��$�e��h��1M$��-�,�\٨����t���r�0�>��Y�R��ϕY��l��ȥٸ�
��]�Ӓ���E�m�hM��K*nc�v~����Z;���5Ajf�p��52���/~(У����2�E\St�ZX��rO����n��^��[җ�2�+hB�UjIΊ^���>���ܿcFgeޜ�L��Z.�o2�>�|�|c���w�V,�뉞�3��ޣ4�2��%J3�V>��[w��nc�h�|@/r�B�c����^��2�u�tì��˞dx�#r�r��G�]�]$�T�[��h(�.8��a%-}�X��v
��"f�d�EEWX�3���M�s@��w$�aD��k�Di*�xs��~�Y��P�ÿw�\N�? �,׳h�a��L@d9�R�UX���)`!�������<z��/���ZZ4�Y��� X7������A�2+P��v�B}�fA}((���^���%�*��Y�\b�G�gN�K$-��v���5�G�}��{w��0��_S2#���"x9�%֢ʘFw}�"5��(p�Ȧ8j>��� J��sq¢ϼ3���j�]4k�T���c���D�G���,��lP�.Y��*�b�����
h���2&~�@��U<�$��� )y�~�I��߰�s�FK�]짼;ov�;���<|����!���1���clH��j�"�����k���ˌ9�_Ib�~����)xG�z�W-�;������a�V�J��-����-1#C�+�v�NX����Df��?髵O4 D�BOTZ�7�!��<�Dk�vպ]ix��Pd�.R��{�rˡ��0��3.��ƌ�3��=���W�|�&& �d��3��:�>'=iq��e��l�M��x2?i�t�<�g��C;I�.�UP��(��*h��T�y���g�yԞ��`!O��4<�/���8�7<�޶���k��I�t�e{.8��#�&�
���L�g�?6eQ/ujE (�/� �zm0}��,;Q+җ`\ wށ��vb!�8k�w��/LJ��S��h�Slq�>o!|,=�̋=nʞ���H�$s������XBd*[ �"J������\��޳)Q�&8=��}�gN�m���Y�Fui�3A��vp\��*tDH�3�
�)�J�5ǬܤpNW��ʺ�%^�H���O�j<�y�؇VZ�'�߲�QIe��HoR&h����&X�y�y#[ۤg�ccS��ؤ�k����6�f���!2y�x��|]�Nz����B�&����s����U��c��l/:����=��ٴ���df�+����	�x~�3xV珛H�^�dל��M��c=vʉc� ̩�2o�TR^R6�Bj��׬�G���{ڳ���7B���`�o�b�QsoH��M���>�U��mc&��|l"�gۈ�6�bt��A�"��N6���������,O��*��B8�����w21�S�z�/�y`�h>8�E:��z�]¨�81��a��.��`�pT��ɟU?#� RI�L-0�{^n&�ٳY�u�5~T�)nl��Sz\�y>O���+j 2zvW8ߐ�kp���Pya���p����N�����H���~g�sz��ѥ$Ӱ�|�$Z�%l1���M�VQ�`1a�	�u�l4��v'��'>�Rō|	��ό���[�K,�9��H*���Nq^Ji� P>��;Y��[r��ݢ��G�TE��֩e�	�#y%j���u���P�� ���Ҭ�\:���*���:$��<XX�uNs�: 8 C�@�H6������k 5��*���J��6{m,�;W�5^���-��K���}\�}�u�Ӥk��Y�%Tl����{���t�l��?����MY����cq�v|Io�Ғ�k�fC�j����n�����B/�ن�특᯽�5�jd���b=Akz����?�����m���30��[�p.,r�]E%l���Ќ��N�u��n�M�!x�JQw�qF����ܯ�w^e���A��'��<�1�:zRQ���5�g��9:cݖx�P{pp �	H�
vJ��������䔨�}&�o�5\������~l2Ozw�@\��̴8��6	2�i|�!"�oV���*�l[$_�5y;�����]HR�� @;�"�N թ7�qP���XL�_#a��XQ�6�ch�'��&���4^L<��1 ��A>�W]#�M�U�ꬄZ�s�D��7�W��mXbF2K �&;��U��-����JKI�ȫX7�	ֻ��n��0-�P�����Έ<a<ydb���h�mH5-yĚ��F��q��V�7���Kd:�������q���e�?��!�Y0��{��{F��'���{EN��:ڦ��!�`<���$]��
�?����O�t�Ӳ������7�m��@�\i��w@N��P��w�]Bu���@	�^���k��"�~o�SBh�����~�U����ٖ�������X��t<(rdۯ�����B����X��a�򐃨�Z�������5����HpC�)��^�r���,9�Hj�+G���Ih	VAz�n�\��n�?�)?��zG#L�?qJ\�"b���� S��;�s<�
�I�c�Xx�=Z=�o��D��ڸ�� 6{РΆ9��T�_�Oa.�Vpl���F��yxቕ�3�$��H"\|�:�a2|�=�o��Kh�l�8��X�05Y�2�+��"���������\���)h�
��hrK7���?�D	݃���9d~�Q�S�m����jx�cM�S�TDpLG���#�ۖr�WW0o ��g�
�ͽ}zDYR��hd��XK~���@������Y�+�Ȧ t�\��G��)..�EP��8�s���q9,�O��M���+�J���O��ƈ��\M���1a0@݋!���V�p��/Ջ�0P�iM�����,�[Lp?�3���$R>��\	���¥S�t����s�#�"]�4��&P��S���r�mK�6	֡^���<�.�-
��c׎п��َ�1��J�$I��'���{������ڳ��⸚��܍u{�00��gY��#��<(�x`f�D�E���G���Dn^�ђ�ȫ��;�-����f�:8�p7��)*~#��zK���\n�HZ�o�r��Y���iv^��f$��F�����h]G=j��_9�0�y�?�wB"F
=���7�����IA�o���>]G~|����'V':������G�f4� 2(�J�I��o��j6[����N<h��O@J��BLU�����W"�v���&��x�����Gh��8��TԢx�W�.3�+a�R}}�����
;��"Add�+W�s3{f߂�>�@R�b?���F��i=��x�w3�y,�]��Pə����_PzR�͆,���gG��9�U��D%d�zyr�{�<���/D����Z���,o�;��s���2�A+��PZ��=vtf��=(�6j�/��?�@�v>X�\����b��g�-����x��B�Ҿ��S8��K8�Z�82~6:�ݱ
�@G���}}tF!8�(Ez�	�L>�, u�s���7����ܥ�84����ȑ�D��M�������	ӻ��߯��瀻�
�
unȯ��MX���oU�%��� �@�~�d2��.�wK�zJ�7��v󋕴����!��]���V݀�lc�jj΂\5�Ħ���f*��Z���s�e��h�xbӔzk�-�a��$��؄j�V�f�9�`4�#^Ɂ?�N�(ڌY��/�f�i����Ե
�aD(�B�@�Z����\�͏ת]k�(
�zN4xk�GPP{R#_u��2뿰MZ�.�Ow�眛����ҡzWO��&�jd��R�P��>"��qQ2f���#��|2ƙ2�tU#gPcCzN���&�PU��(�g�*��/�yH�ۈ�;�W:�N��`ܗ-�O��/gI`�N<-��y�fG�I=�e6<��Q��6U
�d6L�|?�����j�/(G�� Ѱ&�vv��TQf\`����|�v�?h8&���P���\�.h���l��G�H�!�gT=؅�̦I��*!��ƀ$�QZ�R󹾛B��� A"��Ĕ�z𦍽Z)�C�8ؽ��x$AN4�x_�aW\߮fޮQE�� �"D�X��!5��J���n��,��89�r�����h���]�e9�n��B��B9Q�R�e��������|�&����Ѥg[�G1��iQ�|�cĦ)c$��ah��|}�3P�|x_+z!� ���z�aBGǃ�����I�L������2e�=k5�����k�f����9�O�3K�3���0i^�;t�4]��l]kvŶP�[�<����Tm��R��j�6_�G���$�{ի��K/�^�L`ԩb��N�5�-I���w�>�'�ȅD���N8GgVQ!6�0t���̽�^N1���B3����,j�8*I��Bτ5�+w��}S��/��O`x�8)�:
&��8�s���qf�R��_�p���?�e�-"OLh��ڙ&��NY1��uyϐoǏ�`�ט\+y-O~��+e��z�z8��E��6���+�ua��!p��@������=H�tl������w��$�-|w� � ��1(IcMK���{�ڐ���P
�4) �'7C9��R  ķ���	���&\�9Hŏ��4n^�o �ʓVy��E��ʸ���}6T��@֤�	'�#%%����)��@���H�/������%b*wЋ�����WC��	Z�u)�uL� ��מ;^6T�Y��k^�ǥDŖ%�R�q�8,Qz��0p��-Y������v��rҢ�+[�<M:���X���o� P�/�٘�M��gM4.��A�����vw�zH�&g�C�Tӟ5n����/\��;��`�<�f���-dғ�b��lziJ>�RC����~��L�<1ǘq7pI�Qr1!	%GP�H|C�'�N�~#�ɯͨ�T���|w}�F��Q����Jki^`��S����b�<��p:�sR,=��p���jeDc�5Ȳ���p�ڼH΋�JQ�]�a�虾���Xt&K���Ābc���_O�Rf�x\�n!�Ӡ�6g7irP��܁4�OP8�*��Sl��@_K�.;���"� H�� [}"yԈՄlxq< }��0�Z�U�_NX+��~��'uh.���4�'z�dt����A�K�]��,�p&��'�����Dă�74
��Ab��` g� ��XQ��"�����I¹vX��2ֶ n6q�0�C�kĻ��t+�cwu�d�}��c����5��ĵ��C.ڤ�0�]�%&���G:(����QЌ����3Y��T!P��0'��F�xE�{`�]׌���f��\��<�U�����ar�ĵ�mS��J��0��7����.��c���
�2�1.n� ��]�6��sl�V��ҿ�|��9��S]؋�$�~����J0�G�l��x�=�b�x�tW��rߙ}�r/k�}�J�y�i��M�����^��Wr�h�65`��у�a��]^�����ZǸd,+b퍇ļBV^�@������n�Y\�����5�FL�[J�}:be�ĤˊЗ'�s7����d��]X��MZ���)s�)�ϸ%Ф6v������հ�o��_l��.�;<l>_Mİ�3F�b!yӻ"�_Yq$��"��<:`�|!�no8�Kcಚ���X�S�0P!�2�^�����Df������ྩh�F[ۃ%�7��j%9DD~�q�_Z�Q*�m��l�����ޮ�c��ToGQ�'#��rBު0*R���
p��X�YY���h�>a��~�t�@��x�ԯ��R�<t:f�B�u)�
E�~���`s��+i�m�,�cr��3J��V�A�������ڍ��>1K9�@xki�� V��k{�Y��ed�A��|��g�L�!�.w��e0G4�w1��r��Sb$������3"���U�V��^h�G��m&	�X�Q��p�.��l��c򄤿[F,���̅g$䣄�"̒�^Y��V����=�&�~��%��Ȅ���&:�b#v�~���S���,a��j E�����a3����nY"�,�A�fX�;'nT�+V�fe$餫\���K�~p��|�ͨ:*\��VZNU�r�XX�Fݧ�U����M�9����hx��j? ���%���F3_�R��hC�d��o	C>82�|�$9ԭ�V"��Th����4_E2~�zJ�����E�[oP�$ZChSJ8@e�{B�fs��H���~U��Y��:�����xrx��MG��܈T
.���)..�a۳�}dR[���
�J�"��dZ
W�^�3vS���@�QZ�W	#�!=YixxxL�]�tњ��Y/P�<�����˷���>,M������B&9j�U�i�_
o����V�T<�a/߷h��vZ�6���V����#��ujAfO�P�D��8�f��}(�z��J׵���g��cI���\�W+�]���-@NT�ú=��ҙ� ��8���U��2��]���[��ʎ��}O��\��(�냦�>>�& �Y}s���ϲ���q���W4��,��<�ƒ����}��ᘪ�l��3�Vߘd��F
�}��j�G�h�~�6��U�W�Y�0 _((~�߶�4���q�K�p���~v�{?�6���!��e�F���;�!l~�Dj�9f�7�g��۷� �U5��~��D�x}�z�a-����_�����V�����R[�[?#y�����N�Ќ��\��K7f�p�������wgDCy;BEM4Z�O����{�r��k�����_�x&UP�$0R�c�P�O�mC��É.��K�B��U����`�WʡF&���d�
���Á>�3q����W�PFT��f2��wtU��g�@�Cu��丼P��(���*^@A�
U>y� ��R��U|��_A`� ��j�/����q�<h[�"�a�Ik%�e�����'��
`L��?lF�7�j�!�(L �&���͝�Q�z�`��H�wu�v~�8������;�	\�ވlE���rY!2�\=����u�ʔ����e$��
�Q9�ZB3� �A�� �����}��R)��8s�/�s�N���3
�|Y��)�ٮ,:��[+D~��� ��� 5g=�D��ɢ�s�ME'��������`��A�����9�]����ek9��Q\#j�w:8&�y��/[�Y�[�W����ڐ���\T2���Q��&�|�0z�k���8cԜ�C�ۘ�b��o�����A׊�!9=F`2�*�u�Lf���Yu��7�3�>���7u^�2�o/��wv������Ũ>�T��R,Y�j[�����K����{���ʦF�Ǫ`�>b�-x)�R�h1��Egr>��H�#Ȣ�XxuS��g�9"6�|Nt���X;�N,R����ڝj�%,���*�)	B�h�p��wh�S�Lv���$`3�K8D��:��o�>9��#X�F�A������,p�I?����?/�QL�'���u�&��%Y�Եu4�g��=du~�{�\f��O��+`��z,)}8U����e}����a��ApOcf��x��Y�HDD����:i���R�$I��|��,�1���M�Yܖu|�Ԕ�+�i4d@'�U43�R{������/�|3���99ROfH`B�:G^ �h ����qr��R��������XT{��֟��	��N%��"���Z���7���mju���+)��E*������r�F{�u���� y�ʞ6r�6���OTk6��� �� ��ԬI�,���+������$/�����s*����:�w��[ǽ���m1����J��%㚔��Mj�������Kvr�LfA��`C_8��b;nc���j��eۦ������tOի*5d툿b3R:zD򾼍��,�ȋ�	�ڗN��,�pd̅r��%"����*z��N����$�ͨ{����w���F�椄0l���Ks^[tV�����A2<~_:���R�0��RǇ��c��S���pvD4H�,�J�uV�<8���b8���)&������Xu�d�Op�A��\�Hj�n��6��i�D셗lO=�˒�*�Elѫq_�.|;�.��}H�� v�G"�y��_�Aqwq�,(x�U���]X��!˙�.'�X��24�"�����b�A��`]�p�^U�ۊ�� D���7��u�O'b�R� "^J�
|��#�Y���cI���Xm3tֱL�n�<H0yzɣ����wF�>M��zd�!�^ e#�5����yt_���s5�b�4����:��(��0�Ч�1�[�ޅ��!�*`0��J��$Fp�3r{{̊�ۦ�h0�-�<9:�-H�Y�"�'u�'��j�m�b�^�r5������~���٨L�S���G]�� �Q�o����WJ&��@iSxhf���*~\�b���K���ހhɘ�M��{�tr�rZxW�M̸݀2������꨷!�_X���g��(�5;N�Ѿ84�_Y�^�05�E���}D+}>��?1�V�a��{L��5n��-�����pNLϗJR=�b@A��B�¾Ys2���G	���ݯX���Z3�����dٸ��6qP��<�P��k����_��W.�@8ly���KHDF~�Fy.����i$4��"R�]:;�K|\t9o�=K^F՚�cX[$P0k	�2�����<���Y�)f~��Ԧ;�hj�e۞��7�/�E+PD?ߜ�ZV�Q�*mL����p��Y09>��T��EG��#�I�r���0��0�k
�X�3?Y�{h���\6~BF<@L�>���O�C������btՏ��=6�)�E�1��6�i���H�h, 
�W���[�JT��wT���<��R�͕��S1�1�@ki�y VQ�i6K"��@�:O������L���)5�K��o0��q#��O�[���p,�5���x"�_�n�щI��o�mqW	L�<�F����J.h���'�c������u#���=$O���ٹWZ�r�������v�����f=�]����������Ē:��Et*�����(fnT״���!8G;BE��cf@.���y�_8�~�h�0�[�c��\�ZZ�Z!r����l⧟��ܜҨ{�\�Vh��dj�_n�_���ȭ�'F I�ޭ©�#�[Q�o~��>=|��HGVܣ��h����x49�q2��7J��l�2��{[[ª��h��@�\�BB���q�h���t�F]������A�x-)!��WG^s}��TJ���9�.)G�a65�}�{���
1�"���d���W)8=3q`ۂ^w,@�EuA!������i��fx���o���1�P?����)F_���&,�L��27�=�9���U�U�zB�p��1R�<+D!/z��D�ZE����$�q���i�I���NA�!P��'�3ȪfR(>(Y�|�e���5"�ƻq��T�\3H��X�c\N�-�<��'�ź�5�tF�������P`P24sA�S���v�d�	do}*�0��E(A����%>�� {^&s�6��-2����0�B�4<�L�|rb��ʅuM6���L��&3�n��3��J�
+���%�������X�U�w�񔔾 �/v~���莻ؤ�K'_�-�8v��9�q��M�Ď���������l�`j`���u�����ň�P���)/����@x��za�o-xDɚ߼غ�=V����>.�֡<#��5�YN�*v��+��e��fܗ��P�f��I1D^�?B�y�Zm#��$��ȗk�쇺0�jx�bFP�MR�i+Gz��O���M�.���Ɲ5l��l�@�WEdS&���d5Xͼ���>u�q!Ǎe�+�(��2�?t���g��%Cp�В?k�P�~g(ڱ�*٘A��Iy�|x�Tms��=#`R�Ӆ�j/]p��Ʉ�<��支W�\��I�-se�	���G���
;�aLVs?�V�*jVUm(��� }�ɺ���Q�� `-��r�Kvs�8��
�1}wg��o;3l�t�X!�ZE=N��������(�$x$$f��3��ȕBu�3 ��:�;��p�s��)n�878�n��N���
��{:ߤ��O���D����V��[?`�M_��.��yz�(��U�� ��[Y��^ظ���x	�H�eFv�0b���Ўr{p&iC��G\|[,�ܷ��q�2����RZ��W`��2t.��|��\z����������ǹ>e�9��cp�����(��=!���es�����f~����:{��D\3�⹏_�^eI~��!����/v�p���b�c֫T��R��
j6������Z-2{��n�~3���,`
~b�V���9���v�>��&�~*A�&�n�gLB�6���t@����-N' ^��-��%�,�;*?}(B�~r��<w��S�帢@��`�S�8_+�: C���Y��L����4��\��6p�����?���3L�[�L1�&�9Y��.u�b��3ߩ6d?F\�ׇO��W+[�Iz�b`8_������	��ea7EVp����=��Q�H�3�ϼ-�y��-�P$�P�|��v���1�G�M�fܱG�چ���t04���'m��/��R�\�:�<� d������9��H�p��_�^[�� ��������;�&�����1J�T�֚��	���%��/��/�6��ʱ������-���
}E*-'��k���������u�e��D ���1�<6
y�
F_kQǛ=����b���K,�W�&����z�|������Тd�
�q����������Y���6��e���M��r�P|��4Zvm�%�(М�C�E���n>ٌ���� �!���ι�x�f��d�vb�
�z���ȩ ����ڇ?����Pp̡r'U%�����$�]�N��U�`N�6���wsMyF���kE30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ�I�7���~��v ��UWP�Gh1�&�f�
lX��%�`�����h��-r��^���Gr�K ��:�GU7G��YrJ��G�~�-�u��	ʂ:C���'�L�C��̏������:�������w�+X<2=a뙹":4���2�9��&�Z(����ƯOW��aZ8����Z3:�t��7�;�Z#<���Bj�ӣK z*s NNH_8��*��;�=���N=��N�L����AV�܉H���mq����9��Z�~���5L-�I���C��������W�p��⢞dv�ߴ��SO�t�t������v�tFAo�΀��ɨ!��zJ�NFš1mf��9�mYF�V�7v��E���"�>o��Ds�;�i��(�VVd�;$LKh�z�Z�O��]Q�w����(�����9w�_A�}��2��b��4.e��QB�3���
bC���}\�B��FO3��N��W�b(ؕ=
jo�Hg؄�A�\d��х#VW��\[$��"�9��n�1�p�~��dvo�	F�S�bJ��'k0�]���1u*v�tq�2f�od���߈p�����H��-�W�x������]Re8g��vt&6`�6=��
�=�0	Y��r�$�SF�)�%�i�з�m������^@�$r�0��V�A��<#�Y4�c���T���ıąF�Pn~
�sr0Z�G�NVq�l^t,�PAAy�<����6l�k�V؁>�"� �m��C���A$�z٤e)/$��A�{&U.�R {%xE�1u�������z`X�[R���b��ۿ�����Ǻ8NH��z�����zό���+Z���ڸ��1��/�V�+�(z X�����b�����y���fUW4Eh5.�	���w����涪as�']�C�w{�hM|��.���>�@9S_m10�T�)Ȍ�{朂 ����4�g�4��U����+��qҭN�� y颖�S&AòMnU${c�<�'Q��&���/�#����a�G3�s�����\�F<*��]T��/���4"Gg��Q��^V	N\���B<D���}��^�F�W���,*�	���N� �X�ZP.��UN��+�{��ب,m��'���[�ӑ��Z�gi�hg��5����1���z���6~��p+^y��Ik�[JJ��kU/�.r�����ׯ�����/ls8	O�jI�>�y�|�Oe���CLS�1ŷ�ܖ�.�j	bx�H	YO�m�R-�e��i!�.V�6�5[��5��ߑ� ֡c8��⪊pkBXlr+a�� ��0\�COH�3x��{��k���H��e��|�agE.�)��ix#���
��1i����t�P���vEAM}
mRj��h>��ᠷ����7b����U��~,3�*M{ى��$���qśڰ���J*�����,=Y�������o�ٴ݆Hvj�;���њ >R,���|JW��{ߝ��+b��k�</�	�ܷ����4g������<x3X�ܚ%����Cƭ��d�����9r��5��@^:x��bO����jr�g�ာ~wq��������:�i⟺�'Lj�������L�ǔ�פÌ˜0٘\
��a�m"�}p����9�&�<�Ȩ��=OdEai����|3'�߲sES;%�<����Ӱ� '�Wm��HL�,���;��:��p���"L����{V�H�-Pm�@N�'��9�@��w!�B�X����1$i���S�K�C���pd�Ϣ���킴?ĦS� ��aZo�c� ���A��A�Z �ʊ��U
�����;gT���َ�I�m&\�V/V��Iɬ 4Is��� 0��>VS��z�V�P�;1��h��"����Ӹ�Q,0��Ϭ�(ǣ�Cڴlx�}>�}��;�!&��ZG�BY���O�
�iF� }	��B<(�O V�N��W���b6
�a%o����Wϻ�0d��	���LW��\(�'��6���ܿ1������dc>�	�g���N��n���sJP1��v�֞���M��3��	ϾF�ۣ!�Jб�l�Q1sˁ���A�֐e�]s	�EA�#�8&�|X��='a��j�N	&�r"��SSz���;T��Է��D�(�@ѐ}r"[�c���:v#�o��P�R�L{��\��~9����P{Z�� ЂZ1���ʶqW��^��_=3��&�ͮ�}吙G��=��kU`�h?ys�Rwt�j&:y����8�#Wl,�2�o!eCts"'(�sh%�N����"My�;����P�5�c.�4!qq���j����MGs����+iy'������ڽ�<?|���_�i�ú4p9@UY�O'��s,E��yFJ�{� .9��лZ4���K���"ǥ�2 �Q���e��=�>F�$�D�RE�l�*S��hʎ�98sR�7��:���nT�	t��)R��s�`�9-��,�EF6�>5���9���6OzmW}ق�Bp7#$�-��Kz� u��f߆�B��Z�S�B�J0�2T��8�����c���@���ұ�{���I:; �Wi�{�*�M1�y��A�pO.� $��<ʩW�n�i������;��t���C��Do���p�Gے�2J[U'�vPQ��]�#C5����*A�U�,Tn,8t�^�K�P?>�u,cm���AY�S�����4�y����ł8���e�zx�x�䔪d�\�����1[������%C� ��!��I��s��cј7����+a�ǩ�z��u�Su��G^�������w�9u�f�s��"NHM�Mx̬��c^�2CC�ip�l�[J}���Y���fQ[0?۽��i?�n��U��,U���q�ݸ
�J0�]��b������ʅl�PJ LaWe�PVv�_|�]��`)�we��$p%c�ڧ=ln�ȍT�_	O`d8�b��Zz��;9�����l��x�g��F��݌D��c�{'��9��~g	'�\Ίz�������g�I�cuw�4H,�5#+ 0�e�$�ј�es�$���.3{.��� �*TE��Ѳ���V��zS�[�&��ir����\���Z�����YH���zˌ��=�%�U�+m��MD���*}�b�M̾H�X�9��ÛbqU�/y}�f��E���.�Y��gꁡr�����8sb9�:�{0��|"f1.����/�@�TB_����Y1)��d{Z. L���'j����ZU���!ά�m	r�!���>�y|���F?����Uל�Ŕ�'�S&&��f/�����4⦽�G��J���j�o�=<���]'��/,ш4�S������ܿ	���a�<��A�ly�9'm��⇖JdZ�J�	��N��>ہ��Z#@n��j�� ���{��@�ߚ�:�F��X������8/h��5���o�]������}��\���m������J��+֎$����OT����sl�� !���J�[��>71\pE���\�\���ӒQ�ed��N���7�(�	�q�e�2_x�^��I6Ŀ6[q~(q��e��_��q-�ƶ� �CC�y_K��$L���!���d��]��/e��XFM��R}K�(S�������\Ȇ3%�zf֤�X��s}J����zI�K�}����%��I�n�������Vi�����ZgZ�ĥ��c�V��U5-�c��Y ��#Q��d��bz�����)WAv���:���}��#f�z� ���2�A��p��I*����L~|�Ťf���KE�cxJS������-׆a�j����8�d���Đ���I��X�<����ԕR?{���[�Ϩ��$ˍ�4[R�)�_���^L.�gH�b=T�`���,K-��Ft+���|�g(O�l8�<��ޔ�>��AY�Md�t��G�=8��,?����/i�]A�3C����⨒�;6
rܭ��x�\��L����	�w(��?��:�������m�+,�w�)�'6K�"(�y�M3Ѻ�<�v�V�t�c��g�섑��������`dYϴ\P1J�t��Su�`��3���:|��x`dϱ����!%~z`/@�V#j�E���.����n_��M��f6X��A������E��{_z�������$�bf�6̩�V@�Huq#g�t�L+�1��Y� ��0����q��]����&h�zs���?�""`M��8o�x,�w��]�nl"ٜ�/Y^K����mܿ�W���;|H�r�� ј��:�Tv�OI����rMMnW�~��7��X��4:&Q����L`W\��]�8ֵ�����̃�����ZtPpua���"=6��m#9P��&���~%�y��O���a�1��λ3�������;n<e��%����sE �#�rH�٢��n;����N������L:�|���V��H(8�m4���9?�e�a��x�u�\����>������gp�h����ǣ�5��SR`��א7�2������iAR�j� ;<�K����G����N���䋔m�ܛV���2ЩɢM�^�<e�6�ţ4.X��QfV9�[;g"�h���]g�I1!Qb�O��r(}Э�}.���d}4%о�(ݰ���Ր�\B]��U�
EC	��:}���B�rO��zN�!PWˀ*���
MQo�ׯ{�p�D`d������W�"H\��D�<�� ��1y�+򁧯d��		G���N�ժ�x�@�m;�'1��Mv�� L�ׂ2>���b�n���v�W<LЧ��wMA~ҹF�*7���G�]�P"{B��� &9 w�N=]��`4	ܔ�r�V�S�������l�]�%�z�V�/@�mr��י���0=#��2���_킈b����4l�)�P�ƙ�^Z��8�p~q�j:^��M=�	�&LmW��sM�=a'���k��N���s�23t��&�.
�aH8�W"v耨`�!�ҁs���)����h��U0Mo4�;@��}o���W*-qҦ��[�ֻ��M
^]W|�-���R'�n�e�u�3�U?����UG��y�4��SU���'���,�-�y�Ƹ�_�$|�]�4x��ف���谥��C��ؑ�N�3��F��Ӻ�R{a�� ����1�s�s�2#��O�����x�_���i(`�r!-��{�I�4:P���_�
�F�`zc�=�8�pB��[#Z�޵���z���<��3S.�����8�BO�E�:��T뺚��g�u�;�V�����1����� "gi�B *��0���zA�[�.
������q�W�:i�����a;Fa����C���D%���Tt��N�@N�'��P�e��{C+e*Ȗgo�ˀ"T�n�ji�^��aP���ub�?� A9v�2��j��8�{�1�S�'�7U��p"�xr͡���3�ݼ�7Y[n
�u~�%��E�`&�׿�I3��ܚю�̒K1e��6��i	�k��uD�^�R��6��m��+���黩"�W�C�����^*t�CyV�p�KP��ϸ~șY85۫\Sm0����ټ<���bT�� �T�4��{�J& u�U��FJD���Յbd�J�M�W�*�V�Z�_rְ��֬w��m$f^�Ð�il���Tq�_�%d�Ͽ���RK�9��S�U��l.���Z1�<�"�B���٫f'��D9�y ~)�ϊ��@��(��J��pϫ���*C9��|� �@��L�M�r/��/e�N�$E�a�$�v.��W d�wE�Zj���{�mz���[�F��_���`"�Ҕ���j�㛀H?u�zA�V�sy!�K�+#lf��
� LU�XG*�t�kj��X����$b�"����Zy�ϱf~�E�Pe.�叝���h����Gs�7
�L�{&~|�XI.�*��@��_6!��=n�)ђ{do CT͝ɢ���qU�/��ׁЈ�3�W��޲y2��⼴��;�jU�G�{�L':��&���/���M��I�G��3��'s�%�M<�]]�-/"�4k���-�z�C�B	�ZnʺB<-e���g��/�(������v���A	�~�NR���}OZY��b-�▔�P{*2Y�՝E��,o�D�*��v����h��\5�����q��D��y56��[(43,��x�ȖJ ��+����-�bǏ�y���(��̚�Jhky�t5�\f
L��+C���~�	�_�[���ќ��`]�(�ݬq��22����Il�&6QW������~_>Pfq#�[���C�IV��N�K�OLե������'�SA/@DX�i��)��K�:#��炝�\���%�Nf�`+X2��}�l��"�I�T����Lr%�������X������ה������#���\ě�cz�(�-&���-��*1Q���:'�������'S�p������}���fg�&�6K�()G����:�*�_��B~Դ{�lf�,K{(�x@^A������wa��/��_T8]��`���K���l���|��<Y�R5��Eb�7�x��T���k1Rj?W_S^��%g	��>QOx�5�+,A�m��H�t�������g�$l�籹��tc�AO�._ts��D��,���"�bT/���A�,��iY��B��,������9����D��������(��c�Bw���}�[
1m+|,�՝��.6�(A�Mi�����,_I��jKc%���?�D�1�7�*Ɩ��Ϫ\�P�N ��U�=]�V+3�jܰ�����7ϧ�UԤt!�/�`e�v�L
,jİ��j@��ɪwnU*3MiI6Μ��w�i��y����{�V��{����m6B���̡Hk��g:�G���1��}��>^�z�f�����]ն��c���1k���"�Ɂ��q���˭ >]��-"���/�2.a�7��7�%_5���O�v���s��ÕD0b$e�7�<�p������Ŗ�����ީ%D�\�T��6�ڵw������� �ٯV���$.�b'Ǡ�Nҏ�y���������c�$WS��a���(�8tp���=&/������z�67�����̊�<%�H�BR��m3��,ōT��IC����f���=jm �#Rq`���˴d�ed�������H�
^��a|���.+0��y�:�:i�謩�1Q��_>�#"�h���?gx�=y�o"�p�hK��F��e�S�F�Tut�9z��\�V�7�`����S�c���9å-��dHYz-���nx`�}g���O�Q2n���
�h-Ֆ�s�i�Mhj�sF-/;����;�\3�����6�Kkv�5Q�5Dޱ�h75Y�J���wa��f�cB�կ��I:ǅ�W$n�z�Ϡ-=��X&S�ѳ�2����1]�K�n�_TSm�؀s쵟IO�ȸ^�i���Z`�@��_��@�u�����*/�Ȟ�3�z\�Z4�%-g"�"�W���� Zg5�:fH�o��2��̒"�����
4�%��[T|N�� �~o-�zt�A��� ���I�P
��3|�r�!�$�{�H�B����79�XIy��������|1#K�*$�����b���y� c�90@2�(|#\�)���[u���4�6�
��>Mm0_<Uם���!<7`��D=kOA��U����ό�Ό9��a��X����h��n}�Qt�;�ҕ�V&-����U��;)��h����xr�����$����v��U>w�K�A�˱�'l�gv��i�yv!��k&�HC�>s#�#��P��o.夘7�95��M�d
���S6e��֦߄���x���*wmȉ��K�N/��v�e#��*��7T)[6A(6?�V������W���L��M��L=�Fm�u-?�D���ߎS�7?;mLy��6�Lg�=�Sv��-g��O!���qY���M�^�L�A�j墣��%��n<��fAN�>��kY��H[� �갡a���~�x��}E�	����E��� =֞%��q�@}w���ZWR;@���`Ճ�}����Ԙ�e:)�T�&(̴Zj�ƿ�ϗl,�W g˴\q���䧩����}��r`88C��z�sB�<��nI�YH�
F��+%����!o��`�	��<�YS1h_��B�[7��\E�\U�S� I��?��hvY�	&�g[ ��~��Ff^l��5��vT8�h��%��V��yNFY��E\��An5�a���3�}��v5>�A��'A�����Osb���v3=R���R,�av�U������-���Id�����0������v�#K�����n4�.OB��/L:�G�����v�[O&���2�ͽ�н�qZ�4��t�H�i��0Ԫ���@`��6��+�C����b#����yy*��~�c�+��b��oJ�n�HWw�����*�5�9�<���Y��,�><�w,;|��������-�Q��r����C�)�D�������Da<?���QD6��[8#`�	��\�+Z�,����y����S��8��8uW����g+�y��[o}-�<C����F�I[8���]5���<�})<1���~�sq�����������V�r���Zn`�A�p����2�<�RC7�!�Z�0�:K�����1��=p�Sl�B��z|�s�$���B�~���]���F��ꥹ�����O_��n
�s���h�7F��b+ /�X�9cw>@��&AW듔��* ���Kz�K�9m��B�Ke��څ��1��2Ɗ�������a��m�l�2�`�?ɗ8>We�Gz6�ȥbS�w.�_zZI"�:�ɨ
T:�5ugL�GoP�L[��� M�ؙ�/!������T�b�y��� �;��K�����!?vRf&���N&�r��m�<}�������0P���N�a��\Y�4�̩�nj����h*SMԝ~�,�Հ�~�)Z?�-�����c��Mbs��C���#�ܚ�Sk�0����[�V0��7bS�X��ahtw�:̣��C�ݣd�8��Q�A�@@�"��M��J�H�#�a��wNƗ5-�d^�)w��.�d�2��݉[nËڟzc�ߐd�7�K�����s(,¶G�p;�v��Oc'2l���O}t���=v��~ ��pI�)�z�Y)�\a��e��O򫒧D=,��zWp����$�2v�ʞ�/{���<:�{>V>$ID�EP*�r� ��i���j����w�;�s$˹�2Pj��|z�D�?~��Dܗ��۾6;�����Bz"���G̻�L~N�c!������Af�زTry�G����P5��;����.�ی��2�ب����T�j�ɵh2���ӷ��N)�j&��wO�v��nt� !_�2Z���bjDr�|� `��x�0�l6J{���;DѺӑ{BY5\5��L}17Fy3��w
�}/��zvW�g��eVbK�W�@��4(!�(7si�G��C7�U��t\M@َ,���ҡ�ʊ�{
,qC.#��_�jKM�{�HT���L�'��������?c��&��j?�4�RU�'�]�,lw�yM��bɨ���w��4�]Nٲk�i&��\�XQ��L��ziF����.zR��5�q��܏Î��Ns9�$��ˆ����Ro��bۺ��`_{-�h��,Qе�������e�wu�z�J�٩u�B QI#�{���!z�8K�Msx�d���0i%�B�B����:T��`�k꜆�<U׏�s픢N��PI� �G�irh"*��w� ��A�M.[��'%��C�XW�Uii����>;+�ź��CK$�D�
�w�#�y���4'��IP�EQ��]�C|����#�\]TUs;R�^���P�=�u�SF�]��A�L*��J����2�l��d���hy?���x����ku������[_�Q��a%)o��f˟�H��I�d����L�_.��<Wk����0���u�?�^�\#�mM��>r�3�� \"�V����a�^��(C*�@p�y������$Yi�«�J0f����G���z��Б��IԸe���ŠJw���R��ѧ�i��3#J��}W�V�D�_��<cg5�wL?�$7O#Á
l��:����_Pd_�ֱ�}z�@9��F"l?�P0�e����ݳ���j6V'�`%9���~ڒ:B���]�N@��d�n�$�J�����ܪ� �, �} O���4�e#��$� ����.�4 u>JEj�� ԝ}(�zZ^i[����0�y�Q���������4R'H��z�"��$� �E�+���ԅ��Q�gǩ�����V�3�Xćס���b��{��!y��Vf�$�E"�.�؏N/�9���p�?s��}�{w�|I|.�|��kf@��_'���N`�)�{` sGo�.\�n�_U{�,��Vʈ��@���M�Y�y�mQ�MHU��U�l� 'K��&f�/Ok�����ݺGm��q$����<$�]��/s��4�Eā�'����	Ș�ʫ�<>[�� /΀G٭ x�Q�O�fYN	_�DNC���CZ�j8������%�{ۻW��]���6�U���p/��Ih!@b5�jp�V��pE<�jP���Ԣe���c�u�9£J�/�+��@�{Q|�����"à���.�g��=��J���%"�\7������?C�:����7R�B������(��qu��2p���cI�A�6���O�0�l�#_�~�q�ә����C��(�n�KU{LFU��(u��Kwk$��/@'X�g��Z��K� �?x֝��k\�MV%�)�f}��XChg}��L�<��I@Ʒ�������e%�XE�����i���Y�(�Q�+ߕ��;}N�l�ck�5Q-W4��U6�^�Q�G㐥�ْ	ښИ#�)±����3��}�f�cz��?�����8�1���)*�D׳�	���_f�-~K,><x*���@E��{�a/O;�4��8Ώ��v�w������I�E�m��R��S��@�v���P����R[G�_!Y�^�Q1gZ�1��o���WR,{c˽�Ht�5��b�go6�l_aֹ��h�%��A �j)�t��|O5X}�;3����:/P<�Ao=.�ZH�z}�O��}���&��/�|�$�n����(�Z�sû�_��&Mm�&�,��2��Nc6��(R?�M���?�	�\��{qc�B���P�5�J�H�m��Q�����PX-!�{Or��'@3�L��o����[�����4�!,�`W��`�j����{N��z,n� �M��76_K�(}�TK��w�{����ֶ7���66�6@=n?H<\�g+�Ԑ��A1(���G��;ݴ����X�a]��s�T!����6��"i�,��.8�3�^�]Q/"�N/�D�.L�V7����|�m8Og{>��ԛ���DA�eL�?7�j<<v��d��v�1�q?���5D�p!�N�GևZ���:�R�pg����Vﾹ�5÷bX�%���@B��ǵ�mg�y+�o��
xϙL�����pSh=��8�pE����'�� ,�C�����0�R2nI3_��^4��:<��ꅖ@���ʲ EyRϷO��d���U/��0@��(���[����^���0G�0yh� :Z�<����Q=
>�g���h7g)�,yo�a�MK����c�S���T恻�5W�L6'��7pM�`�!�fS�h�g(z��[�d���-a�Qni֓`�:���u���Q�!�5f�ω-�:��d���^����&��!O�c�;������s�H�kg���5u_*5š���YV
�)�ᵀ��T�<��Gަ��f�UʰnA;��Q �ᤁ�&DD�$��2!����ED��R�nm!�S��DVß:��ɀ�i����J[@&��J�"���f���4�ȯ.��a�Z����B�"��D���ɺ�Z�p�gF��fyt�o�)���"I�ȇp��4����"�|_�h�1υo~,ktO���i� 8quIs��
��9|���!����u���l�37ꅳIJ�O��`?ę񚭦�#���$S�ր*��������vu �0Q5�Y<0#�>c�Tq�uE��4Z�e����>>i�0�Ui��n��!�����Xk =b�&T��	6xϝEν�^ײ�	X�VB���廓Ɯ"'^;�ߘ��^���7U��5Y�)M�hXD0���r����P� �$vm0�U��>�X��r�_\��XE������I�%�X��"u>�D#�n�P�for�Hߊ9>%�D��$�ݰ骜2�}e����o��F}�ԃ*�$��3��������7�e���*��7eY�6rZ�?����^
��O͓WQ�؄��>��LN�Am�H~?a�rD�(Ǒp`r��B4>ƒ����Lx����,�~a���e�D5k#���^�a��R�Aj������a ��X��S�<U{�9�[ ����Q8���mx�%E�ޢ{�t�:���J N��%R����+�)�Z�,;�y�1SȒn˟�
���2맥�'(=}%Z�� �ixl��a �m(�����j.�R'��8?8���K��B�6v��hYyqF Y%oX����oS{ʁ�\E�-U�SB!����[��\v��[6��^� ]i?��
h��;	Wa�[Q���f��@l30D5�\�vEU�huj��s����Y����7x����5�����q<Dѐ+� ǹ��O0��e'�Ԓ<~sS���3=�������a�r�YBB�ȳ`�ȉ�9������\���ivzq׫���?��.@�R���p:?��a�m�|�*v.��[ �"�gH��������q�����}Hn�5����[����p�'(��<�~�وKbtʂ�f�Q*z�e�,&��7b���o[M�n/��wX���I!z*����R<��*�~���dA�oavw}n|/3'�z��:��Q��c�҄އN)��S������E�?t]�Q����B.#q������+�i�,��.�q�9ð|p�$9F)2�8����/��+D�\����}��i<�Y��Fz�z8ܸ]f1�ʍ��)��f��fs"�o�����<���֣Ͽ�Y�`x����Xs�R�֤vC(0��k[k�%��fV��E��1^��p�ot���zm���5V���~$��]-@F����'��Z�3��|���94
(D1�d�/��86F%�(+ь:XRMRw���r!AD%X��D��>��Y8w���m�=-�<Tݠ�R��b2���c���ʜ�i>m�72x�?���>�u�G�Lc�C���_+��.��YyTK�zu���G�'EL�|♱<��J�u!� ���T�cI��@n�e|�ň��ܴU��!�f��_�rķB���o�/s�H"��a������M-�E�˩�T�����َ�Me�
uq��Q��o��k-ϼ�}Y����b��CsH-������3�ABw��^կ�`W0%�Kb���s�tH������&�Ԉ�N���	u	@{ʟ�@oJҠ_�42a��]N��-gM+� kwm�׉5���閇[�@�о�c'��d� �ܖ�a�n(��G�`pL�U��cxҁ�~���u
t]�=G��~^MpZ�$��߯z�qa ?'�gI�CӖ=Ҳ�j+�^�+���j�����/�s/,����{/��$Z�E�gp�Ψ)�i���y�����,ys$��c.ɶ8!����~�و��j���@e6,��ÂBM�P�0IF�,�~��<c�Aΐz�\�2�f�òy!h��i�P��!̈ܵvD��s��#F�ع����jS��&:;2;�x����Qvj�8w`;v�{��\ ��2��Tu�DCF:�����k뭝9al�H���:�-����Π1ӶM�R0�o)����D]1α�?��L�����G"t��^�!�i�7ˉ�5]�`"k٠/+-�.��=7�ȸ���Q��O�JL�7Û����D���e�f�7���<�����mȡ���Һ �D.�p���z֒7��S�w��M��,57�V�zd���bao몧1���n�a�y��ק��h� ���U�o���q���p�GA=n^0�� ��V:����k���e�J�$`]R���3�G���-�%
ܗ2u#������ ��fR��n�zGAd-]0@ױ�{�����'�f�Q�=m~�M;0ry�y�͔:E�6��?Q�)>��u�QV+gT}�y����L��K@kGʯ��S���TQ������8�E���7[&{`���t�S%}���~C��yd$E-��nTj�`�+�j��<�Q[�� %,��!�-g��OB���j�O�6����z��K}�̒@�kR'g�7"5 �q@�DШY!������@�ˢ?�NMXQ��t���҅��n˘�|���/07&/��o�2��ǻ�A��'��n8LpSI0r��_~�%.���i��'��!F@����%����A�*�����V~�Z�oC�6'"t��p�Tz�Z�!$g��nf$�o�,�\��"�u��s 4h��Ԏ|��t���o��t����d � c�MI�3�
��|��!����b�c�7�<7��IՊl��B����X��#���$n2^�K�O��=G�\�`�0�o����#�7Ҩ��u*	4�@��fw>)�Y0j]�U�ga�y�T!�Z�W�k+�X��5���Hv���h-׽2�X[畊�I~���?��c;ǭ���0	�J�B��ܠ$�)��h����+��r����+�W��9Ovx��U�>�\~�TR��N��C�ʃ��U���0ᾌ$d�>�_;#���PZ�\o
i���a9銡�)_�^���{�ܜ]7�eLIϿ�I>�d�*����Iq�p��u�e�g*oWU7�k�6�	?�������~W|8c���)$rL�όm�/?l�>D�U�;;��wv���ՓL�:�/<sމ蠽+�3�޹��Rp�^v��j���)C��J-��%��;��ģ�$2� ����=���
8	xl�(EW����͡��� �$�%�Ē����Zns�;>�ͼx<�Y�ß��Apu����(��5Z�}����l�,�������ձK��9�����δX8#�֫_B��]��k9Y$B_F�%�"9Z�3o~���e���]�S�&jҝ�$[���\�-&���j ��x?��hҳu	�4[\b���
����l^7�5gIBv0ӓhX�9�hh��K1Y���¡ ����5j@�����'���Z�Ύ��q��;�']���s>��H��=.������a��J��:�S����8:BƬ���=�������gvE�4�֡���S�.+*���:�'��lK����v�I�[+懈��J�����Mq6 
�~uHٞ^��Ԇ�����Ї���|b&���ʾ*EKn�@���mb~/o�E&n��dwc����9w*m牏2�<#�k���T�Gxť�|w�D|����E�ve]�QA0N��)��)]��^
���*�ޠ��?�2�Q�����#�
ܢ�6�+�1,^��<�"��Lx�H��8���ژ5+O+�7�}�_�<%�B�Fe48'8k]��ʘ�)*ڒX��sM[�<�ʸ��-�p�N���dC�`�ےh h�}�d�� �C���w�o�q���5�1)bp�+���5zX9���	���=~/�]�KFl���+��0����1��$-
ӘG�o��Dd4F�c�+�>qX�D_w��xJA�����	���$l �'ŃmW�Ү'�,�6t��X�2"�o��X��ۘV�=2m��2c�?%">3;PG��-ȁ��ӆ�_V��~����s�T��uC>�G�}�L7��|AT�uER!lq��ĜTH�`�U�s�p����/e��T��F!���f����ro�����&����]���\��z?�8x���\�s����[�DW�M0f�� ���:�Z�d��.-z��?���"b��WC��_����}�1�� -��G����0��b���Ǟm#t�GW����O��9�����-B�@�S@�J?����J��߼Fazs�N"	|-�sSb�w�	މ����Ԉ[���{ןc2�pda��s���E�(�VG�p�'Zhw�c���������pt�w=Ҏi~�ţp��G�V�?��a����2\��n?�=]�G�4dT�L��	����2��[�/W8rܘi{q�$��E,l��h����is�&�F�{�VjͲ�$'���"�C�>� 3�~n�C� ���UCh6i�Y�PB����;��̗�~�G�c��ِ ӯը���y����t�P:W������7,�����9��cj^�ɑ@2Z��饪dTjW�w�]�v����� ��2�
՗�nDδ��"�Ԩ�H �w���j���TW�bYt���	�>W1L0�����ct���G"�Y[�����+Y�"����3���4>�T�y������[����@��1᠇o3�򋸟���$D��X�AN�q�@��e_��ҧDv1���I� {_�;h~��l�"�b�=�$=o��-h[d֚�f�����s��KO���s|l�g�ټ�hP9*�#x�� ��}��ŗo���Z���~e4�N��I������p�Ul��9�AGڛ�U��Tf,N��3.r`P�x���M��I���(- �������uR�B�����R@͋�B:aIg��I���e��#u���:G!�G�p�F9V!O�C"�)s}g }�GQ��\���}���O�RTg����G���Y)�pQ���\��l2��G�9ͫC�`�BZ(�)���n~^���Tz�w��E���Tt���[M� ��<����%O�O_��AU�=�%U��������5(U����Eu�j DlK%��2>͢�am�!�߮��L��P�8h�oj���Ϙ� |��D��T��=1/��@��/S	�GH(ޑl;vR�F�$92i��qV)9o5�2�<�(�G� Uր~�c�t��I�Kk��l�l�~�k0[��O'h�xL�/�Y*k����x�����|�%=E- ���b�x�0�صg��k�#c�^�X����wS��$w�H*�l����*�_���d����Α��
��9��V�8l�f�K5�����۷Ƒ��'��9k�/~է��V�h���3: �ƕ~h�Q�p��L��OV ^j�����y�{��eJ�i$����W&.]�� 3[E��g���/z�N�[�{��e��e���.�H�BǛ�sH�S�z�I��+���&+��v�{�)��To�g��,�*"�EX˪m�q*�b��&ԭ�,yk�f6D-Ei�K.Ͳ��UiT� �7̦s�yF���{ަ�|��.�H��@��_�C�����)�C?{�+S ���U_��u�Ub��]���D���a��y�~0�t���-�U�c 31'�}q&�/}Jϰ����NGt�m�X{�ݺ�<�<�]3�/��4#���9����	����ry<�������0}�G"��x���m	FB�N
�ۯ!Zڸ�wB��V���L0�{����Ǩ����n�}wN�H�Hhh]5ѷ��]���Wx��1����]��kZ��n�ݥJس7+ċ6�b{3��D���ʎa0���b\��J �?�,B0\���OFJ��6i��d��tМ�S���(�"�q\�52̈́񤌕MI$��6	O�������_��)q�⎶L�cC?+�g�K��L���Oո�R���/�5Xt����N$K:��ІF��=�\�ɲ%�&�fD[/X�:F}8��I��X���L�5�%�L��?��]�������lـr[��@&U���S
�c2){�u�-މ���<j`1�Q��������y�l����!��(�1��>.}T�kf׾���������>l1*z�Գ��C�3�f��zK3-�x��Y�m�[��a�i���D8h��r�~�:���a�������1gR���H��[���Սmw�R"�_�, ^:�{g����\nne�,�/C˄tY�ՕjB�g��l�>~��9�,H	At�Qt+5�����L�gV�~�/W�1AV���!H��r�֜�]JwVΦ�P��)d�U���w_(�t���g�mކ�	[m�Q�,�bB���d6�7	(��[M!�Ⱥ�,����x+c�����+��k���K�N$#�b�]P�� ���c��Yٔ��3Gu��hD}�f..�_r�\!S��`,���6j|��"ڃ��{�n�M!(�6�R@�/ S�;}��{��<���N�=?��Ѓ�6�t�Dq�H#�|g򘊐zݳ1��7���`��k� ��_��]�*���G��sn��E5"�#��:r����B�e5�]8Y�"G��/��>.��7tr�����PHOn�J��Wi�y
D�$e��7Y�<�g��F~�}mr��Җ<�D�F���t���5��/�ʞa���w�@��V�Ҁ��Oab��B����k��O�t�u�`Y���Yq���r�ӎ��_�Op`ID=ʛ��w�|Ų>��q ��&:�\w�i)� ~�RYd�3fL��EPҊ����q�����Q ��R)F��Vhd��-�V�ר ͯ �­�û�L�0N��yO��:!ͣ�a�HQ�Q^>@����9�Mg0��yVܾ(�VK�f�ʋ{S@�T-+���cf��77B�`Y��h�HS�[�خ(���d�d �d-H��n0��`W_u�F��r�Q7Y!�\�"���-� ��+�A��:�+� �鈪\&�i�����$�k.� 7�	5�fF��> �Y}�������TE�E��_,�α�����&�nh  �X�,�L�&;���82��ƻ�+{��n�=5S%MՀ+E��]�pX�il�E��)@mWq���]7�MC���	*�V���2�fZ��ݣ-"�E��\ɕ�j Z�&g���f o%oHu��8{�"pY�w�~4ę!Ӱ��|����`�o��)t�(`��a+ ?nIZ\�
�D�|`L�!s5�3
���$_֓�7�_I1O~�]�@k�4f�#Sr$J�֧������}C<	)0�V ���3#fѨ���ul_�4a!���si>I�0���U�Vi��NZ!�����/k�4������D�D���D*4���X7��;���H�	�.;�mw�EH;孬מ�m�|r")t�6h_ˉ��]�r`k��N���|hv�3>Uɂz>/����ɱF�)��Y�z�O1���w� �b>+��#�#XP��"o�'��J�9�=��5	:C(�����9�Fe���������i&�[��*/�1�z������e��*K��73�6�h�?[�Z��ָ�v"�WX������	L�2m��??�5iD�K����W��S�%�ڪY�L*�'c��.���ɦ:�rKe�0:^R�x���Sj��@�%(�&35���O�#u�� �u W�	��L�f�xH��E����8��P*��| ��A%�Sy���i�p`Zʔ�;����a�5���C.>��y�U�(�S�Z";r�p��l䰷ء#�nՍ�6�a�:��T��*�8��2�WBe�Y�&�Y �Fg��%������oZ-��O�����S�i[�y{>[��\��n�zk��'� G�?��<h.��	�U[������L����l:�5�=XvShh�+��D�[�1�YרY���d���
5�І��FY�>H���.-Z��/��=��'�%�y�sO(�X=
�k���,�a.�`g��y���#���d&��X֍�v�Y�ײ���&��.�H�]:�~���}��ÓvU�_[KH�N������u'\qs��yLCH�8��u�bם�S���/@��q�`��bې8����*��������هbZs{o�n�y&w�����O*��[����<o���3:���V���9w亙|vt�ɡ)�A2�Q���*����)9��H��b4j���?{#lQ�	����#���5�+�,:�ޘ��÷Y��L�lY8-1]ٶ�+����4Z}��f<�M��3�FA�8��]����L)�D����s)�)q�ʔ�׉ �*���`��C�����Y�Ҥ�|�C��;��S����$�˷1�cwp��ٹ���z4]���z��}3�~�ɴ]a��F����w��A���{�'�W`�
�?͓�[K� 2�FL��+���X9��w�t�TP�A˷^�L(a�~們��^m�|�p������6.2~:���^��7Zz���mn8�2?��?�1�>6�G2L�]A��/�_2ǀ��_��#�T�uU
G'p�L҆��:'�Qj�!���⮐�T���1/���;�ω���U\�!��fޅ��h$rK='����v��o���h�����|Z�$��O��]�\� ��M�3H|y��8�)6l�-VpP�w�$�Ф.b+e�Czg����Y�ا�׻�c����0l�b�F�zt/��nY�Ae]�[j��,��	(��O�@�ԉ.-J�Kۼ�5paVNoN~?-�}���wt�o���ΰ�[&U��W�rc���d=M��hJ�(佡G�NOp�ND�c�I^����c�td��=.�~؍�p��2}���ag�9ʎmO�J|E=�| �p(���( 	e+������V	�/3�����h{�p�$�E��*��pmQi�AE�"Pc�z���-$�c���01��t���A~ʢS��X���6�B�õ�KBԒ:˗c�s��~ɵc�Fg�aH��(U�jn�y�����$�P���ܼ�y�������`��~�~j�� �m��2b#�܍��tj��	wev\�&L� �-�2`C�[��D*�e��ʕ�0L%�$/�ӊ�FB��r� 3��Y�`���-��F1�v�1{
�����U��G�Z7Y�0N���+�_g��*�3��4(b�y��˹N�NL���.@R#��|�&32�/�{4�N�D�~i?Nm��@0.�e;Q����1�S:���Z{;(�Ħ2�H�߾�A� ���W��h7&"�=d���H׬ύ�K+����g�i��k��F�9�>Mx��j�]�����U�!>�c��2�e�-�NQ��]�_�,~��9�$�;6)��&�0|�N]ym3
`�i{�s^��I�m��< z����f����u���_Jݨo��g�:�K5�ʗTY���[�|u�aH:#�LG�ǲF��O���~�ٵ
g��Y�Y��\�Ȝ}�A>Ov�1TCh�	�1�~�)[y���\��H���|k͇�P���C6��)OenZ����z�T%T��q���̛� c�y@��$'q��u�#E^ʈ�UU'�f��cْ�b�2�5Ӭ��Y!k.j|��K�ݎ�d�m��}�6�����
��8D�j����t�)|j�- %`�^�:�8��o��i]b	�0tH%p���JR���Āp�i��zV���5�|��5�~E��gl��\V�cSH��%'Hk2#l�ґt�����0�p'O\�x����uk��W���G� z|~�2E��Z��r�x><M�!�
�iWi�m��Q޳�ϰE�D�
(5�� d��Y��l����_��7]J�_����,N�xM����W\$ ��q`֛��v���w�G�(,Xim�`���C7������6���,T>�����oJ�L��V<�Ɔ�.�k�`2�d�D�]�M�OMہ.TM�Q#Xх%�2?�����w��˅��7r���@�:j�]	��+rR���<�~�.�}��B:K�����]L����ԋŔ�,M�B���~�����3�Ha� "B�@��7�9���&���ɧ�wO_`aab㸦���3BiI��e�; JO<��@�J;�ӫ� �]�(��HgM��2WU;��+�Ӧ�����L�p�$��V��cH̀my���|9ās��ใ=N�����]����ƿ����Zp������~4v���SW��|�n�OG���\�|�Aw�t�Ŝ}ɰ[��.��V{��9C���bma�2Vʰ`��&�}�{w��-{C��{�0��V^e�;,nbhZv�bp���{Q�]����/(����g��}�~ľ��\�<��տ�B��S���E
jT��>�}d��B�ЅO;N�>W��؝�V
r�Wo�G��IPd�S�+��W��q\cD��*�����1����d~ԟ	N���j��/I�e�A �}1�fv��.�тw�j�g�縔��LW�F9�0(�������ap����S]�@A��~��&>�۪=����E6�	a�r�e�SNz:�1;��q�T�󺶿'���EJ@a�r��2�^����>�#��_�k�2��K���;(Ĺ(N��Pv���{%uZ�1"��qҢ^|#�=ng�&q{@�xFX������}kpc��㥮s��Yt��&Ց})�8z�W'Cy�M�w!��ys����d]�� Є�JMԉb�@!��k�k��*��'qW#�ڀ�ͻ~��MoHL\��:EJ��'�������X�?wq����~r^4��U�Vh'x��,�ly�ʴ�v�����S4G��Ƈ������["���C�`���BF���_l�R����ܣH"�8ԖsM�i�W�f��ǹ�$�ȉ����N��`-x-5���@��������*K���zH�ٽb3B��u#T:�O�z�����ʆx����/9�6Bt&7��QTP�d���q��z�P�Տ������"��E �qkiկ*�Ҳ���8A+E.�;�;����{�W�SJi�A�����;�ڢ�tC��D�G5��	ۍ�8�
'�3�Plτ��'C�5����4�Ti�ϺJ^�q�PZ$u����~bA�1(�W��/2�:��3�����|���U��x�zr��P��͏�U�O[s�g%=�%���\"�IX�i�����&�PN|�V��� �P�uɠ�^3ಿ�C��*+0∣�Nk"��J�(�� �~^O�|C>Xpb���'G�#0Y}�P�A8�0z�M�sǼ�+�t1w��e���H�3M[J���/dkQ���҅��YJ�>�W�<�V�V_W� �%�%�w`��$�W�Õ% l�����,c_�6�dsps�;���!9Qj,�Z�lӳ/D��!���2�����'�N*9��~"���gŊ�5����p�̶�^��؏�c��AY K�W���T���H�Le���$
�F��.��< 	�E0�u��V����z�կ[����{<�eQĿw�����(�HĞ�zf�B�8���E�+(�@�h�0�e�X�=���m2�SFXؙ���/bջ7Ԛ�Zy���fc��E6��.:�Ïb>��8,愯�s}���jV{��|]�>.&D>�%�@-
�_;$a���[)k�{�D� �@���w���D�U�	�ܹQ��l���Z:��Ky�:<�ᷙ� �U2�&��'ߡ;&*�%/����/��A��G�&��'�*��<��h]��/��4𺮁R?L��I	\�_ʿ�d<�.�����U�����z7�	�NW��ۜ
�Z�2`㤬<�#�ږ��Y{�m��:R��m���R��
X�u%�h51"5>~.�jt����~���w��y>���3��M�}JE�+�ܟ��Ƃ
������?��c�Q@J��;�9P�\�}����w��N�V�@RX�V�Z��(���q	ɪ2G�y��I�-�66
9c%�� ��_Uq�l���Z�C,��.�K�lLZj���,�_!�s�/ �XaɊ�nR�Kg��Saݝ)�O\�˻%jjf��X��}�5����IT�P�7��!%]�������"QX���8�?pT�H�b5�� cܧ��y-kD���Hh-�iQ)Oh����&F���g���豵����'X}!��f����ٍD5L3֫+�b*�0�'�&� �f0�'K@�x�^�����H�"aCۅ�Ⱥl8�p���Pċ�܍?0R���������R���g\�7���9�F�Rof%_�Z�^ǅg�d �_5t��u�,�[3�ѤtFe��jtgA-ls�͹<�K�9�7A���tk=*+�ɶ�Od[·�/diAƴ�n�E�wȒc?MR��=��'��J�� ����(�DɇG������QmP"X,�@����6�(��MM�����$�	6�f�cℂ�G���I��������}CϏ_�Pl������u���3���U�����!όڅ�)�9!��0`*A�����j�����O�n:W�M��6��<ү���� �{z�G�/���jax���6g�UQ 	H�0�g?K�g-�1<73�ە�O�pՋ�L�lDV]:���h\���`S�Jз"��w����2{~�r>V]�I"�]r/t6�.`ـ7�+r�����	�O{�D�@ߛ�ƛ�D�:e`�7��<P���S�Ȋ������Dw
��b�?������������>E&VJ��ɰ�bl���3��5��*_����ݰ�W�)�����<�`J���p-�=7�������_:.;������WU���&'��́Rƭ�3s�����N$a�{�K�T8<�"i� Y��R��׷c��d6O?i
���}V�<�.��q,������0[��y���:n5��NZgQ'K>mLq{���g=��y���u@�K�u,��0Sm�&T�n�^��!�)��)7���`F[�� �S����{��R?Wd��-��*n}�`D����)��Q���ɝ���-p�+�x���g}��:��}�w=��}��s̛�k{��$&�5�Gcɯ���Y��l����I�U�h��O�[�7�.���i�in�n{�e���8�Q&X����?25K���$��7�n��S2&H���NB��]�)i�Zh�?1�@:�}ޣ���ĕ��9�35C�<0v�7�NsϺ[�������z����ܲ����"���� ����DY���!��tYe�2N$=X����.��$ \��E�y{��ܰFBz�,a[�!��WӞ�X�q��,k���F���H7��z9h{�k���C��+]FԻ&��[��P5��l<Kb�xX���}bȋ(��{ey�VfvR~E�u�.Qc���ա`9��w�s�79�D�{�l|��.�&�"c{@��_.z�5��)�	�{�x �W�͕}Y���\�wh�Q��d��1���LY���#+�A�e�V'�F4�4����:)ka��o"V$w�3&�9�Id&,����2(8Os�Ea�p"���h3֫L��W;��-<���ާ�ӿ A ?'<��H����F�>;=@B�礂�;h�LD���V���HakLm�4�ږ��9�S2��R�Q���$� G��wMN��Ѝ�rp���:�+����.ȝSk���75"�N���}AV�����D� ���:��a��M���]�"mu�V^���JFɛ;���u<���M���פD
�V���;@eUh�3ȇv|D��1�Q����><(��6{>�{��}-�о���������_B��$��1
�`;�ݯ}��B��O�L�N��WDE�رJ%
�o�u5tU��]�jdP
��?�%WIP\w�驾�����11rG�(3d��	br2���F�CY������1��#v���R䂋w�7�I�҃�u�)�05WР� 
�zt��`H�����u]���T����&R�����=�����	u��rQj�Sb\�Ŵ	���8��!��(��i�@ ��rAR��r��)Q#�e���C��� <�r����~Z�~pP�/��G�Z��̩�q�Ko^�=��r&|���YU�6,���k����"gs0�!t!_&i�k��8I�W;?h��LF!�Es�{L��J��}�#���Mh�B�T���ɥ�O��tDqk�H��:��0�M��pW:�kK��.'7ܨ�bh��9�?�ԟ�N�`����4c�U�#0'`,�v[yuo���2�pJ�4����(�Ƒji�0����t�t�,�aF����XR�A�ۙ��ܷR��� 1sa�M��ƿŻ�Z����\�`AV�-�D��T��-#`���l�5�*�zܤ����BH�#3����hz�+x�u�C��3�XkM.�Bo���+T�ug��̜�#�dZ��C��=��xM ��fi��*�6�(g$A?��.���O���kl�W�V�i������ ;S�� tCs?D�I+����ۡi�9�j'�9P >3��Z�C�/:�/�x���NT}R�c�>^�1 P��Qu����6A����v��C���P2��t��������Tx������!���h�[�Z���x%Qd���e3�pt�I�(m���ч�a�d��Nz�m���5u�ƌ^�����>}�f�PD�Y�"a^"�Y������4��^�CR'�p�7�*ḷ��Y���Փ�0�k���׼N-�7���t\����GZ�J�ɱ���`�5Q��R��["�J��rWK�V�Q_��W�9c]�A5wt��$_Vé��la��g_x��d��y��1w�+@�9�k�nEGlgj[X���ũ��PXƒ�8'�AS9���~6��br8�	��v%��Ɩ �rp��#�!�� �&����w)��\�7eK��$E��:.�O� ��9ED�i�(�m���z���[�_��X�"�y�t��վ�� �\$�H�`z���L[)�D�+<(���U��yr���8v��5#رX�b���b��u�.\^y?"f�F0EJ��.�id�v ��a�e是sɪ�y{�ڇ|q��.�p(�.@���_O�|�v(�)*�?{��] ���V�͌��U��3��a��2��Wm"t�y��"�u�R�x�U��f��='s��&>��/>e�����-G�a������>�><LP�]��#/��4�~��#�	����,<f���0�
ΨY"�(c�y�%���	��Nk���0�Z���8���7��M��{%����b�	:6�}�ӑ.P�	i�hI�5��I�~����{���K��56�3����a�aJ�c	+�;>��/1��O�J��	5��O�e�>J!�=�M��\_	��S����bN�ԑ�j)��}�(��xq��m2.c,�@�IŞd6ʝ�w+����_0dq���J�C����.s�KB��LnD��PI��s��L/4��X�!��kKK�R��gg��"\�Ni%�Oif���Xk�<}�"��d�Iha���W�%K[%�&��b����_�6��P��S����v`Ĕ��c��;��-��}��A�CQ������ٺ'l��{�%rT��۞[�}5��f ����\�!z$`�����*:!����x�f��KT�Lx9����s����aW��\��8�[�ğs}���'%L�:A���|R��۱�H���D��Eލ�w�R��_IA^�>�g�@u豭%���,:������tڟw��sg�pl����G�M�AH�r3��t���>��]:��cZ-�ͮ/x͐A��Ն�Ì/Z�wt��)1+�^Χ�a�����D��ثn(4MɛPl.�!���Um��,س5�U�6U(zo�M»Q�gZO�{����c��a���ƺ]Z��p�H��.��#3�P��B������d�O��3�4����I�J�� ��=�]!T1�`>0T�E^�j݃�ܣv��"��n��BM6�GI�P�z�|����{l��C��0����6��+e��Hd�XgS���[31P8��o��cD���ה��L]�Ÿ�|�ِ)�@�^�U"�wЁ>U��'�ˆ}@]y�{"���/�.t��75�B��:��	O�����TP����Die�eto�7�m<d� �G�Ȟ���_����D���v�֯�����b�����T�bV��]�Ib�����Y���[���0_��i�=r��2���tC�� )pA�h=�D��=����O[<�H<�k"S�*�}��/�RZRB3���ņ�_�bpP��$�h�.��,� m �R*�ݷw��dʼ�}*ӬX��P럃�w��a�J0o�y�zJ:�)����Q;Je>������D�gQ7y�����K@��,=SD�T!���5UfO"�7�@Q`�yO	GSB�T؏o��zd!YA-��Bn�q�`�������3V5Q�U�]:���9-���6���.������s
��Ea�n�Ѝ[�/n�k�w�@.5���]� Y~.����s��NĢ|�V*�R�o���D��}�/ni��yQ����Z&lN��LB�2I`����b���n���SF��ltʟb֎���?iDA��<�@N45r��GT��P��C�%��	��V%Z�W���!�"����ɕ�(0Z'�-gnO�f�(o	l �J"q���c4	���|��ԝYzo��twH���} `
�I�|�
�l�|��!���b��ە�֔w�7�Ir U�����)��;�#���$+�%֨����u�������0ym�сyP#� ��|��umΠ4�p0��>f�0G�U0NO:�!�a\��¾k(v��N���1Y��ť���2d�ڵ�X�ߊ<��l��J-2;����1y�ǧ�_/��]xJ)u�_h��ʱȣ�r�yW�)r�(��v��jU��6>05�8����	��`8���
�JӋM���t>,E2#�GsP�d�oG�d�p�9fR��F�<P����ZuPe�F5����&��X*𞎉[Q������`�e��*��C7�ш6��?�	��qP�w�Wy�� {@�f��Lv�Qm"n�?��D�7y��Tf���fdT�N�L��>�ަ�Ľ�զ;�N�D3N�^�l��z)�j>-��F�����Y��ڢ�dC��a�� �6顺n�'�Qx)��E������>У�4& vK%9��$#�Q��Z���;7F�Y�8��C��rl���p�ͽZ(eԺZ#�@��9Tl%��9�I��8U�.��"%Ŭz&b�+m8v��s^+BƉ���9�Y��;F(f{%��]��o{�����UP'Sj����=[��\��M�j9��_ B;?�w�h��
	nf[y�_��N���l[�5�vm��h5%3��(���k[Y��>���죹��5'K��d�l){S+V�񐳖1�>�'ɄԺ�s{>�%4:=��,B���a/�z���D��1����|�A��v�
��!$v�~~�ӯV�g!X.h�T��>�:g�-É��Ĥ��vV�[(���ܧ�R�����q����:��H��I�|Lԃ�Q�9e�Oc�dDi�.�b����|�*�4t�%�$V�b�w�o���nWtw����qX�*�ݝ��Q<��V�-	��$Uw��Vjw���|W�ɢ�Ub�{Q�~���C� �)�}�{_��C#:���T?�N�Q=�����#�ޢ#	+�Sk,+�ޙ�����L�pQ�8����W��+l�����}�D<�K�$�F�B8I�]���ʵ��)�i����bsJ~������o�
W4��5߁̬`��N��dQ�zZv�5�CP�w�;C�
�ߎ�?�mO41�c�p����;�1z��v�]��\j~L|]B�rF�R���P���|��G��i�
Py:���_�XaFMϷ+��Xz��w+?���JfAl8��c����;�$I.m��ͮdo����Ŋ��2?
M��&d�8��:B�m� ?2�s?�>���G��>Z��0Q_S�lMƫ��Ts��u��-G�L�;����M�r�!	P�YT%ܤ�ҽ8捞ŰD`�?}~'!8�Bf?ɓ��r�ܫ�����W��p(��A#��Q�u��m�"��σ�E)�FJM�,Y����y]����-�1:�8�F��R�b,�OC�R��������iZi�|
��"00M�<b�ǛYotp� ������!��Me���:��w����@��A�F~TJ���\��a�B8N?�-��U�\�w�O�]���B�[������2cOycd �{f��8.(%p�G0I�pt�^�9c�4��%���t�Y=o.R~9Y�p��֕�D��=aH�Sʏ}��k�=���E�A���8�&x���H�W��/T2y�5�e{Wޏ$��aE���(SQ��i�3��C�g���-�Tl�$n�ɋ�S�`#���ce~������@6TR;�6�kBu�Y�X�o�T�v~�yc����� �Z	y��ZpyI�ˑ52P�Dq�`��w֥ԙ{�K1�����kj{�N�Ny�2c���R
�G�j?e|w�3�v�x+�p ���2�ۗ|�DDk���9���������.��'^:�sILTLKY�����}1�75�O���"b�V�|G�Y�}T���+66�a�k3Ү�4����z(��$��Jk�pJ@ӵn��M3��2�\C��O�VD�S���gN� n@��]e�D��[1ų1��R>{\]ҩD��? �ޡܚ���h�g�>1���L���K�US�P-�R4"�5��mH9�|Bx����BڂY�*��մ��G���
eʀ�NR���~'%�m��)����]�ms��K�� �N^��3+"`�N���*F0   �   ލp�F˸�$�B�H'�1�#l�����
�޴Y�:��O��d�����	;F��lx���RUO�=SLP,�ܴM~��ibӪ��I+N�V��v�/\���J����޴��:�)c"<�$�s�x�0�M��:�3%ءm�Fi�EU�D�"F�`���KE$4?LQ<>�6m�S}�hY�(`��y5�[16v�uꇮk2��b�i���ǎ���dQ>9/�����pC&C�<F�$�2���ȓzh���U�N(>�%C$�Ӊ9,�ц�k�P��D���7zV�
p�H��\��8zl�u*�;�`U
iS���ȓq�p�s2a�/Q����%M�Ɇ�A�>���(`�����-��8��I� ��j���x��@(H��.�h��Ҋ�
g��@��1lL��ȓ$�
�ÀmB5_5�x�FcX�d��ȓ
��12�H�����S�Ȣ����i��$Z�Hڕ`=&@aaD&lŇ�Iv}bgȔF�841�B�l�F<"�g�?�K��P�O�ꦹm�\�DAbI��������]?2�@9�*,s(~5�A3�I@�<�p�>	���U��z��,]U"d	�b}ba\�'\,�Ex��gk\���,S.v���(���yR� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��                                                          .    ލp�F˸��%�R(O5f��p"O��Q   ��p�>I2�P�?)����S�$�F�8u"�7��   �   ލp�F˸�@�r��9�1�#l����_�)��ToڬrN�'|W�DCĢ�M��d9����� �д
(Ţk^h����i�z7X��ߓ|!���GO�>�.t���'?C�h�獞Q�'�-DxR�@Ȧi�geVE��*u2pg\�*�<�Ύ�M�ęq��n~�`��t�n|lڰ���BZ<u�$�E[��]���F�\�4 y��7M�!d��D(��$�޴D0��Ol�϶B?�	�`��'@:�(�̓��y�U�B0�@���=�Dp�N��y�o���⡳��C% �4Q�w/7�y��Fp_"=��d9{������˺�y��̗x�jU�C �'zpZ�����yr���y��Y]_`��!W��y���2���΁-S�T�q�P)�y�D��j�B�t�SSU�Q�@E�y�e�J�� J��D�q��I��y�\J�R�@5�r ٳ�5�y�ϔ(���W$NA��b��p?���g�8Aw'�
���GP�+|҄�Į�OHբ.O�hS��{Ӭ6�4}�'��u��O��`��Jə�0h��É�>x"�8���(�`��Q����>���DJ��pf�����7Hg}��y�'��eExB+���) ��H�:n��XÆ �ybJ�U d  �$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ������}W�pI��럔�O�����!�6o���&�X7dD�F��O"�OF�ԟ0�*u��-��'~�Z*��m�Pl�I�L1��Ɋg����|B�Ӡq� �(þ=��jH%Faay��"�?1��������T̃EmE���M�$��?k���O��$;�)��45v4q`��_d�,�Q��q.C�I�D�j�h1�7r� ņ=m�v�O����&�')������ �*K��Q�\":Et�r�'���''��1aEP�G#LLӷF	�e���	�'�H�b� qԴp��%'d�Y�'���� � ?k���d�'=��P�'��BIW<;�����(��:Ǔ"Q�|r�dYZ� 2�"$\�
�AB�<�M>�0�-�t�'$2P�TL�7;1�l���0`�u# �)�Ɉ]�����`�(�ƊhŠ%iff�	o6�O)�B�'Yd��a�o/M�$/G�~D~}���   Y    �q�5�oN�b�ǐ�o��h�"LO�L)����u8�.�6.��Ȁ��'���!�@�,np��'��k@  ��*��v@Ȭ�7G��$\*�h�'��'|J?I��Ą;4�dHӜN��� W�!�B�I�x2x�ƒ�?'�@�aF+�Dp�G�/�d�w�V�$XI�!�� ��(X�8��'�O���%���v��C @��ct�${�"O�xP&�D�\\òϟ���8{�����=G{���?���;J|�z3���jM���c�){��|r����I�	�$����8H�8���|4~B�I	# ��g�֓�~\Sf�\'{�PB䉋AW��I����t�RAL�T�,B��I
I3E7���@1m�
�&B�Iz�8����+�~�X��FC��;b��E���}��锠7� s
�>T���@��E�*�r�'�a}�	@�Wt1a㪗���k!\1�y��V;m��P#E,xa�����yRF�8�֐�P�Ipc��I����y����D"5�	�jz��g�*�p<���	!QTڸ��i��7����E!݊'T�I�1�2#<�'�?������ ��k�K�b/�i��L�I��(q"O64�2a�br�Y3�I����S�"OblK��^�:���A�*��[�D}��"O�D�!��M~M	%ɓ`6�+�"O$9ծ:F�ج�Q-
��u�$�>�6�)��"�j��B�"��<Q��ӿ ���'������'aB�|J~"q�R?�hL�"F�/˴,B�g�j�<9pN42��@�L�5l����-�e�<Qc���9�(�!���-s뼨���Be�<�G�H�sZY�sH-:���`�d�<9��̅1��0�j��)�ԴA��]�,�������O6��k5V0ȁ06Ɂvi��(%f�ȟ'���)�gy§+-�(�+Ō��0�0�˞��y��
_H��Z&Kړ'f��;c���yr��7���Qǌ�&�x5�b��y���zL�T�U�zRȈQ�A4�Px�i��P�B1
�kM԰���RG8$D}2�J��h��= 5�33Ʉ��L;%C	.#�9�	럈��	B�L�xr�ćdThm��/�TN�C�I
��!�5�͑x���� �}\�B�	�z���K��w� �b�2��B�	0{bPs��*O�1�`�#���$q�'���2)�� 	�p�J9?�4���'������4����O�kCL���@�H�Q��А^5�ȓ簽Jĥ� <�ܰ2��-2��y�,17I��]^@�cn�i�z�ȓ'�hM�3Ğ1S$���G�3)�9��b�t�և�,.*����W8D���O��Fz���B }֬���;bB���G�W���I.;z��	���%���$��#���
�Fe1�T�?�Ht��"O>`�W�;b�(( b]5�ư��"O�y��*�
e���3P�[%[�m��"OF�¤���,����� ��iW�!�䜄v%*uX ��e��!�㇊�e?qOn5F~R�0�?i�`[?� YsU��v����M�h�|�����4(�(8�7!q1Ҥ�Uo�
�C�I8V\<|��#�.+Q�pBr�&yS�C�I?+����/�4u�T}��-V�8�hB�I�X�Ġ�aK!J>HQ��i�WP�B�:b�L� �u�dsI��N� q1��	�@��}rS�Tc\�j�;F��=� ^:7���'�a}����D>��Ui��%xũ��yR��;6�p��F 5Ƹ�����y�/��R�e���Q�8ih�g���yr@WLX����	9��ɡsOF��p<a$��(I��e�g�E��Bq'��r.���$�|"<�'�?A������sX"� W��&Ic���%[�
�!���"2ܤ��Kܐ_%^Q6%�)IO!��;�t08�	.麥cu��=�!�c��l�雡7���ɷ@=X�!�X9�����˝<`��|a P�n��?���?�g杏Z�Ez��I�B����f:}�D,G(r�'�ɧ�{�P���n�����唸s�Ą��'�4|9�Bá0Qf�C&�ZH�,��
8-�3�^�I(`U!*R�[��\�ȓm���Pu��{��;�pv���J6��ޮ�|ucr��XmX=�=A#���)0���O�T�� ���&48��᥍2P����K���"|�'C����T(V���ЧC�7�\�R�'(A;f�cҕ��HQ�
���a�<�tJEd���� >B50l˷��`�<�F�Z�D�>�H F�	m#q��a(<ٵ"�jk��!��DR��d�Q!�z*�>QA)�b�OzlR+�-+���Qiܿ6xy��OR��,�O� �`"�.�"# C�'��?#���a"O��s�̒n�z�8$�U�Q�!��"Of`�t��T��!���F�#��:�"O.(�7��?���zpԻ],��p`�'��<I�8M��` QoE5+��t�B�M?����w���D�'�S�#��̚��,P� �h���%D��Y1�'1�n��L˔3o�`�4"#D��Ԣ����P�	H��t�%D����l�"!�&�4�C?u�b�C�"D���D���vH�p�V>���?}R)�S�'�x��w' k�8x��[�p���O��O��d=���+,H4�p�"W�A��1�(���y"��=)W ����Ϫe�0H���y���)���^�cID�0��?�y2jХv�����U�p�*��X��y�a!��f)1Rhrm��3�'F�#?A4#����c0�ԶH
P x���/U�vE�G<�?	L>�S���d�F�0yy� � A޽SJ�$!��V1U�"w�Q�|>�Xƈَm!�d^<\BUJ�J��!Q�-9����6�!�䁶�M�&�3w�`<1�F �i��𤄲r3��Jv�K6NK�iQ���f7`�����>�`��^�]�p�CQi�+(��c����?����>�ŁO=K�^4cH�9�����J�<��$��c����$�:��8z7J\Q�<a��Ԃ�ڸCs�֭M�y���AK�<�� ��&� ;�H�*EHEf�o8����ĘZ��-:#�9<d��)�.+V���.���S�����j}�l�:$V���J�|ų��Ե�yB�"_ҬA��"Ց����t���y2��%Q4mѥnX0~�`��K<�y�.^�_�J��@5u��TrԨё�y�)`����Lץi��!�
\1��I�HO�,%�"#�0mKvd�A ���R�>!a��?A����S�S?Qi1C���(�	�mC'��C䉠D
廓 �o�������TY�C��* ��h��Y��Y�"˻bC�ɽU�ܝ3Ԭ[�ww���B"K�.=^C�I[����ה�Gďq���x،��ÎD��F�9b�LS��ڭ_ � @ b:l$��6�D�O>�O�@�A�I/b�*�%πx�L݇ȓ0^28���Ymp(!+P�t���5m�Ȳ��

J��R �TX�ȓ���9v��-8|��$+�6��(�3�|�
K�
z�7�YhA���RI3�g_N�G���žn������Y�����e�S�Mk���>�a+V�BQ|�A'�2�ޔhg�R]�<qp�K�G�T�
�!P*E�дo�[�<Y�I�K)���&o��(`u�R�<15 @2!���מ+��QB�ÿ+�x�4ʓK�����n�%�rҶ��-U�����
��\Gx�O���'���}Ғ��2��`AwBx�B�<vSڑ!�D��SU�L0��ӞiB�I�WS� ����A�Hl��(8a��d܏h0�B"�ʗ|~��� ��P!�$R� eq �؜	l0�r�L�.(�F쑞�?�!rg��q�mS��<,�r�`Q(#}R�ڮY��'Tɧ�'S۠|%�]z��m2q�B�G��ą�F�8PFo�$	�޵���4D2|܄ȓ1F�AiCU�ɴ�G�
!��l|ip�ʖXx�H3��8UJ���e8��pa �$h=��*��@�Jx�=�b�	ma��Č�:� ��"�եu��	��* ��8�	~��"|�'��g��cy�Ty(F��X��� ����%!�*��AG\	z��Q�"O���D�
/6T�f�\�F�
�"O��է�+�4h���YF�u3f
O��s�zӄ���� 	�	 3��O>Q�퓲*F$�� A5wrb�9���E5�)����?���.�9`<Oa���ƝV�B$�ȓ ��Z2���`pIfM�#2re����x[S#��7�`�j«�kz���	s�`Z��u�����	�m�ެ��ɻ�(Oh�b���:���ak�d��D)��Oj)�s�i>���ß�'rxe�ӽp2���)	<�Ib
�'c\A�ĭ��g��d(Šª+����	�'
�=!�[���P�t�_&#�F�k	�'�]�#O�slŹ@J1����'���q�9.S� Q ���R��H�������ʃ\���3����������	��ֶP���?�H>%?刅'�'��i��KߩHw\p�<D�ڗo΋lf�,�&�4J��p�I(D���a��J8*yBb�۵h��qGm%D���3��63�L�uhg2  �� D�����}�� W������-?��Oԑ0��' �*7/ͷ#�n��U��f@�� �?�K>Y�S���DԐ�N��F�B�J��P�ҽ�!�R@?�1��B�~/@��*�!1�!�D���!�b��#��˶LC�E�!�DY�K ��ƌi�@�jǱ#c��D�%..q
��4H��ף�aYr����_��>Q�pND�y��J�9�|�r2���?���̰>7&ޜX�B<:�fX	��J��g�<i�Y�g��T�քӦ\���µ�_�<�W��	ne�)�5-�	J���s&�a�<����n��z!�˅w��I��`8�����$� ��mY`ױq�
���lN ����D��� �IS}��H]��ط�֖'?���$��y�ϙ��0!�f"�2T��Ś�
���yB�U�V])����R�J]�'j��yFU�YEp9 PF�Y��R���y�dO'C
�q���G�|�Y�CN���I��HO� x:��?Z��e�7�\%&䍀#�>1'�Q�?���S�S4<"��6b	�T $�(�Ңp�^B��-�F$�q�X�] �� ���r��C�I/[\�܀��� 9�i�"ϩm�C�Ii~	�v���]ZD�I4ox�C�I���7�G�bf"��$ȋ$�㞈��䖻��!����]��6TNh((uc�*��$=�D�O>�;�uy�M��AI�t��"+����HBJ��@$9]rԊ� j ����[����l�o�~Q�B�cq⨆ȓb��ߊd����#��RQ�p�����]���1J�#[���Z�/�q'eF�� �mC��q�@�C	܅Z�ng
����O���.{;pi`��,uzd���dB�c�!�����`bB Ӹek����K��!�D�|_>y{�C�XL��0�@ԣ|�!��p�rT0���	K0)��I�T��x�.7ʓL~а$�	Y��� "G���F��5Ex�O��'W�	Gf4sw�Ì`�Hl F(��_;C�ɞA����RCˌn�
�i��L4�C�	1YP q�$E!���	��)d~C䉸CbXqI�'�l����� J8�C�	Jx8��@E=��\�C>���'��"=��e�lb��Rj�M^RMʥǟ^�D�	d��D�O��O�Oa���u因L�a�"NP�x�Z�y�'��	�lҦd�J ���_$0����� H�p0�I==��$+�Ɔp���K7"O��)e�H�UZjm %��{۲���"OL��a�}�D*�� 1P��Y�B�d�W�'�Dm��XѾ�xW��	CIx�"�"6,\��'U�'7��Y��i�_Hq4BΌ^UN��� D�(�ɜ�S̀���jiI&ȋg�>D������s)P�!-�_�����1D�`�Iڨ)�� ;���y,1�rJ.�L#M�>Rp`����E_�ѻ�dϯ]jQ����9�'�v����$��ĉ!�"1xt�p�'��'ۦyˠ�ȺO2(r��άP
�'�",�/B,R1�LS�@���P
�'V"T�HN�a�x�z��Ikƀ��	�'xs��/-��P���c?H0��(AQ�P�E!�/�$����r 9R�g�'�bT��8���O����Hh���.��q�;9�Ԉ!)���ڝ�Ak�O�2 �V�g��j��"]�E-h�IŏנG�:	��ҭ|I
)��'���3�j>�3��č �ԉb�M1s(Q���W��e��O �z�x��i>�Fz��_�}�"l�vf@?y1�ɂƎӗ�y�L4wH�y��tR
��"Ĝ���Ɍ�HO��}�O\,5�����G�8�u��E&��=,����Od�D;��~�R(�
�bU�͓�o9����Y�b��$�/��B��=�U����<Q�ۇ_��`*!jV�-�H�@)��q�Rف6�Ͻ!��� D���<��^�(r�%�F�%��u��Ń29�����D{�X%�P��9hr>i�I9:�!��9��1R�6O� cc�ʘ`[qO~L�'��O8� ��O�z��dM[��(��PfG5, ��SѪ�O��O���<Q�OW5?f`�Qw��C&�Da!gN�<�d���;x�j����*���i�)
E�<�1���O+ ��S�5�z���I�<�҆� K���/[(�(�k(<����K*NP�e
��;t�z�B�>AS�z�O�.,)�h(Tz�=�`�3_Bl< ��O��D8�O�4���[,XР���E�/��m` "O$���ϴ-�&$��j�d�a"O��Je�Z+W+e���z3�Cv�<!���.2m.QH��L������/�s8�HB���1��2�T?xr2���_:����/NX������IL}Bk{Y�����O[Æ�� ,�݆�v�D}�2!�)	�M)@�� k�l��ȓ� �q�N�8�tY�(T.��A��5CbuJB$ΈFH�� ��ڙY��i�ȓL�ʷO�}�U�V��(3��O�Dz��ǈ�yF\�p�nN&wi�!j����	#3,��	�X%���p$Y�.Z5jY̪#�%#1"O��K�h�s�S7o�;�Z�rR"O �Ƀ�&q^���ϓI�R���"O�Y�I׹v�j��X�,l0![�"O�]!)P?Bm����!
��$��d�z�'�x�2���}(Q�3������0@��` �'e�'���Y��!"ޘs$�0��%K����\��y�.A:�J� �,�$_��q֌R�yr$L�`��@@A�!���y�!��y��O�,���q���_T1� ��PxH\�	����W�v���&b^>	G}b�Ɩ�h�&s�`ĩx�ؐA��5n���ra���	]X��q䯐�3�
�!���&<�n̓w� D�Bw�%qy�$ ���bU�m�4+;D�@�$hK)~N�Q��'Z8�Lr �9D�x"��?,(qUH��1�����8ON�Gy��V4M\�Җ�N�M$x��.�y�"A�A "  �    �  �    e  �"  �(  9*   ލp�F˸��%�R(5n�� �
"g��{�� �� ��a�����2G������#*
?#>!���>_�X�C7	9�"���p�zpX���
�Ф2Ӥ�;G��7*�{�`�P��H!%a2h�0��d�*�&���p��d�ȑf�`qRs�D5P��aF��u�d����ۼ�b�%�Bh��m��J����A?D�B!ǫ�i�$���Ҧ=�<`*H0d-��P�G-��{N� ��T�Ü
K�R���ٰՌx��(M:p�ye�@�@rD���Ⱥ��ޤR(�,S獋�\⡃*cX��ĮRUbAQ���;�hY#.D���P�C�T�Z�Z��H���L�W�+D�P�@�; kq�
�_ߨ(�6�5D�41A��5׸̓�a�GvA�O!D�x;���'U �SM�b,�a�b!D�pYH45��q��M������.D��K_/�,Q���T�-�fT��D,D�X[��R(m�j$��/T���;�C6D����k�`�q���ҳG�9���9D�$I��j�6|����:��U�K3D�,���G�V~��d�^�*�j��b,&D����/�$j���"�# {�y��'D��0� W�KMn�b" ��Ɲ��(D�4�2���yѰ�z�ϐ|t�y�wK9D��3f��+�-@��$fk��RD(9D��1�K�V�\��Ch�d�x���J4D�0�rM��L� �XD(K3VG"|��+3D�`i�"��6`�s�ĕ0����!/D���S
��@+��b�i߃U�ԡh�l"D��ȑ�������[��bmU5�yB/����q�&��h2MH��_�yrY.ޭq!'I�_���-��y���yЦ�3�mn��U�2�@��yBn1e8��SwK�qr�t���<�y��@..i����D#d�J�#��S9�y�
@N�m	Ǟ�ɆmI!Y��y��Q�}~& ��
�����$]+�y�E�  HA�-^(&����B��y�%F�T	6��-�|�PV��y"�ߤ�jf�Bfh�lQuE���|Ms���<a���uԈ(*�Y���ĄA$�젡AJ�8)�h��N�(��}�J�8!�̘F�T�OG !b�)By�D!#��0f�5�v 2V��#�CB�p=1��Rv4]��d߈R�L�*1dV�'̭�V�f��9�5��3s��X�'EN�� j��@�L�y����"O6���X0B
�MR�)[�iӜ��'�"���4u�2�4�.9������ʵ%	#��c�_�6/v`r�%D�lQ�&y@�5"V�T�J�� �I�%+rѐ0Oʵ�6����R>	jF�0���L��G�9�	�$�@B���H��瀟 :А�W���W`����i���e 9^�:�x��+1���ד9z�����'Sje�&(Ÿ`-�XD{beƐ~n�j����zY(	K3*P�y��8Dzv�8č�\��4nZ$8!��ϩ2Ġ�SטV���	�RhBR-e0��h'$ԙh�)��ǹ�y����{pX{� °x�
���Z! �B�I�m� W/.#�dP��=n����$�  P��D5\���$��|
�� |�cE����|v��iEJK�/c~���I�#��1T@�� か��֐��f��
O�Ybro">���c	A�MV8��DʱH_4d0r,�-iK
��SoΕ0�ў��p(�-Y
cO҂bv|Ԛq!d�|���>=KY��oLC��ӀaIx�<1J�gʨ�I��*#����t
[ɟ�z��D�(�3�i��n�0�1Nu�"|�)'<~5�p,EMR(%�"J��yR�ͧ�	I��k��%�0c�5eX|[Rϙ�<�T�P/s�9Q)��1'��W i���3���>��YI¤�32�} �#<r���>D4��DL��\�4�Yz��"c�y�6n��&���D�\aH@��� �x��Q�S�8\ўpЂ#_2�@=`1N)~��T��)f��i#C�&~��]�$苸$��HгB�T�<aa�I*_|Ta�Eɩ`:���2jş���C6����
��Qac�a�"|J5FD�#7� �0��%I��G��y�m�=9���Pq�ZPQ�}2�ʛ�]�fܒ��U�<a�7c�<Y�/���T��БBǘ�`v��?��|0��S�}��[?P�(v� L y�#G<A�&�s�F�T.M����'z��fn�,)$�IדG��dA�o���PWز�F{R�5��Z�+"CTպ����y��0:�N��B2Hj0�c�P��!���d��<P� �&0|�9�s��8SҊ�eNh�C���@ɋ1���y��ݳ=�8�� @�( A(��[{hC� ��X4��E�P�!0O]	5
v� �W�e��
"�T�Q�d�|��f�fܓY�x��z����D�b���
d�������Q�Q&�����!�t32E�1U�5a����]~l���X�0Qp�qT�Ϫg��� ��Y�?ў�9T+D|+���Nli`�ji�Dq���J�d`���Ͻ]��@�d�T�<Х�$@=j���C���I@����H֧�yd��$�t��ҡr�"|�DeP KFl�!E����;PoQ��yB��>+�������%���훍�y2#ӅnH��밄÷2��Q��镬�y�� ���˂��>�����N�y��/����M�4,� !q��y�!S�,����1�Q6'X(��#�0�yB��&�V��0&R1'�`��'D��y�@�5`�N���&�"!��Y�$
�y���)�N!Z�����c�
��yBDV�|�<$31���	�Ӂ���y2eD~r|�E�9m
ڬ"����y��Z ���o[,1o:m��K2�yK�B����v�*�,�;@��yςX��x���;�"�`uF�!�y�R�H���u/��WzbWܒv��C䉶r���/Ū0�,����H�C�	Z�^�rF&�
X &��O_zB�ɿD��< 7i��2k0���f�+j�.B�I8]�&���H F�-�V儆\>�B�	#;������j4��ץ�CK�B�.?$AbE��_t^��s�O	��C�IT]�<SE%H$Y�h���L<txB�I$?��h�,"��)�Ň�kJC�I%F�$��l�=n|X� u���C�I�96�=�!
�;z�na�nL2T�BC�	�7�	�+F�S6���
I7-��B�	A!��k���>йh�xB�B�ɚ �(@�A�W�r�}au��z�B��2�F�K�-�U��Ћ�A��C�9ch��覭L �X��#�C��&5��eؔp.  �PhՙrV<B䉣G�����Ԑ9�х�:B�I��,��eO���n�$�B�	�S�<a����p��9�F߇>��B���Na�"�L�*�4���M]�!�B�	.<�ݱC]> 9�v�	NZB��0D�(t[s.�?���:�B��nB�I2���C�4T��40���pDB�	>b�$k��0lV�n
'z6B�	�m�^�Xqi�
ilĊ�I��B�	�IIb!(����k�<H����E4�B��$
�L�K�9,�@�x�r=,#
�'�Z����B���E@W��T2�'_$XQ  ~o<�S�-�l:��'���׋ �5:���Q�M��H9��'.m�`�ْ@���Qǅ40�'�Y�dL\^�(E�+�C���)�'<@<;��w�*�b�@�1�'F���g�3����ƒ�y�fI"	�'����� Ϊ��$p6-Վ����'�r�Y�8ZB �<&e�}��'Yj��aj_)�>�I�˄Z����'��en�pŠU��!T�:�z1k��� ��(�*&
�H1���OY�J�"O�	�"Ã�v��i�ϔ�]��(��"Oj�q"��!cq(��}l���"Ot@�i�6*�6AЯ
Q|V�p"O���a���s3�!i���`ڥb�"O8U)6�8}xș��#UsF���"OF� ��4{�*1��b�0S�b�y"OVB�d��)0�d�A�D�<�[�"O$3A��;��b���N�P�"O�tv$yt��锧��-ܞ�G"O4`�7h!/-�-3���3�$���"O<`�+\�K�P�TK��l�0y��"O�����K�D>���Q�M�b��d"O�"�m͉��Y�Gk���"��"O�!�2)��rBN˕�Vf���3"O�	���gc�)���J�yJ�"O�xO�eo�0���81p�p!"Oh(�W�Z��H{0��/N���P"OF=#S�à5[T�x!����}h�"O�8	e�
8z(�䐲"�s' ��f"Ot����s�,�R�7D"�|�"O����ݱ%���1�J_��m��"O^A����7�6 *b
�D���V"O� �5zCHU걎��=Q��+t"O�ˤ�:���:ĭZ�F�r"O6|�4�Q�%e���f��D��3�"O�9@Y�ek4x"6�N�1�̥�"Oh	�p����5h=����"Ol�K#D�u��]�$O0$��%�"O<i�2MN&F\<%��-)C���"O���'f�%n��|Y�P{H�Qf"Oz���-��;���c�?���`"O��"�]�Cyn��0��{:����"O@������kфR�`'���a"O� �N
7;�$��#��	 ��a�"O�i��"�;6���f�U�H"�"O�؃Q�.1�
���L`b0`�"Ob�C ă-�4q@�^n�(��"O`�7h  "�![��&6�6�j"O���u�P���U�E�F\���"O�8���?	=̀c�O�4HVfe��"OԱ�b��P�x��C�J#H*�"OR4���#h���nU)�|"O�9�b>{�:�PT�Ϻa~����"OL��"��{ޚ�!�N� L��s�"OJ;��NeFʽ(r̝�w����G"O��C!΀�#��y����(�s�C�	-mGfl�a@��S� ����D��C䉔s4��2�Ǉi3� Ð	�i��C�ɿj��a@c��=0�d�tb���B�ɽi�H�!��ڃjv:}rT�@"��B�	2jj���+#Qv,�E�=5��B䉜^s�J�O��b���L8�hB䉲e�4�2a�
0�Z����~C�G�¨���l@�II��W�ӬB�2��r�G�I�t�c�0
�B�I�S�.�R�B���ےE���B�	L��9��_3��4�uB��ڤB��;__��;�D�{�()kD@w�~C�l�d�с���4�p� i˰C䉕 "L������0 v"U��~B�ɫW[�l!!h�'j�v�h%$/U�NB䉆rO}�%����@�����LB�	�-���#^�nY�i��'��ٚ"O� �$��EZ�p��i&8pQ�"O��iqHS���Ԁ0��%����"OXy+��^_M�d���J��>��"O>�p��.[
�@�I86� *5"Or��d@�*xLT!範�Q�� "OvTIf���^�6�9����D	NYrr"O
�q����T� ����Vh�9hT"O�ջ��[�x-0�Jחs ��Y�"O�yBD���0,S�`�^=~t)�7d�(�q��`X�����8-����\1F�X��$$D�T�դS?W���2o�-G����� D��d �/b�������3Jcp�9�>D���$Ӳ�BnX�x�.��=D�<ڣM�:���EX"�V���;D��H��6{ x����>	Bx02�M;D� 1N�^1� Y���n�b8�;D��qb� |H,C6I�;.X��&;D��
v-ǲy.Ԍ��D�;s��E��#D�����B��x�A��9rж	H��+D� X���m�xͳb&� r���a4�-D��
7�6s Du���ӗB,J��/?D�Ļ�-��Y͞��,9"�Ea >D� 1��L�h�q�ޏrZ����F6D�8'�]<��J1n�2v�Dȑ�3D�<���Ϊ'�V����.ifn�A��-D�8�@�D�Ay�h��|d8�2�,D�`'��"FvZ�z� �7]Td0q�,D�L��o�7&�N�:���|��H�c)D��"�ǝy|<�&��MJ���j&D�����
H5�EpW�F1$�z���8D��	�MT�@����	l��i�� D����o݈L�P͑��[�<�(&�)D�ܒ���P��ãR)c��,�-D�����1u�|�4�N�B�ȸ�4-D�T����Z��|a���ue¼�Gk?D�J&L8;ԩ�D�H= ~$�7b<D���`�K@E��\�Z�*��$
8D��R,�#F��pA�R��[�7D���$"J$f��5�K&#�Ay�5D���/�v*f��c�J�A�TP�J3D�x(bjѓM
2�9��ƘQM���N1D������-�ܑ(� ��6���#�"D���e�+W/��@�1"�H����>D�̛��|]�(�TEޚt�|\��>D��JI�
�0a�#G��l� D���E��]��:���`!"A�)<D��c�G�
2=�ti�N 
�6�x G7D����>�"�z"���~��4�Bm6D���A��J�tp�g��0{��dڑK6D��i`L�g��a��B�YF����2D��n�2!VuCQɌ�zR`��$%D��(!@�~�JWI̠!N���	$D��ZBAڜ �R��C`]�u�b}8��'D�,�'�"M��)����$��	���&D�����?�N0�BLm�Dk#D��'�h$��I��Y� �4��!D�0�C��>Lh���P�1%���i"�?D����ׇ&��P�'�!z��q��/D���D��.yh�X"�xm��g�)D��JCkR�8#�ApNەe��|�b"D�Ԉ��&K	�0�(�ђ�a D�tҕ�sFDLA�% +8}r�(D��������� U6k
��0&%D������4`���(�!gF"D�� �����W�LhjJ�/K��U"O.mp� Fb�i��	�2}��Q"OԼ�W�7v���dϑ�DP��"O,�z�KϾ�LXzvm
6�<�R�"Odh8p!�R�����@j��S�"O�L�.}���	�<V�|��"O����ýJ���+��[BD�;�"O����TU1D"��W������,�y�,B�_l	��+�9i� BqS��yr����P1A�OF�_Z�� A��y�E�=6P��Do��Q����y¨y�(M��M
�fOd0��J�#�y�K.:ؼ�81�ε^��a�7���y"��`�����Q�	@i���y�d�<}���ƩU�US�7�y��A��V�j�ܸ-���jZ��y!D�8>�AԠ�os����E��yBԗ>��q6�c�4}��'��yb�C��1�CM:Y����j3�yB�~��hS��M�d�.�#�y��7�*u+c�]�Ve"�X!aM��y��S+���bO�
S\�Ya����ybhƝ�줒Ua�/6�Ba;P)��yb�8Y�(�*��Vw�x S�LB��ybB��x�)��D�o�E���N�ybLG�ܜ!���(z�$���i	�y2	J���510$�����(v���y'�L`�0��
y>�����y�"��+!�ax�F:�|I7����y�$^R���q�"M�P^��7����Py�,���B ��:UXL��lj�<��̞����A�RV�mj&H�z�<9R+6)Z���`�%��`�3"p�<y5'X�,�y���ֲ(���Y��C�<�� �(cH�#��&]X�,�o@�<�EXX\=@�����a2�c�<A��W*k�
�"���fP�+�h�<��n�[:v����R�6�sb�f�<��N�w|�@�U�X�u�,p�O�L�<S \�hp8�a��Ї?sPk:T�HCP(G�Iݼ�����O���vl!D���U)G����#œ��m��N>D�\��� �j( �5|��9�1D�`�6�P;W H���E�i�.l"�$D���c�Z��� Gh�(}��]�@�"D�b0��0fuP<{aVx�)��-D�B%BS�&q���A�|���%D�z����Z�RT�2�;� �(%D��;�`

$����g@?K�<B�a#D�0k�IOW�J�hGݻ}���8#�$D��s�Z<&�2X!��N�hj*(�2�>D����XCp�A$ɒ-��lK ��y��.;�514�!$Ǻ�p����y���<C�R��eʖ<!��9�w�]��yb�C:e�l� �Ҍ����u��yRL[�g��0W�0���
ה%�'4BD�c�Bƞ���0wE>���'?����̾8Y�� �Q�p����'itt���XE��#1��n]F�;�'!Dts��X�r�N��ǣ� ��z�'q&E��ӷ"dUqlH���x	�'����5旄k�RA`BJN�y�x��'�����[�2�j5)���X��'��@�2%��pn�d#�N��(��� ����퇲�::W��q��� "O���D�3~K`y���9*^)�"O�0H��BlB��e��:�`&"O�\�ō��t/�1˷�V+T�D�	"O4�s�
2҈KWa��ֶ��C"O��$ڸ�j]�Ҫ�N|� �r"O�u�Ȱg��2P�uO�!�q"OL�#F�ܮv����[�$j-X%"OV���N·WV���&�	
)PsQ"O��@�GE-i�#��3�<f"O�M8F�%D�ȴ�@�?�6`
5"O.𱀈���� #/3'*�ss"O�A�PA�:�(�`���^�H��"O��A�F��oN&�CY�Z���a�"O����V��j�l
	h��P"O>��' ���LmR�ͥ"�D)q�"O\�R��g@�ux�L�{��%�g"OYYr&��2�%����Z�d���"O�@�!�eˢQ6�L&ǂ8K�"O�AZF/K�ߖ� �M�+��Q�"O�Q���	k���B�J�L+�
�"O���'V;��(xG�Ȍ�$��"O앀���6d�8���WQ4yz�"O�5£�¦-��<��F�LZm	"O9���6~k�xq�!��]b툠"O����m2x�z�(2�F�"G���!"OH����QxVZ��0���D �I�"OU�B�B�I:6-;BO')Ԍ�T"O�Uj���X�^v�����	H"OZ�zP�
-noX�%�ă�x<І"O2\:���-^��Hj-�5���z�"OT�#��2�j���T�#&�l��"OV���X�X�����2l(H�"O��s���(<"�}K��9&�D��"ON�Q���$g9(PIc$լ[D�H""O���擿@R����߲q I��"O��s�[�^���s��W	K�>݁""O��s!��c;�4��G Y�p	�"Oh�+������d�8��"O�-$���mP�sW斗A�DP�%"O�iu��i�D4�%�����1"O�%��ÁS@� �2��j��@"O�#��K���q�@�/T�u��"Oh�X��ٌV-�<:d)׿���
�"Op���C�}���]ܾ�yd"O��HPNQ�D��0s��M�>� 9�f"O|@d��?��ht��.��`��"O�)bs�àv{b�f��B��E�a"OJL���
`�����
u�$`��"O��Z�-I��䘣*̩IG�@Q!"O`��tN�hG`�'�
_E�dɤ"OPaA5�I�(��{��A7�<�5"OJ)��
E <Tn=y!�W�P�B"O�!�F_j��0J�%�8B���e"O@������^��G�ˏ<�����"O|4	a �Og
P�
�1V|FY�c"O����F�����E�Ce25�c"O�9�l#3����@�5
X� �"O��q/_�ظ���"FjD��"O6�#Q�8�N���.BP(�{�"O.����ۑ<�D���D�� 1<)�E"O���EO�j< �s�&B�d���"Ot5K�)Qv���e��b���
�"O�#�A�)O�Љ��؜@&n��"O� dqҶ���@��BX/}�J�"O����Hڞ1�e+ É��p��H4D�����B�~��c'�B�"��d�U�<D��3��M>������=hRI�a�;D�T�!�O�V�bs��')M/!�\7���P��5���X�HA|.!�]L�ȅ@Z;�(,ˠ�P �!򄔕H�^�ItŘ�ft�4r�78!��\�E�Д[��Sc��b�ח|�!�S�K����N	VV�	)�JJ"]�!�d��xIP�AR�aCfU�2�Ђ:�!�D�Ue|�㇩U
�J0KFR<!��=B/�����eD��	+�
,!�Ɏ2# (  �   <  N  b  o  �$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*��D˛|�<!`��
u'�H��J޻&�!�dυ^��ؑAo��%2Y�6

9.qOR�lZN��Mt��4�?	ٴ!m �zG!4d�Y�N�$w�N���'�����t���|��F6�X�EQ?$Lƌy͇#*�L ���,��� �� c����@N	o�'�!&�[-%�Y���sy�6Ož3�)����Q �q��\���ė#e�e`���|�<�(M�"y|� s�ޠ@ؚxr̓8�	ϟ4�I���$?Q&���2H�r
�{�h�$0��E�;���#l�c��<�i�1=eN���^/c���)���Eʑ%4�tʴnXyib8xFo�SV���.�L���'�a}��@�~�|��e��!��la6ê�y�J�TQ>�@�D>d�I2fbݮ�y��G�lw8�8�$�dBe�b'J�y2�(�D�{�	�*Ye��B"b­�p<���	��$(����]ZRX�G�<����:c"#<ͧ�?Y����� >`�VݫJ���G�0,��F"O�-�dEI��]!�`��{�@]��"OVx�"�X�IQ�+�[V>�C�"O�����J,��*��ۋX��ىC"O���j%��e����@h�I1�>1%�)��Z��iH@�X"'zz�8$�	=���'�
	{f�'B�|J~Ze�&]�� Y�E�-��`	A�Q�<9'H.,Q.�K��R���-���D�<yE�5.�>�Z�h�-G�&�8'��<ٳB>̈́�z�MN�̵ w��E�<���͗o����bDɲ@� �H���jܓ!����@E�OT-���ɶ/�ja�י�8ȠJ���,'�<�)�gyҪ�E�R��H�4P��`��'�y���[�>���@8�d8��?�y�h��b.��;Q���?VNpsP���y�-�`��
�@L���[��E$�Px��]0*e�3�Iӥ#� �ic�T� �F}�)֎�h���jc�^[��jU&ُx�P书kO�t��jX� ��*��t9L��yDJ6D�Dp�b
/o�	Ѥ�
��Y$�9D��v��:�2���Q >Y�3N6D��Js�P���a�gl0�T]�'�9O�qEy�oЊb���C�CL,H�F<"�����~�j���O�i�O����>�6�ի
H|���_�<&��P

o�<��L>B���R��W* ��*%�h�<Ar�۬{ �)ըɯc�6ap'.|�<��)@&dd�Ѓ���x��g��r�<q���2��2��ʻv *IK���g�$
j���O�HJ���SQ�2Q�]9hn \�I���MY����	M�)�)R+7�T�@A]:%��J��žS4!�Dˢ:IJp�HŬ#_N�2_K	!�Ǚ~�*�ҁ	�=R��(�l�h�!���C�L�����?���
-E�!��Q�����O�:1!H)�ՊLiqOjE~r쌥�?���h@x��C�s�
�X�I-���|����	���p��	�:��ɸ�.%��B�I�<�e���q&еR��U��B��n	�K$i^/~��%�c��-�XC�	��dHqAh���ʋSz,C�902����&�*z�䐪� �*<������e���}�pO�V���1��P eD�q5�D��b�'�a}b$+#�Fh1c	x�dD
'�^��y���:��̣Fi��i���`aL��y�Ê:l������ȦVښً�H[��y��}�L���@��&�����d���p<ɦ�	7c�Ȁ��R�WT< �2��	�o�"<�'�?!�������dc 	�I��$�e*�
{!!�$	٘��7#����qE
ík!�$��Y7����o��������Hg�<�Eo[�@$(ۅ-��i�\�<�fK3te���p/�Va���!BW��o���O4t��r��>r��(^��J�����S�<��J�)���n=���d$�Ř�	���`C!�N�x[&DrG�� ��)�!��$$!�G,t��KWOV+�,lKA�	�{�!�ċ<c�|a!��R� �6*Ʀ�i�!��3a��'&ħd��1e��w�qO�%G~R�?�r�<r>���E���Q��y��#(W�|����則	��#��Q��p0��$QY�B�	�S�RM'��
��hS�яXB�	���Y���ΈS�J,�5�L4M��C�I�p��Г�mϸ=?V�f����Cቇ{��s��$jH�}�τ�1x"0�B���F�}:X&7��|IO��&�L��6@�s���'�a}
� <]8��p�<��$��j���ۀ"Or����0��qd�!w�*cf"O�<id�%\q���mE/-��ܰr"O���'�]���Ċ�Jת��q�'�У<��G�:�|�9�.�%/ �B�g}?	f�����'f�V�(s�+'*&⩘(Е<�u�1D�TB�-ʊ lT0��<m��H ��0D�P�3��k�Dx��W�MBv��1&4D��c�&�p��h�c�`uv- Ў$D��*���m�I����V+|{�$}b�.�S�'� ��ͫk�lD:F����]�O|$s���Ob�D<�����ƟL� �8�I+����i�yr,-<Q�#I,�������y�ϼj�,���Oʨl2��Y���yR�Џ*���@�I8�ς��yRE�30J 8�n�!5��`���'{2#?a0L�꟔�SO,��e�� �/l.���A�_�?!I>��S���DG�V�v��/�E��1�b�	�!�Q.M3<4P'����;R�œ0!�dٜVV��bN�Vњ�0�ʂ!���1:��e$�d�	�,��d�P�*�A��(r�t���%�l9��DͲn+�>1B㪄�4>��r $y�����?I���>���,�ĉf�7zQ�9��m�L�<��R���L:�(C/)�t���-�G�<QaaܛN�~Mr�/��)�ҩ[$��E�<�5��Q�2�S"M�)��h���@8� 1���M�8�ٷ�!Y��X􅃑X��d����џx��U}�V�"2�ቖ(J�j��X��yR� `��g�����2�N��yR��D�p(�A�G�ϖ�ʐ�X6�y¡��\���b%Q6�HTB����y�gO+�P�Ӈ�gБ�����ɟ�HO�``��·$�Bu����%⒜>�ة�?I���S��+�;u�%�~�c�I׹C�C�ɒ}8��pMR_���ڲ�S�6H*C䉩[��X��ݾ1�l�"�Ơ!"C䉝M��J���>f{'�F,P'C䉜|�b�k�L^�Op���bI9UB������J�E��'H&zb�C�%��c�1Pr�	�#{B�$4���O>˓&�� ���Ds2�tkec��ȓ�<	Hƈ#��:��|K���b��%��
�A����@���`�<��^H �`D
�R���A��v(<!� L�
}��qF�G&��B�Ù&I|:�>Q'�Ee�Ox�z1�
�f�[�`��*"0 ġ�On�d$�O&T*%c�2k�X9 ��sc����"O�H���=5� �H0���"M����"O�$����%ԡx�l�HR��yE�,���GCíR���*I �p<�T�(
�t�_�G�`LT�8^��	�p�#<�'�?���$�/SB�+u� /e$��	gけQ�!�d�F�3��s�N	S�a	�G�!�Ĉ"@���r���[���nӫs!�$K'D��mi���f��U�s�Z<`!�D���4m���k���Ak���s(���?��i\�:�Px�1
�,݆(#�>}�˕bY2�'�ɧ��ڙZ��(<B�ݐ�ǔ�D~���J�G��g&詐�AGG����m�@�G*��Y�X�!� T�%��`��\���ZŇX&�p�{�LI�}��ȓp0�p�&tH��bQ�@Y�Q�=�F��)�<�d�cd�3C�L�7R�y��G���I|��ǟ"|�'�h@	�&��rg���Waދs����	��� �,�ĩF�=�n!5Ċ�4p�"Oڄ���Iw��ɂCҍj�J0z!"O�{H�9� xs�'ԪZ�H��
O.@��}0	�0�A�1;D�3��ؤ��O�  ��Jx���(��e9U�R�4�\����?�	�6`�$ Q 9m�2(鑨C$�Vh�ȓ),��b� ��hÀ��Q'젅ȓF�,]�!�.���#�g�#b<���Y�1gف~Qʝ��բD�����	#�(OѰg�[[t-@
֡˄�O~ ���i>��Iܟ��'Mb|!�k��M��ic�΁UW����'q`$�G֪9�X� ��]%:t�ʓ ���bTe[8B�i`��OE�}�����!:E������'Z��ȓ� �rʕN^ҌH �� EF���OBYFz��T�I�Oc���Sh(
>ҕ���@(��	�/낡�Iٟ|%���D�f抋D�`��(K�aJ=�2"O��p ���r}!2�3T�t=�q"Od]iai=B��0�u`�82qr��v"O ���l�P�0�Z��YXO�E�D"OPqx�i�Ŋ�.�?�P�#��d`�'�����n��"S�Q5o.������n�R�|�����IX�`	Uo	��<����Z�C�}�.�C7�H8�}]��X� I��yr�Ūu�l�����(���&Ϛ=�y�+�<z�%"E]�B%���kϮ�Pxb��r�v�)�GͿL��!�7D�%.�ԐG}B��#�h�F�1 l��y4<�i�+tn�1i�m�ٟx��wX�$aD �/L��2C��#$��Ăr�?D�HB5 �=I�x[�������;r�=D��b�	X}��Ф˯o�Xa�g�.D��#%bΑs�@`��� IX=I��)O08Dy�L P��aFލ|�tx�oP��~�JЌ�O�)�O��d�>���� �����:������UE�<I� ڄd�X`(Tb˵6�>a�4C�u�<	�"Ӝ=�F�� ̌9W����q�<y1��>t7��qF�E�;%��2'd�T�<��a��h
,��F/L	z��q� �I�d�g���OZt�h$`,'����B�;;`�i�H��� ����蟨$�������B�}3ESsO�9I��CF"O�\��'N/Z��F:��Pv"O�)�4�!�XT['���$,�y��ө1� X�וg����c���y§?}o �h�٦a<�8����'�b"?��D���(Y�	Nz�$��N��"aB���?aL>I�S���Y�;K�U��n�m�^��GԖB�!��*���B#�QM�]�TZ�}�!��T��)���%k��A,H�!��|������Qz6Da7%�
ǡ�݁C�2�Yv'�:}_����68���"��>1�*[�/�a���9��0aJ��?���İ>��e�6| tR��@3x� Q�[k�<��K>I��A+r��n�����Fh�<�&�L)�J�ӅN�(c����%\Y�<	�f�
	��DJGO��$�L�����U8�!��䐀-�V�#ǎ3 F�a 0�A�aP��آF�������Ik}�h_$����>Ne��Q�y�-	� �K�O�Ęږ��1
>���(�Vҳ��N~�v�Z�^�h��L���&k��@��KQ(N����L���7���9)�U"f�B= V���O��Dz����L(����C��>����� ���I�T���	ٟ�%���D��p%�.][<��P����0*�"O�����=�j�v��v�,���"O� 
� ��O;��h�H���L��"OJ%��(J�(�)$f4P1V�!�"O��KU��9lkD8�p�/�(+S�$Vh�'54�"���` �I�9!��lz�*��Q��tJ��'��'���Y�����*�P �!��)@ ���6D�8�V��cZ���Z���3S�&D�x9�k^?TABUQS�V��0%D����5:h�	��˔j��1$$��;ף�J�� Rj[!_�h�2�o��!Q�,Sc�.ڧA1X̣��v�(<h��7����'!"�'��5r�O �p��Th�esL�!�''XL��͓{���Yu݄aB�]��'�d�S'/�/5n��˵�L�)�n-��'(�J�)\�U����L�������Q��x�� H�l�'�:�8���Y�'�	������O$�%���$�Ev�ᐕ#�*�,�R#&�ng�$(D��O�d�.u�g≼����O�)@xa�+�?S�@I��/�l��q�'�l,z��9�3��(����Bl@�i��dI
�5�D�Ic~ҩ��?�'�HO��+$�K�>>�x�@W�,r�`�"O��嫛�[�*��$�Ƥp�����>I@�i>I��[}�) +*Lx�PЎc��YH#�w�RH����<�����$��OBv�͔Q�&!�p�W�`����\�E���h�n�8Ơ�{u�'�N@4
ֺ�.���Z�y���J�p̼-SC놪 r����'˺��㗵I���y���h�����=�?	��hO:b��8�oV?YXH]�BS5�t;�+D�D�G,R�3a��%TM~:����'�I��M�����$7n� �O�����0��c�bA�|�"`�`�����D�<���?9�O��ac��,7�n8АoȨt�H�@��fj\�R���r��y��",OlhaC�'�N�ȡH�km&q{��O%*�8�K���b,�k���X�l���O��d�>�c�ð}T�Zr�B?oL���ɂr���=�6F�Wㆱ���Z�k�t��łU(<�� S2g˔��Ѩϣ~Z�q�敲	�@%{���'1h����w���)�M^,#����j��@���I�	�O$�d;�O���Q��$U���`΋zm6�X�"OXi��ʚG�hXW�T�P1�"Or�H�DNT���͈��S�"O, ���I/ v&�a5�äD�F%���'B��<���ƈux��'��4��DH?9�B�h����'��P��q�ԍV��hRJ[�<Df-/D��ѵd8at�)+e��Oi�J��C��sH,<�7&ň6KT)q��=a��C�2P�R���֟#H2i��fZ��C�ɛHp,����#���s#�-Fx��'�"=�B��1*��YG�)��p����^�dݽ,� �$�OT�O�O5����%�O&ԡ¯P�]��=9�'ph9��-X�#Ґ0���I�HGb��'��ͱ�D<��H�����j�\�
�'��� �+^9i��l*���-[O���
�'��H�7��:�
��O�`T��{�{R�>�R 1�I�9® ��Z�_��m�'���.g�Ԛ����?E�,O��a��T�=�	�oX���"O�݊��*���6c��/M�(��"O^p���$2��M�1Œ�왚R"O�-	�FD�;��KvDժ�"��
Oh�i3�+:CvY#�3E�z�R�a ��O�AY��S�|��iQ�
(9"����[% ��U�O���0�Oz�e�ʈD��A̲��{�"O:�qDl�.~L���n�1��t��"O<�s��TIZ �!�A�f�!B"O>���M߱RBP�k%�L*-�JDXE�'8��<y�`�@2�v��MZ<u35��u�<�Ca_0   �)D�B����mX�����?sF	���?YN>E��@I�%�t�`$S�����=�y"L��.Q��U���sU��9�y"M��F��()f@[2d( E�Q��y����#p�9R�Z�Q�������yb��
I�"��擌 ���sD����d�'����H� 24�#p`���GȠx-<��s�>�d�O���<Ofhq"�2q�)96�[(Fe�q"O*=�P�ٲ:���M�'V |�"O��$A��T̂ÆQb��ٷ"Od��_!wͰ��G4���'��ʓ:�Pg�9r�E{5,��D��?��.Kw���$�'��e��сs"<���LG��VL[��' !�V�t��U��Ί�&�D�F��	W!�D�Q��	Fj��@��ځ�P!!�� �pD���n)���E�H�b�"O�A�$b�9
t�e��D�{���퉀��V�(�$l�i�##>��e�Ԁ�0�O��)�O��D$�O�zXڼ��ЃO:��'
F�^��C�I�^��
�
��;� 3t-� p�C�	�$�TY�!�G[|a1 ?C`C�({t�$��N�����Eßq�zC�	�bXHPy����D��af �0q��d�j����H�3���P�x�oʴvrV�@b�O�]���Of�d7���'���CO�X/�(2����+��C�I��H"&��w@ -jBI�rd�B䉛q��h���îU�ʙ��dT��B�I**��\�BͦS�p��lS;6��B�ɇx��U����X#��)@L�{���_�����o'}��.��aW �Xu�����?	��0<	v!��p���W��**�숹ĉJC�<����3$�����O��Hũ�y�<�b�ξ $�mae��@��lPTky�<�!o'1�P\2'耆;��E��}x���*O�uiG��<E��@RL�&����]����ğ�'��|:!���$���&�LK�<���Jm� ��t��\�
E8W�9teP�٢�Y15s��?޴��(�b>q�5Ϛ�(V��j���{�dU��E4?1��OvQ�v�>��yb�/�HDڗ��7��X�E�)V���������M��9� }�K&�I��
��UB �$P��%I��]d|�PO���'j�>�*	֬��cNrȈ"J�2d)�@�2}Be7}�b�����iC=N�VA��fؖ].B$�Շ�0d�����(g�0�����&P�,(#C_ �,�f�ޜ�?95�BM��F�$T}��Bs���x��;�˚I�|��U����-k����?]"$!ӡ�^��%��!a����'�~"�Į���|Γ;��m�'�^e
s�T�T
2�
����(��n�0�� \T0�H��#}�1����-��/��(�SO��?��뷟�� 1?��yG���~���rd���Sc�)d�����8�?�F=�O,$��̈p���;F�(��"O�	ɔD֟.��R
S�/��S�"O�h0�fP%4�r`
"�л-ٸq�"O��*���Ь���K�<-��Y1"O ��;�:E�uL�:./��X�"O�� DA�(W��\�g
:�l"O��v���J���2����=�
sW"O���P��	SY�`ɳ�f��"O<�I�ݧ/r6�!�ߗ��5��"O`��oJ9.�<�Q/İ>���K@"O�����̍m�BlZ��0v��=��"O������8��r� � ;y�UF"O␊v�^6f 3�M	&w�h*A"O��������hUƦe��ْ�������<��ş�3�R�9�(��'�'ߦI�Kة�M���?���?����?���?����?A6���]��a7� jf�;Uh$��'�2�'�2�'�b�'���'v�ݷeV��FK08-H�s�e�#�7��O��D�Ok�i2�'{r�'A"�'tV����Ļ���b�C� �b6�h�d���O.��OP���O��D�O����O����O�$ܾ����ªh�f��+�����֟H��퟈��ڟ��ß���ٟ��tJ�z��}Rd���g%YJ��]n͟h�I��0���$�I�P������zG�SfEܷZ\XYb�
M=\J0��4�?����?����?����?a���?���q��E��̨'�Y�M�ܛ��i	�'���'�B�'���'e��'�4����G��44�NjF�And����O����O��d�O��$�O��D�O�a��j6H�:��5��{��`���릁�	柬�I۟��I矜��şX����hL�?�B��1H�!AS���cƟ(�M���?	��?���?���?9��?y�#P&U^����k��N��R���?_���'���'�R�'�"�'�B�'��͋.+*����ȾSdL�sA��=u27�=?a����"�2�z���V��+f�N7�i�O���?���D�'~���*'�b)А$�J�\Qu�I5�r�'\�>�N~j���,�M��'@@h�6ƚ�U}��ʦC�0 ���S��y�O6��4����*R(���CV"M-��{W���]����<IN>�G���O�� <��%�[,I",R<N	�ŀG�d�<���?��'��S�>�\�OI�pF��$�{\���?Y�/ �*:���������<OfX�c�*����%UoV���T���'n��,���
O��ֈ0Ƭy"��O$��'��Iɟd�?y�'�a��(8�y�Β'�����?���?A�6�M��O��S��Xw�X2ԠA�l)ĸ�	޺'x
ۈ�D�O˓��OfN���2h�L)S�nר$�\��/Oީ�'H�۟l���DU�W����Q˗\���+�%���O���h�<E�dj�.s����e��l�P�,�G9�@�,����O�,z��X��O��Gv�bg��in��p%�o��1�ߓ�I�<)fWY�I+�JR)FB
|�@ޟ,�It�����O>�do��@�L*,���!��G���P��e|�6m8?Y�C��<�Se�Ӆ����N->(���`��8�"��C��І��Z0
)�b�6��3�0G���'3�m�>�+Oj��;�	�D���BA� �Phw	�>�I~}��'��'R�i��	 f��D�s�M�~�J$9�X��kZ8s�d&���<���ɣ;xt	��C�?�ʙ�3�pZ�O�A�'?��'��?�XG��((���zt��<���<I+O����O��	m�'k/�  ��ES|��G�	?�L�V���TxpDQ��zy�O^V���@��'Z���+��&�����EKm�!�'�,�d�7,#$��jZ�$� ��S��#P�bR�X��u����O������)?j�[�k�y��a����O��H�z�7�3?�vʇ�P���Sg���SNhha�Xz��f�ß�?-O����W�JP���uƈ��dhıg�����O��?��	�<�f�6�ƙcD��8��x�4(�� �	�<��O����%P�r����A��<ٳ���6L�����>ڨ�$ϓ�*�)�'��'��	e~҂P��i��ME�]贼x
����O>��'��Iʟ�IϜK^9)�M\�[a�`�v��D���d�O��dw�l�O���vd�!~z���N	�zjݑ/O���W�Z�7-�n�S+��d~� ��i��W!�Q��D�l8�����7D�k�#	}<��A�۞Ib�{SF�O:��'��	�x�?q�'9*(ҒD�`��y�H˙I��1��?	���?ї���M��OX!�p�P���$)S�
��3qJ�$#�p�J��>��'���|�I�����֟����J4�(�)C>k�ޔJ�	���F�'�<듰?)��?�O~"���8QӲA҇[�D���fV56Ԩ+O���OT�O1����Ί�5�����%�-<(`g�+w�75?Y�ȅ�3����U�	Yybe�%H@�\"s���ZҢ� j^3�b�'ub�'���'w�I���D�O�x���R1���d��p%\%Qk�OX�(��Iy��'.�:OJ�l�y��T�W'J X�p=2�Mf3�7�9?Y�+��B��|r�w�b�`/�Gej):HQ�6,�c���?����?���?�����������D�fl
$i�	,^2e9�'���'�v��?q��?i�y.�-O��3Ħ�?e��|��@���?���?�2��9�M�O�����G���
6I:�( (`����'$�'|�Iɟ���ɟX�I�\.թ���3R����mؼ=��ן �'�&듭?y��?)͟��S �O�d�!������4r�\��'"���~�fKD�k��{� �F�&���I�/o�D�Xސq�ָ<��'��������Ʋ�y �Z��ެQ�#�)%�V�����?����?����'��$�����֪l/���^$"]4Y�#�?���?�����'��	ڟĩ"��a��xs��ҾCt�Q�C�yB�	�|�F��x�J5FL�AJ���ڍm�$�S��h�q�a�Ɛ�?�.O���O����O��d�O�'57F�Cs� :~�ڣ��#�:�O����O�$'���O
��g��q�@�1��,�EP0��`��O��$+��%��-�$7��|#�pF�OV�0�aJ�q�6��PF�|��'s�'Q�ܟH��6c<T�ӱ��:J�J�� �F�,�i���X��ڟ4�'�����$�O~%�Ph�)r?4��G�Bi�`��<�	`y2�'Zr�|2	ͩ{r��0P��g��ȓ G
��	��v@ ئA��t�A?!�'�p�!��?d�$Yd�'�`9���?I���?���h���	��%��K��F!��@ ȚWޞ��W`}B�'C��'��O���X�j�s���#�\��D�gj���O����OR��t��7t���f�?uz�A9^��|���,�J� C�.�O���?q���?I��?���Ttn��m�0J�����@ @+/OV��'
�Iܟ@���M�ޔZ`�.\n�j�jإ��d�Ox�$=��Ǹ.�ֹ��Ζ6����S�̢_.�@���?����Ek�Z��'u��&��'�(4��A��P��dIa��� T{��'9"�'��'��R� +�O��)� �Ir�o�O�L5��%��P��'�"��<�����d
���C̈́��h�SP�
1����iF�	�+>Ĝ�P�O2�p&?��;/RΌ�t��6q[ �ݿ�������P������I���Y�O�H��M�IHU�G�L�w* ����?���g��	���	ş �<��[��*%�0�S�hh��%���I���I;�xl�M~B��n�Z�I��	Ө<+£PL���#���۟�0!�|�V��ݟ��ɟXbÙ�D��ic$� <˔��QDCԟ���yy�)�>!��?y���	�<2�z@�##�JA�碖�R:�Ly��'��|J?ٰ��B�:��3���+@�[���j%��
>�I�?�B��'&.�'���C G�P���0��2��ᢢW�����ğ����'?��'�f���7@*UC��ڒCӤ}�����EB�'^"�'�O�˓�?!U��M�:��um�l3����H����:)�7-;?�dl��[�L��ٹ��i�?;�h0��`Ώ�7�R�#
��ı<q��?���?��?�Ο��JC�L�.�j���h_�Q�b81S�>a��?i����<Y��y"FUi:.=��#P�No����]4�?������'J�`1۴�~�b��]�F�9 HC>9��1�C�O��?ɥo^��>�xQ$�L�����'�����P8I�T�� ń�2i��'���'O\�xj�O��D�O&���3t\���l�6`T�2�(��D�>��'�2���%7̦%��)�������8�~�P�����Z�(�J~��L�O(�'T�����7f�8�S�!Q�f\����?����?����h��I�Xb��˥�6.^@$��C�#m�,���j}B�'��'o�O6�,%�T��Si�JfI6��#�O��d�O��ָr��6�1?��I���' ����Ip�y@ߐa�F�Y�d5��<Q���?���?����?��a7/n2�r+ڊ&��+#�� ����}r�'�"�'R��yB員P�! �dI+R8b��3N���ʟ`��^�)擯obt0)P�U�s�!���
�Aw�ʯ/$�;�$��N�OJH�K>�+O�|�GNơF����!a���&��O�$�O��D�On�D�<��\���-d�<�RjZ;̈́�0�ɨ2�6�I⟄�?,O��d�O 牫Hrj�
V�ӟG�:<�)R�v1hu�6�Imz�8���>A�;k�	�f��E/z���$�;Y����L��ӟ���� �	�O �Q�p⛠,�<�ҋ�� �C���?���2���ڟp��ԟ��<�i�-6�=�0.I�4�<���^�Iʟ���ܟ�ۀFYԦ��'s����+�4sf���@�d��u"@�w*F�y ���%�,�����'���'~�Pk��RNk`ً�$�k�̢"�'mBW��J�O��D�O���1R��߮A�Xs�nuԦu*��
Cy�\���	۟�&��OA��j���6�Y0�Q|��ĈT*Q�����4#C�	�?��g�O�Ol�WAߟdy��1
�nd����O����O`�d�O���,�0�̀�+�FH(AOW�?����c��?���?����'t�IßP�2��S����b�ߞ���V�̟����-�ZmmX~��Է=����~�3� 9a'N��tDS�vi�|�"�򟈗'xb�'���'��'b������Zc��Ё�Kh��I�'4��'R����O��I�Ką�ǉƠt� ��fO�!�8�D�Ox�O8����7Fk����!c��y��DF�V��]�0�Kr$X��%Mv�J�����Oz��|b�[N�I�Q/� '�Z���P�>�̱A��?y��?�)O^��'C��'bA���8���&J���)��.)��O���?Q���Nrޕ ���w�mҴ�R�42fT�,O܉۷iB1��ȱ���Sb
2c�<i&�}���զmm�(�#��0�I��Iڟ�F��8OL���L�(�XB�,�6@����'�'jX����O��|͓/�P�1蕯�*��"5_���I�����:V�M֦Y�uG�'4X�dU*E�����M�`h��pG�pL&��'��'3r�'��'y��`�ϔ��J5����U���OH�D�O
��8�9O���G�MQ�AքW�{�:}҆�<���?�L>�|
!ȝ'���7/��9�PԩŦ��	�(�4��	-6��@`�O�Onʓ|b\�auk��)�M�֌�>�
pJ���?����?���?!,O��'�Ą�V�0����2Qi��C�Zr�'��O:��?q���y��FE�ٚ����9��ѧ�	!Q��H�4��d�=�����O���Vm��'g!-�� ���Z�xL��'n��'���'pb��k9x�SB
|��Z�
Z�/R��D�O��$�~}��'���'P1OrI�r	C:D� 0"���\#�I�a�|��'��I�<�}o�~~r#	.��8JW���r�$�k�C;P�ީ!����*ן|�S�������	��T�U�P���g��u `��o�����yy��>���?1�������:?��1B%N"be0�q���CybT�@��۟�'��Oqt�B�5{�U�#K�(;�@01'I73����޴52���?���O��O�r���;�u`��H#.�SRm�O��O���Oܓ��ʓh�
� �B&P:����P�9k�>1���'f��ԟX�?�*O����'�h���/
�_��|��/ú��O�A��o�~����+RD����&�:�Ϟ/~�����)V��@��'�����T�I����I�$��o� F:2b����	S�E0T�ʲH�	����I��$?�	��̓d���s�J9
,���d(:P���	C����O�\I�4�~&\7����	�5r^��V��?�?yC�]�-=��D�����O|�K�KJ*P�gϨ3+PE�B��J�L���O��D�O6�XO�	�`���R��ި/�8�B�*v�vL@�^����d�O���5�d��+t�Z�ۭ���v2M�vʓn��e�u� ���4	���hz�3O�ƫ��("~M ���y�0�۱�'�r�'��'�>�̓mv��jd��?�%�q��)}ƈ��I���d�<9���'-�4in.�'�[;	�XP��ۗ��'��'�4,��i��I#F<��O����	������p9�`+7i�?L��';�I��4�	П��I㟔�ɶ%�
�F`��5<��(�ڝΠT�'5Fꓹ?���?���� �PR��%o���ؑ�7	�W��ܟ��?�|���9>w�xcw��, *~	������u'8��_�i�x��2�ړOr�vn0�dYw��y ���&�:U����?I���?i���?�.O���'9BM˧e�4E��i�.x���E�U���'��O�˓�?Q���y��R-HJ�1�%�k�|�Y����s�,��4��$Q{��������OF�.�.!5}��dT,3�u�7I��}B�'�'���'~��S�a��i0�6�X�1A�P$uC���O.�DI}B�'�b�'1O��	L6#�R��5+_�@�a!s�|2�'��	5R:�oZc~b`H�p�J@�3�بW�.D�d*������D埘z՜|�P�0�	���	Пl�7J� ��E�p�æsߴ��#f@���	Oy2L�>����?������c��$��@:&���`X�j{�	|y�'��|J?��5��9u�l�'Â?/��%)� ��u�^�0�Άz���?��U�'�\$��� 
ɂBe�t)�l�'N�.Mk�(�ҟD��ܟ��I�%?і'[��D[����BJ�֭�ҁ�<4V��'#�'�O���?y�F�u��̳�qKX����?�c���޴��d\/!�A���'Dl�>0����~�H��OA&�?�.O��d�O����O��O �'j}H�2a�0�*M�"�N#k����O����O �$:���O��{�,R��A�nː�ɹ�Ɲ5:)4���۟('�p%?� ������� ܨ�4 ���uM�sG�P�I�z;��'��$'��'�B�')��3%��.���������%�'b��'?�\�ta�Ot�d�O���L�F�TMy@��bml��W����Ԗ'���'4�'�	��KG�Rv&,d�r�JT��fLY���oڥ��'**�	�<�v?7�ε�c�{v0�33�����	�� �I� F�d<O4�)pA½;�����Q�e�٩s�',����$�OP��Γ	-�M�GnC#<s��y�I�1*�h4����4�	ߟ`2UE�����'~9�1���?��;>&(�#�ת��!�W�~fJe%���'X��'��'���'����5h�\�H�h��W?�0��U��c�O~���O��;���Oq�gN� ���f�D�H�Ti���<���?M>�|BA��;��,҅+�kA-s,�JuUcٴ���A�_f0�A�'��'�剮u�\KtD��|@�b��V��y�	��l�I���	�p�':���?і��<=�~�pG�6��@�����?�����'q�	֟����<�dOP DP�*��G�a�X�@�Z�JiG�iL�I$Ǡ��T��˼�w��(^t�լĎX�ԛ� şX�Iҟ(�I蟔��П�D���R n\�@�f���꬚��:�?����?��[�|������M̓r�5�dj��M�n��Z4��$�L��؟���%N� 	l�v~�|3��XL�(E��Ұ��;7Z� ���	�~2�|�Q��Ο<�	l3ǂ�O�V�{�.Uk�z�wˆݟ�	myR��>!��?����)��t*	Gޏs�,\��T54n�\y�'|J?�e��_~���Y2\�܂�,�F���2a�����f���$'�T�&h��hґ�7�#;�QJ�A�П�I��������%?��'X*����$�JOnƆ�+P��/J2�'�'��O���?�a��J*�0#b
U}�H����?��ʞ��4����
-̖�����ħ0�4�1��Cv9
T��!_f@4��Ry��'�r�'��'�Ҝ?A��?mh܊�η4�0����F}r�'vB�'E�Ot"�'A�D�$Y�5[�,zg��cA�,Q�b�'T�'��OB���Ӽi��d�&[5�0��D?��Y6��d�BCQ����ɛe�'�i>����n�s6�*�B���A�0���������џ8�'�듢?Q���?�M[.6��6��(��+��	���'������IU�i�6i�$�$PZ�N͇?漸���<�@i;^�l�H��I~�O���Ʌ��d����ȑ��V
>h��"�&I���' ��'2�S�<� 2����,}�<%��1�,� �'�H듨?���?���5O�a@g.�;OrT-Z!��2�PI��'F"�':�Cx�f���@��L�T�$��|er�R{�&�+G
�`ݠ���|"R�<���(��ϟ�������B�5s.���/S�%��j$N�gy�A�>���?����Os��Y��@K�^x�TDM'���gY���I���&�b>�#�mK8�1�%헒-��Xխ�HtHi�7?��*]�8���d��䓺�Y^�bS�@>s���"��x>��d�O"���O��D�O˓)���<���]��āk����%���h�$��	{����d�O���x��H��A�x�����DLX^���Of�b���U��?�$?��;<i�6N֧~�����:e���	ڟ�����p�	�|��`�O����5&M�h��C��r�@����?��Eu��Q�D�'�1O(�!�䂁8�����KGΚ���|��'�"�'HD���i?��
7�xaP-ȍ:�:�bW��t7ddB�Î���<���<)���?a��?p,	Bv�yp'=h@�2���?9����^}B�'���'R�ӡ&�Ա�P�&T2�s	� B����O��D<��~: �!z$$)W-�(u-� ���t��p����r�.�����O�]M>��\
E���Ӄ��<a3�̪�O^�?����?����?�K~b,O�X���};�)(��\F$�;a�3����O��d�O��d�'r�� Yn�]p���7$�p��ƮK5Q��	"��o�z~�&X7@Jh�j��Ӊ"2��k�K�e:q����0�$�<����?���?����?Iʟ�:�1(�Դ ����]��U��>����?i���'�?Y��y�`
�*l
����W@�IbC��?������'z�z�j�4�~��B *)�8 F�ˋPa�,!Dσ��?��b��dE���ϒ����4���� 6
�5x���i	Jup!�Y�B���D�Ol��O:˓FE�	�p�	���j���x	�L��j�����J}�����O��|��Č�n�u��+x]eфPuy�-��Y8���i]��OQ<��I]���H�V��Ik ��	��j��y���'`��'�r�S�<aӨθG��������8@���P�\;�O,�d�O`��;���<��ɔ@�J{���r�)7+����O��WD���4����-<�Fy��'L���qS�$�h�#�-T�j<1 B8���<���?���?����?!2��*e����g�O �����ĘC}�'Sb�'���y�5E��)��K��8��D4V��֟<�IR�)��5?n`�iW	Ha��W�FC|��!6�
�u�&@2��O:BJ>Y*O��`�A&/r�T��CG����Ȅ��O����O��D�O4�ĩ<�W�d���M��'ug��Cנ�.ƼY���|�?�,O~���O<�I�à Un�ց��Z;_⼹��v�h�k� ���%!�'�yg�9:=���� e�4��&D��?����?���?)���?ъ�i�e�x�A�DQ�I��@C&�>^��'GR�>����?1��'�|�ϔN��1W�N0�.%�I>1��?���q���4��$G"H�LkA*�t�%�t#����dBk�4�~�|�T��ݟ��	՟h�����{/�[
*0�٣nGȟ���cy�e�>y+OD�d,����@���"�/�<M.� �my�Z����M�S�I��5b�%��J�%7�.�����;
�ԠX�捅R�M��X�pΧ6b	Jq��^H�+��J"�
��ɸ����4���������$&?=�'�|�Ĝ:6&Ze����+!��9@�K�W�BR���������OUGF�$g�|��Ëb�
�p`�O��DڛJ��62?�"�(�`�OωO��Aۑ
�,.������0@u�u����D�O6�$�OF�$�O���7�s��7v���v+����A+��X���d�O��d�OZ����D�OT�IH�
�ۣ��E�a ϖ5���O8�O����Pw����>!$�Xc�0��	!��V��F�π"f,��'��'��i>)�	�m���AȀ	3.t<[��(<�����ğ�������',���?����?��l�G�ҙc�`	}0 �APN���'���0��|�ɣhR���rB�p|H$�A�xz��'h�!!�.K�x���9�O�	��?�s�`�l�T��1puH���k�����O��d�O���Oʣ}��'�"q#whңi�.�0%��8>1��h��	iy�'��O��I"wb�xsTBё[��h�.� b���O��d�O\5��GӸ� %z�k5 ���]� ��m8A�Gh�Dȧ��`2X�O�ʓ�?����?����?)��v���6N��l�5�kGt�����<Y3Y���	���IU�s��LM+rm�X�cR"Y;��("D�ey��'�b�|���a��4�ubP�Q�(��d���h�%��DPe% � ��N2��Oʓ"Y}�F�ІK" �3��^@\����?����?���?A.O�,�'��l� @�����\�L���Yv�Q�.��'��O6ʓ�?9��y�Dt+�qp�H(z��S�/U!5��0)�4��dپC��$I��)kމbSJL�;����#с>i|5����O��d�O��d�O����O~#|� ��p�
S���D�4a����v�'���'u���?y��?��y�_�e*���� �q`��
q�þ�䓱?	���?)6�G��MS�O@����[U�~Űa\�=H�i��1g�q�'��'���x�I��%4��̓��^�Sp&��!��)Jbz�����p�'����?����?a͟�=V�_�^�Y�3�ۿwjly1�^��'*��'�ɧ����"p&`[j��L�G�9J�+�%vx7�,?��=��	m��� 2b.OA�򐮔Zt����'���'���'��O�割�?�L;��-#R'��4�T� P�П�'���Ķ<��MF�x��G/"�i�4��N6��k���?�����M��O�i����K|�fj���pDĜ\Uz��f ˟0�'r��'R�'���'��2\������^+vu�sI�I'(�'z��'6��	�OV�ɐ|���J���B�h��1`R(D�����O��OL���q[�Fx��	�+����,�8��N@�n��>8�,��'3�'�̟|�	�(��4ʤ��M����L{�^!�I�@�I⟀�'����?!��?y�AV=�ʨ�C!�@u2��1�^���'4�Ο���`�OZX�"�ϻ/��<Q0�T�#�N��'��G�vC��I=�)�
�~2:OR�ń
3��RFh[YZ�'@b�'}��'��>]Γq������P�J�jg�K�p���������OL���O�㟰Γ<1�����2��u@���,	}���ؕ'?$t�ļi��	�80���O4��tH�-Tx�)��]�xm�'�y�	DyR�'�"�')��'�/ϥ?����f�뒍M���I���D�O����O������d4��B��xה�Ej�8R����?Q����S�'q㈉q6m��-�b=�uCI� P��j���Mc�O�@���\��~��|"^�l���*`���8�LI#0|V�s�aß���ޟt���p�	~y"�>��}� =�5Kٔ("�!�k��O����?���[���ǟ͓\K��u΃"(�v4b���"@J��j"��Ħ��'� )x�SN~��w@�,���ӍaR�\{sJʸi�R���?���?���?	���r�b�%$!*@Æߍoþ4�$�'��'Zh��?����?��y�Mi�zXp���n.�cB������?a.O��[�k�b������	98��%�U�P�t�c�%�� �$�����d�Ox���O�D�4$�4���s.�A�q*!Yv���O��C��I]y��'��ӞYԘԻ��#�~��d�7�����Ox��(��~����%������ެ*D��p��9_�@8A2�ʦ%�'��D$	\?�M>	Rď�����(�{�|y�Ú�?!��?���?)O~:-O�5��,�d@�U��0�-��%����<	���'��՟����Y����Vf�"$8�ɢP� ǟh�IQn�Io�w~�AV43�����L�S�|�R0�'C;��e�,�V�d�<9���?a��?���?�͟�}k2	B�]AK(�t���J
��IџT�I柀$?�	柬̓H�nA,��!��֝3ֈ��IV����$s�4�~�'�3xh�M�	DF�Y��d��?�1C��P�N������$�O���C&�tJd��!F�1k�)ϥ����O4���O��=����|��8��R��z����k�:����A����$�ON��/�$�"7�T����@�<�@ɚs#�87�˓i��
� ��9��|���ß���=O\m�t��0x=���AlÄBj A�'�b�'���'��>=�7!�]R���5a�~���/7B*���I+����O��$�OP㟬�e.�Yz�/�9[zt��E�2W�|���ş��'a�!���i��	'nk�c��O+�y�� �C�P
f��r�'g�M�iyr�'i��'���'}�#�h߼	 ��J�B����#3剏����O2�d�O
��6���6-�PLje�2x,aV/R-v��ʓ�?�����Ş`m�����96�:`�H<<�Q����?<Hd�'yx �SƟ��֑|rU�p RG��w��˕c�[�0�'�ɟ$����8��ɟ���jy�>y�T��#�^�0�ތs�и��`���?A�BW���Iޟ��"�*#U�� v^����h��(�,�Q���'�\k���?}�}ڝw#�d�s""6*�i�BK��n?،����?���?I���?Y���2a�vAZ;K�������E������'��'����$�O�c�@����8�(�@��9dr$��6L.���O����OKVJ�F��Ё���UƦ��PH�Z��N�$
�PQ5�'�n�%�����'���' HqǇ0#N*����.&��'m�V�dP�O��D�Of��%���K�ykU��(�T�	�JyB]���z�S�)�.z~����'QC9�(;w�U:G1���=2&��W�d��w�N�I+RX1��Y)-n8��+��f�v��I���ߟ��	C�SJy2��O��e�_�z��<t��YԨ	I#�'��ݟT�?�+O��DN,�ܱ�J2� �kCګr!��f����4���;+��9�'4�0�'RQ��AѧX!D4}���\7mۀ@��[y��'��'_R�'�Ҙ?� �]��@�(3�J��T,��.�B�s��>����?�����<����y*�!L�j|��eF�+�� ���4�?������'����ܴ�~��L{L�T��aB�$1�P��A��?��$F5f,��
����4���$��Hv� ;Ͼ!EL�2�~��O@�$�O�˓L��П|��̟|�D�<�0�rE� 0�TL3�( S����D�O�� �D^]�N����	V�a�	R�r�W\%�'��x&\���N���*�3Oj��S��l��L����`	��'T��'J��'X�>�͓;X���-Fr�0)ׁ�0'):��	����O����O����1��Y��ɉV��`A�9#b1������	͟{Db�ۦM�u��8$�Ԯ�'lΒ]S�����q(%j :"�`�'�t�'���'$B�'�r�'�$M� �:o)n�ÃG�!nF��f\�X��O��$�O�%�i�Ob[�r��ikk`�ڠ(����ן��	b�)�S���,�$"5��&B�T�
�H�Q�M(.��'MP�+�bM򟈸��|�R��Q��H�(.��0�B�o����#�L�����������	Cy��>����
࢓O@�]Q�� aքy����?��W������ϓ��i2GA��U	b�"�l(�%D�Ħ�'�`��a�E|�O��C|�&%ajE�iU@H��]=Z=�'�R�'���'�b�S
{Vu��@��A�8.Amr�b�'���'8���?I��?�yr���~���oN'����1�J����?�-OD(EjӖ�]��m�A�G�M�~p�-�,�bQv�[�RFp�D����d�O���O�����@!�dX��B<��,qB�)�d�Op�@���ǟ��Iޟ��O'��J��ӏX-�YPb�D�VQ�+Ov˓�?��J?E"�+�9� �ۗ+�L���X@#K$	�@��6��9�"��r�"�O��N>Q�"�cHR��W�JI����󋍖�?����?q���?�J~�.Oր��!6$Z�(w����j��30����Ob���O�8�'.�gNr�,AKg�F}a�o�.kK��'�@�R�I�'�,AJ'"\�͟V0�ƍ�%l�6Z�b��B��?�.Oj���Od�$�O��D�O��5 l���:$j p�D`���O���?�I~Z���?��'�F�0$b�	i`<!�פĘ%�p����'��O#�ْ �i��d^����B�*�
��i���T?\��%����ɇ)4�'��I͟h�ɢ<���&D.Kƈ�g�Q
Gb����ߟd�	ٟ(�'A(듳?A���?-b���D���� 怌:z�b]�?/O����Oj�OKS�r?8Z�	�-~B�4򓨌 ���'X��%���������D�ZF?��'D�����.���OW/p�X�9��?����?���h���I�\Z��h�/�r�d @��Z}0���\}b[�d��}���y�
P�R΀�Є��%vTm F��)�?)����䛏R��7�8?Qb��ef��P��vd��	4$�N91�NC����L>+O&��O��d�OX�D�O���KT�Pz��:S��)��|���<I�_���I⟸��v�⟠�J �|�w�˲Y-"Iyr��wy��'��|���ۮ����_a�r�T�C2"⸈�i|��b�G��`$�ؔ'ءa����ȓҠ�=B��%�'�R�'$��'8�Y�l��Ov��S '8�e�EU�)��I!-�5���OF��'��'���̧z�BtS%�"q��I�4v.p �ܴ��Q,҈a+��)y��бo@O4djW�� 9��H�n�O���O��D�O����O�"|�F!ҕ^�i�3L_fgD��2i��X�Iԟ< �O>��?q�yIK����h��e
J�����䓵?�,O�T��#~��B���!��Q�����^�0�\�Є���<Lt�d[9�䓾��O��d�O��d0pk\�9��Nx��Hv��
j���$�O`ʓc�	ϟ���џ��O]BXʡ��A�t0r�a�]�-O��?�����S�I�(I� T�T�ic�L2�J޿O����!G͎G��n�<��'2k~��X�j*��Q�k������y ��I�P��ڟ��	h�SQy��On��2�Y�//\�#Bɛ.k��A�'���'#�$�<!��3!x��E� �-�^�`Х�0!��9j+O�0��o���]�d �RO���Sȟ���$MƆ@	���P8s��'I�I��|�	���I�����P��@�^h`��ρ�{�:�Ⱗ���'���ş�'?���ş��k���z��)0j|̳P��?�X���Z���'\��s�4�~�θ^�ʑ#�!GjԚ�˝��?�k9x�	1����d�O��$
�(��s�/8=�QAİCr�D�O$�d�O�ʓZr����I�҆�C/c�ISE�)F�N �2m
o����O$��4���(V������O�`�Dm06�SN\�>�m��!J��Mka����CU?y�'�jY��L��B8XIcȑn�t]+���?����?��h�<�q�`X`����M�9A�!�q���W}B�'�B�'�O��	t$��S�3�� � ��w��D�O����Om��bӔ�Ӻ�0��AG۫,f��%&�9N�>i��fմ{��O<˓�?���?i���?q���� ���!�uOj�C�^�C�2�Aq[���OB��O$��(�I�O*(�7��������:�9�3E�<��?�O>�|BB#E��(�c�O�:b��Qy��}�2����C1��us�}��
�ڒO��6.��,P�ҕp�ꊱ6��h���?����?����?	*Oș�'C�Ix���K0j>!�)a�dʄ5���'��O�˓�?Y���y¬�����*f,
`D%��F�R�bڴ����D��8S��.�����e��ŉS���t���E}�����O��d�O���OT�$$§Y�m���H��A.��zԠ��ǟ��I�����O:���O�b��"�܀��x�������4�.���O����OT���s�B�Ӻ�֌�dX�@�W)+?�b���#?x��r�1�O�ʓ�?���?��$�M r��iTQxb΢5��i����?Y.O� �'��'B�?Q郱XDb�ͦ>K6XH �)f8�	ay�'��|J?�;u"S9@�a�S�$m�8�wO��~'(�r�8����
�+�O�,�I> ���~�؅ a
�=%�	����?	��?����?iO~)O�����P\a�)�*|Y����̔�:
����<q���'��I�0���> � �Q�D:��̟T���s�ȐnZL~Zw^>X	p�O�d�O���Q'�)!��I(����T��E������O��D�O����O�S�G/�?}龁a&E�-k�0�m���d�Of�d�Od��b�D�Ov扎'9^�Z`
G�=k�P��ʃ+g�<���O`�O<���Q���lӤ�ɻs�"h�t��9T�1Y&N	��]����s�_�f�䴠���t� ,@E�ޝ3C�U���LpH8+&��!��y�`�{����Ɣ]�,�l�RPѴ
��$���8&���0�G��	�B	ˎiuzL0iV9�"a;W�L'��)t�D$^dpc�P,F,Ћ�LP��Y���ԕ��6�<P��	�#q�����$h�@ ��@l�h@x��].p��"F�+;mԤ`U�&5�t��:T�����OX��91�P8\�}�Ĉ�]æ��ď$�I�E�s�䐐v�d8B'
��j�$���[<wdh�E�$z���� �<��@�m���B!��d�D�*��X#]�F�����u�И��FP����2�(O�1{��I��\�$喠|��z��X���@���IYv=���L���e˱�
��(0��Ҩm��J��Z��8�rvIS :C��0��D����U0Q���p��1�����L� o��Q��N^:+�P����h��P�:E� ��u댓r��RK��>��d�ݗh�.���*�����Bg��t�b����O����O�Q!�$�%D�X�P%����I1�j"���O���D	��@̧�,�q�?��Q%�"U�x���Ry�'UR7M�O��$�O����j}�M8Xe�f�7"��8(7*ט1x�'7��F�y�|R�iO>�¸IU� �&9�1C���u��')6��O����OX�$A}R_���P,W��0P3�4����TĊ�$KOB���O���Fh�<@A�o�)T��(��L��j6�O��$�O ��M}�_����<ѓ(��d��Й#,D���4r��C�;ݜ�yH>���?!��O����*Č\>s�0d�^"�?����?q1[�D�'�Ґ|�A"�� r�<���pAl�?�剰v�'���I��Iq�D-��J� �� N��s�0�B����?�R[���'��|��'��@!7@*j�$�� �
5@�h 7��y ��'N���ß<%?5�'$j�'W8t �!�LS�m-ty��Yy��'r�'���'�>T*�9O.h��]7m �����
$hWW�t�Iߟ��	]����	�OT1t˃!l��u�$Y�����O>�D)���O<���+�@b�l{��ܴ`�.��B(��Q��?y���D�O(m�O��'��e�>vH�Pҏb
�%��M�I��'��'�^C��'��'��C�H�r|�"[~޾����?;�Z���	��M����?���9O@��I�@�͑u�ݲO� N�O��$�OJ|�a-8��{̧/�L��FQ�B���Cg&��|����� 3�4�?��?Y����Qy��Gv� qb���R���חr	B�]� �O��?���J�4a;uM�Q�k�A�q��4�?���?�j��Igy"�'��D�(��=hQ�
zެ�Cި'x�Of�0��/���O2�$�O�I;��/=Z�D+�k^W,�"A�O,���OvH�'?�Iџ`$�\@!DB4!3�Ǜ}�!J�(Zsy�G|8�'#��'"��?���#7L,&\� ì- �)�F��O�|'�l���(%�h�'I��ѳ�����R� O�!e�p�'�b]���������u��J�.��b��x9d��,T�$Q�s(�{y��'�r�|�U��🔐�\�0\��e�09�~����`y��'�B�'��O+����Bg.%�l!2�B��f@�k���O���6���<�'�?yΟ�Aؓ�@䲉H0L�"�PL��'O�\���'�S���I޼C�C��-����MG���
�r�	֟��'iHչ���Ryq���F�
r�2b���B��˓��D�O��D�O,�$�O��d�D��t��?<��3�k�g�n�Z���?�+O`@��)��M��(A�@�����7��d�O*��O�$�O��S��C�>��M�C�F'BX��d��A��ɦeb�"<E��ݰ
q�I;��/����A�ƿA��'T�'�]����� �-��)^�]D	�n�c�Ɓ!��-�O��?M���<���/G-��(� �;��� �����	؟��'��SH��_,B%AA'ąW��DӖm��zM>�G�i̓�?.O\�I�~�����l�<�⵩��8r����<Y���?�"�'��+�,�!��	+x\�e�%��&������O���O��
|�S�4p�ӑl��n�*�j�ت˓�?������4����ʭO�m�����ۧ��;&v�Ol��<I,Oʧ�?�ģ�xy�l�C��9��q���_1�?����'��I=%.F�'�ꩉ�2R�j��y��x���?Q������Or%>�����æ�]c��h����9�h��#-�f��y��'r���'Qp$���Sn��կ�+:	ny��'�	����4��I�Ox�$�myR-� ~r��+��J�sݐy{�jD��?�/O��d�Ox��ȓ��A�1�	c���Cćݤy�.���O������a��矄�	ş\��O.˓:�1����d}���c�*G�TH`��̓��d�O��?U�I�k����(�!-���B�kѓ *�Ѡ޴�?y��?y�f���ay��'��� Zt�s�]�%���{�AF$Vq��'.�ɒ<�@�%?��ߟ�I�}�Ĕ�Tbҙ^-�TJu��ynȥ�	��I��$�<1���l���͋~��O�Į,2�,�O��DJ���<����?	�����pz�����R 
@�ȂuCȡE���{}�V����ny��'Cb�'�XQ���'S�: À�,|9�H8�I��yb]� ������u�S�����~29��)/t�~Y�E��Ȕ'�R\�����p���bx
�|�^eA�CE�fGv<st(ϫ+��	֟`������]y�O'맿y��K�F��˂O�e�>1��k_ �?a���$�O����O0}�S��;��� 	��x�zɱRF������O����<9�*������ɟ��!w��@ӷ��$�$$�p��Py�'���'��h��O˓���W&z���2TH;{��XGK��?�/O�����m�I������O��������aX84���p ��O���O�p #8O�O�c>�ǡE�)Ĩ�RjT(������O(�d���	՟��	ݟڭO�ʓ
`�h�Kޱp`n��&�.,EA�:�������Orn�t?"�@�-�.��'�Iɀ6��Ov�$�OD�$�P}S����<���W�|�>hc��3$=F�((�]�\d�<���?i�F���j�����*h�|lh��?���n��IYy��'��	ټ����椛�hX1a�P\�v�՟D�	B���ǟT�I����I��|�'�
A�$�_-��9aIբ^���'�t���D�OF˓�?I���?��)���*a*���X6�l����L��-̓�?���?q��?a.O6�$N�?�r�FԮ 4�9@�~3 ���OT˓�?�(OV���O\�DW�#o��?
�4!�g�Ʈ{yl��E�߶
v@��O���O��$�<�'o��S�dr����(\藢h�0x���4f�J�d�O���?!��?A`oT�<�/���GM�c��Ի�_�r *r	����$�'�R��~���?��&M@YvkS�8\x#��F3�\(O����O��H5/Y�	Iy20�X5���b	$�!#c�j�v�Xp�':�	���4�?���?A��J����?H����F!abؐ�!�TZS,������������<�PK��#��l�y`1 G1BJ�$�O�l�����	ɟ���
���<��'�.N���U0]t�(��U�?1���<����!��ɟl����7BhYeNE+(ԮVd�?�M����?a���?9P[�X�'�B1OR��`�в?؜��K6h�r�(�Z���'�8�3�O�	�O��D�On�2�뇺g���C�lɴ*Ŕ=--���'�2�>�,O���<�w�F`3��O� �@+oK�Qj��,O�Ԣ!;OH˓�?����?)͟F=�CŏO�������a+��'�R���D�O�˓�?����?�`TMt���LH�(,�Č[�)�8�'�"�'kb�'��i>����K�`�&���X���U�c����tyr�'j������ݟ��@���F���8�xm���YF=��[��O
���O��d�O���|"�W?�ͻ�򥫅�^�-}�q�@�d ��	⟈�'I"�'�"ݜ�y��'@��Z�	�5�1%�%p_n�yD��k���'|�U�d�I�����O��$�O�U�c��I'�m�v�I�<��N�<����?���k��Fx�6��I�le���1�I�\;�0�5�'~�֟�s۴�?���?��	m��T�ē�'ůT��Q�2�� kan��	����ɵ�.����*擜-�\����Kތ��ʓ������OZ1l���T�	П��I���ĳ<��$���\�emV+��3���?�B�s~�W�������$�TQ
=~Z1���-�N�Cf�i�"�'q��'0����d�OF��B��37�J�2���A��!��D.�d��h�������O��$�#A�����Va�=0��7�8���O���C}BY���	OyR9�lI��Cy�AjǢf���a!X��QSiv���	���I˟��	}y�cO"��5C�o^##+Hli@%�f{2�>)O4��<���?����� �M3�B@�v��b��L�|�!����yB�'�R�'G�W>іO�,�	�:-!����!�X�6YЕ�˓��R����Ny��'��'ѸM�',�}(e�E0d���JD�0�R�'�B�'�B�'��i>I��8�kS䮊2��h�k�s0��$�O���?���?-Ĝ��M����(-ju1 `� ^kF�
�cDHb�'*�V� �I1�ħ�?��aF��oC�"�&��Cǂ�"����O>���?�1� ,�?1J>��O|Z#�Q�d�Fʪi�&q������OF�ow���'���<ie㕃MN��f��;n��R�m���<���L��b!��O՚���LI'rk��
B*�+T/Z,i���?q��iW��'���'��b�p��
H�ńp
"J	�l��bF՟hhp�b�,%� ���]P�p
C�ւ=��DoA�h]���5�ir��'��'B�O6��O��%V$�9��Ol8q�eTx����9���*`����f��O���Y� ���	vMI5Q�J��`�@7�@���OT��[K�֟,�	sy2�0,1`��)1B�t��!���V��z����D�'��'��?����݆+��ٚ2m�%?Ju���F��?9H>���?1��\��@��D\"�r��l��_"�������O6���Of�����=(�]��(� ��hd�$XN��?������?��p��1��w[<��&ɟ%��|�SL��N~tԢ,O����O���2�	�q�ӷ`*��I3�Q�3�6 ��)F=h��1��ğ�&�4��ğ��`BA��'h��j��"�u��w�t����?�������O�I$>���ǟ��e�_�"������l�|����]�Iџ��	'O�2��O�I�|��!ΩqEBI�$�B'�u/0��Ĵ<9���W>M��џ��/Or5ň�Ka�h[ /ƽ1R��J`�'��'����'��'�1��lyэE�2�Z@�g-:}ߺ����'���e�����O��d�O���>�`G�L���s$ =l�r��d��?��Hܝ�?�N>����'�8�k��R�~E
�YSj&<j��7�sӖ���OH�D�O6p�>Y��y�!�J���ဥ�w�D�
4�?�L>�A+T:���?���?����XQK鐒��%*qo��?����?I&�x��'���|��R�4b��R����|�Bh���
�ɧq'1'�\�矼��N����#=>�hf[9�X������?y�xR�'tў�͓�bY����boJ٪�ꄴ]8Z���'������IƬ�+]L��J��8���P�B@G��
��uJ�\��װ�8ᤥ[+�?��?�������	'!��e�S.�pBDa�W� p�l�8�?a��?!�29O�<ر�*rnB|k����e��,_�d����ӡƲ|MH9ـ�Z�d󊥪���2%12������ūv.Z�p�T�2Q�ͤP%D��KY6�J�*X����q�B�#��5",R
����@꟦ �t�[SH^*�eA�(]8�6�+s�H��e��q�t���D��HO,���#I�=bH��
C�ܔ��e,�����!�p�'NB6K�f�8�I��u���#R��X;��2'�įg�l���i�38!��t�"yff��&KŸa�����\�C&�6/D��Z�/*����#c0��#�ͤz��Ģ��'�P���	�'dlЯZ��2d;@*ι`c�h�$��$`\z��̘;�a{�� .aAC���Cڼ,�5��I:��}��G2lOZ0I��''2�i4�A�� �����JX�Z	q��d5,O��f�_B��cCZ�q:l�I�"O$�O��fT���������H�����<9��B�G���柜$>5�C�ߔc�2 �sh�gJ����N��?���?����eD4� ��Y�������m��r5�#L �@�n�7��׫*��,R	Iہ)X�Ī��w�c�'H�h�ˣA�ע�if�^�]�!�>�'k�ɟ��	J�O�8%k"�)]e�!��!K�̨��3$��bw�F$є�(R�[�/؜���$"\Ot��=�P���Z��%���C5w>lx7d��7H� T��>���?�O���'#R�i{~]	5d�P��d�B���h}����gc�qD/�����nҌ��O��6�U�Ę dd��L��m�Wݾ�`��w'����H��	�
�2p�uOA�ux���&yna����?A�O�Ц�xb�hA@�3@xBPc��:~\�qs`a4D�|����,m>T��*A�l2��0� .�HO���Q#p&�_	�I�f �*�����?�Eȇ�V�'�B�'��	՟����L�+ޒs-�,C��A�`�1Q�i��Y[�h�R����
:LO,QR!G�x�v! ����O{�a(װi�4A�٦3�~��O#LOHz֩]�,"�Y��Ir:Tkſi�<����?��d'�Јq&��
�*\��8�U�7~!�$�;bx�ф-jp�I5��fQ��3�O��i�]g�O�Zւ�E6���K�.P6e����[yR�'�r2��8X%��+Jͱt�:\xZt�� �z��х�:a����I�eIh�)$.Ц2�� ��#�i�R��R&��G�h@� ��=����@��¦5لb�	l���Ȏ�8�
���J7���<� \�����*b���+�� V����"O2L�v
[�h��#�:/զ0��$���d�<��+�����'b��4�L�&-�D�#�R���*ݝ%C����O��(y�
mX# @�IN�����D��Yk�RAM�&��9s�����V��`"�4P!�	A1�i@�lU�(���'�H����zɱOfD*a�''b�v�(�+�IP�NP&���T��h\�k��'����"|�'��Y�C�ݡ\��U8բ�>��e*��Mk��i��ɵ,������lpp��C[�GC2]�S��n����'[�����O0���O6Mȥy
��0�d�$:E���RR7�Z�;���>�nO��N�<y�4�| ���z9>E�0� �ƹX3�D˶���d�77P2�<���y� f ��G�4�����Þ$��OfLo۟hЃ�>qp�Z� ��f�Y�`c���r��'�xdص�PP��GMXp� D�{�Cl����'��|�ڴ@vyq#�(EI�|�R�ϿX2N��ȓ2��!��J/f^F`���E�{�����R0�"W�Z�!�W)]t�0�!��m���	[�&DL�'vN� �&�ƨB䉶HK�iD�
i*m�V�9(�B��4L(���!MY7�.Q�l���C�ɯ�D���̡"Dx�#�!˴C�B�ɡZF�d�F�����%���H067C�I�@�uv�N^O�{�H�� �B�	7[=m2�Ax����iG� ��B�ɬN����aKσbs�$1�ψ���C�	�?H���f�Q5��L�#�)M>B䉥y�a�eT._J�̸g�B��B�ɚ\1*�� ��x�Lyj�ʔ� ހB����E�2!�#��%1^2�"C�[dB����e��� S�"pC�M`p�0��^ >�� �g�vE`C�IHf��TH� <�A� N��pC�$ˬ�����N��0���ܒ*�C�I�^b:�Q��J"�d��4��E� B�I��05����d�dd�4��6�0B�I'�t�G�@�h�Vt0vK1qA8B�	�n�&9ð�*	r:�H�IHO��C�IWH�SvG�sv�1�dM�W��C䉾TOD  �v7H������@B�	
Y/�� a��W��Sr'�:@B�ɉ@W,17��$��5�)I�VB�ɉC������:~g�U(�'�`B䉂3.��PD-L�P�A�v�M�mK�B�	#d����ʾ$TjMI#c�X��B�	)6��h�b��4��*��nԺB�	�#����A/N;"�T�7O6Wk�B�ɖA�P;Qg��OY���$�
fbxB�I�Vy@�j�#��őB���LB�ɹP>��� JLbi�w�*�B䉍wV%9&�>n���@�ظs�TB�ɺu�`�չR�r����pR"B䉗)�>e(�,�1@*2ܓ�NC��C��<X�\��l0��E�7/��C�_jT�G���!��0�.C�ɃL�;�fW5ed.�Ab"�n�BC�&(�������R��� gC� .;p�C�L�.X`ȅ�mZ�w��B���40b�\'aF���ԍY�/7B�	�et�E��͍a	~�8s�
-��C�	�:������V*�I�X��C�	�ob~�Z�/$	76� Vʐ���C�	�AdL:��
m�H����Λ�rC�I$%BQb٘7e8-����T�>B��;`{T��Di�i���k� X�Kk�B�I�;�,����C	)����ƊŹM7�B�)� ��T��Q��k2핍���"OD1�G��1�rݐ�c�b���P�"O�AC ϑ)֝�b��7�!k"O.�+�O\0q�Pк��S#N�T"�"O�x0�"K�4����W3 �J�"O@܊�e�0(��;CjH]�P��"O�u���KᾥT�� ]�R���"O�8�p�ՀB,�5nպ;�6��"O.x�Gj��}���#A ��"O(A	�����L�+�\+�"O�����Z�%���1B!$����'�0�L3<"��Kӿm�b���'�|�գ�E�J($��w����'����GbYgЌ�Ήa��@��'UJ9�
A�G���2�/3Ú,(�'q��a2�I�[�z-c/[����b�'��Y23@E�^Y dHEJ�)c�'P�勰�N��@��B�\'���'���:3Ϛ�+�#�-FX����'� m ���vל��%��0_Ҹ<��'�&�#�H&{@q�Ġ!�Փ	�';�ѲP�G�c�*�I'���Bd��'��Px��
�(�H2� �
B��}��'`6��� P�u�4Hp��F1Z���'�6���B�%��)��L�A8�@�OhICB���p=IR��7��z�ƍ�|��#L�Jx���c��&�|��6S�6\Iy��?�}�v	�i�<q�HێZ\
PQ�mY�x3�"ѧ`~��[��b�{e�OA�u�!K +*���d�Z�(3ai��D	q�ܳ�����>��M@����b��%���@�Y<��U���\�4�q��A�Ύ}ࣙ�l����OP]kB�����˷X8r�z��#��)��sނ���T-�8;����ۿ�h�Z��@�y��|x�ͫ��(GH�y�@Ɇ?��P�%d]�9���b�\6�M˰WO���[����QZ(�)񩃒QV8���$ zdb�ˈ!^2�u���E!t@Ĵs�&4�����>��쨢JK|e��r�A?�Ą�SV��K�$U.K|�F�ӝKI|ʓUD�ͻPD�H�Q�/UFx� ��%pʸ����&L��	�B��5��k���J("
_�k&ލ��:�" D# ��Im���Γ.�h���ǈR�(\�w����eEz"���j8X���E*L$�+�~��	7' ��7G��<t��bR��<aဉ|���#'����<�%c�zܻ#�Ac^��*�g����܍~}8��
U��Mv�'bZ��z7'4s�XU���a�<�I�B<�B�J�<	'��5�:%�O�;��QG�ˊGmD1N��k�.Ƈy}�A9��\�q�N�L���"je�ͪ����Bv6�!©� M��c�"�O���3��8��*`�Hfr�2�Q�hĞ)P��W)�-�T�i��'�r�	L/И�?�A` �GkD1Q�
ޠq� �"@���Ob �QPIZ����]�C��'ê}	��[�Mi��� �N�_��=�'�dZC�E��|B��Zy�P��f�G<�i���&�R{ 1�f'����l|�%�B
p@���šB�u��"O�h+��K���m)u��#R�4Pg4!}��'E��9`�/�3�d�!{��� �V�0>0A!J�c!�=c���#0jQ>(��p��B&�HiV�
<���
�pa@E�fn�!���xT� '����>1�	�a7����(G�=!�h� O+哣��a�Q�ّjl��P7HK�k%:C�	�x��u��l��D��@�	4>_Td���ڷ�~R�3zJ�����S�..�E}��``F���@4��	/�!�G�P��ѣ�d�T���Z�~�|T� ��/;`�I�'�v�����D�'�*q��G=U���UDP!R�j��ӓER�z��+h1��I�Z�[ �S��nTX,���H#D�����ar�+�$	+:���!�I�,.1�s� �ZQ?�vƇ�CF��A��
m�� �=D�x�A���f�P}�w�]hq�$z�疤�N�@V]�D��Dъ>�>-R��w�<qv��=4����ؽ^)��5D��V.�qA���3%4Bd0�M�;c�r�sסЕ{�����+&n��HO�e*��
"���K�$�J�Y��'��+@�Ԥo&X� �A( 	P7&�B�6��gC݄ �eC�LD j�a|2�W�VX���C?r��Z�≇��'��j�I��|!z�e�i<^����.g)�tX!�O�&\@�Ap��P�̘[���'�Ĩ�#�{��y�u��Cb>�($��;;���7/�&\ET&ӎC�̸�3��S��y���7Pf��M��;�����ǈ��y"HA4M�\L�g�F���� hKn�`��+E�|�h`[��ھ����^w�0�bEߥ��'r����6<�h�'$�%C2H�� �xÃ�2]��d�ɫ7�R�� �zi�o�4S��B��;!a{��Y�"(4��J_�b̶��k	�O!�q�� �H͛��4�b1�-�3=6���%�3�.���D�n��]��"O
�;��Q�q����D�D�]����t:O�#ǈ	H�^|�(�M���F�>�(��	Qh��b�\�E���A.6X�"Op�饏Ѓ�@(��S�r"�1���X�`���9g(�H��L%����'rqO�M3�k�1������V���'��2�.;[���K�A��dB��oO*RO>؀���c�)�� ,���I�5�9�0���yW�$����X<�#>!�Ɲ�d�o�#{�}j�kG�h�1Z0\-B���D��j�����+Ph�<�V&D%]���숏{ ����d?�B嘾dAl�S�N� �0Aks/WQ>q�7�Е}ن�Ӆ�c�~�u�/D���uL�f�hX��㌏	3X=[�`��[�f�Y�)F�<���Pc�1 �z��*7�7fZ�艑N��d4GM/�O��
gLN� g�]���o��z�'�,���K��Y�U��p�ψ���=a��v7Z1��I�`�J�����Z�'���H��5#U��jE��!h�4��'E�(���Gry��Y�"ϴD~̈́ȓ@�NA[7LC�
��}�g�C0Z����'}��c�l��AHިi��>I;�I6��:�eɫG#�@(>D���N֛Ū��"�
|��6�S-l�n��`������'�0m�0c>c�	!)�S�E�$���C&�58q�<���4aZ��&Lq��ٙl'x�s��MҠ)������f�'b:��4�\�7H8(@	�\��xX�7L40pi]���'~+�ɞ'`�^p���H�GS�(��g� �j�aƱn#��b��W�XŠ��=i�,bQv��)ƘG�*�3f#�>�^�� �<I�!�d��+�M0L{�� J&�Xq�!���]I���!�H�$�bt�&L�4w!�F�����n�*#�6\sdnQ�}y!�Đ�|��ك� ��2s �2�!�d�"���$J�{��1�#Ix!�%P�����f�����%ʣ(R!�$M5;E�T`�!V��A�0��	!����Q��rm�)�$T`��_(�!�dX�8���QҩV�^u@r�ĿR�!�I�CfC�kg���%�?o�!�D=mDt�6���2\B(�Vi͎P�!�dD��`�g �4|J 4BBW$[�!�$�u炝�J� b^ȼ@�B��T�!�aҪ�xS%��8^�uŁS�o!�[h`*�	N�4^�����Ƅ N!���
c�d	�
˛j;B|�B�ȃZ9!���~"�jFK֎
@T4F?�!�D%�|U��Fu.��6��W�l���yΪ�I�c�$P����o}��؄ȓh�$�̒�2�4���o�ʙ��}�f<!��
&���F�؈v��A���0�Z�,��T�#��Gp4��ȓ�H��u�%l����) w���ȓn��u�p��(#�V8��N��;
���� P8�E���y׬ܺ�ŴC8�ȄȓT��(�wa�wqXM��lR6y����ȓq\�qzC��+	VE�FjŻee4ņȓ8a�Ak�@X,^k�x��B��{��ȓG��jդAr�@��}�j ����|跃�t�ds�蘃0�����4�s��et`�z f"�ވ��S�? f�(��^ hᙶ����P�%"O�Q
�n���Ik�)ϴ{*,��"O\�""Ĵ-Z���h�_2X"O��1.[r�ܰ8��|p�А"O�3��:y��҇��+YG:2�"O􋕭�=��<�`MS�R3*��V"O��wޤ���T�PC�"O��b� 	+@\,�Ǭ^$���"O�ܘ&!� ��b���[6�K2!��@��X@qL�"GWPҰ�;v4!�P�#v��ĉ�Fb�3���U�!�Hؼ�:�N�A\�-9�`
�&�!��!v"�YZү������g!��@�48��!!�Ү%��- �bĻe`!��A�F�8(�m`x
� S�
S!�$ԋfr�dȢm�DP��Q�g�!�$S�a�L\�I�Q90����I3!򄏯R��!ZWȌ"W;$�J�m�,9�!�d��׊�b�*@�[d�sE*\�p!��ϔd�X|�1ɂe
(uIǮHgw�p1&o$�O������t�Ȼ�K%j�}�r"O��
�/��I"�:A��W�~�<�0��𲵨� YZ�����w�<��%�x�hE���Zj��cF�s�<yr����, �:o~0r�p�<�Vɕk`V! u��D�9:d�k�<$DH�xh�dK�r�@�Zu Ff�<�A���(�����*�X�Ԯ�^�<���U�󇑏�z|�`V�<�`�hsJ��ы͟CB�(SOU�<�B�<^���3 (�20�~(��R�<!a֔<3���$��6��`�"K�<�3��
0dTs�Y�1
��h�D�<� .��m� ��Č`��]|��C䉔�¤���T23��,S��[*2�C�I�	}ʵ�R�]Eh�r��OB�I-k��IɳB� e� ��E��g�C�	�N�:�����0����*�"�C�	�-@b,������Kw��

9|C�	�9�d����0<{\̰�����FC�	�J8�(3��Y���r��I�HB�I�x��1�����l(\%�U�C�D�&B�	4U�\��G
�M�RA�6jA(\XB�	�f~ީ�u�B)�
X��GK5Q�DB����E��x$��aP�	?( B�	7WB�TEZ�j�Us`C�`ԠB�I7)'����'L�MQ���erbB�ɾW����34�H�n#F��C�I%s����5_�$9�n-Y'�C�I�Jl1�'W:9?h��g]�O��C��4�"1��nͯ(�$�p��ڍg��C�	T`�؉&(('^�t�>۾C�	�-G�1*3�ϵt��k&�קhh\C�	I��8��S�إ��Է|�C�I<	���'��)b�����Ed��C�	�6Z��R4��9P, SFĄ��C�I$&v�0jF���6�:�P�h����C�I-O&8�YE��b{���	�)PT�C�������ҫQ�TǗ�tB�#K�:u��c2i�*M ����3w4B�I�[��pS�Ƣ]�V����S4R�C�ɝ7��E�&�R�O�D��eP?��C䉫<0ɫ�p�Ѩ�ɓ�L��B�	E�v��եқ^y�8���,�B�)� `�[�-"�p�G�A$D ��"O(|���
	f��Yg-֭Y&�t	�"O.i��!T�V��!�"�'U\���"OH�Sb�#.9Q�!Q��3��O-``X����z'���! �}+r���,�!��Z�UFN�	˷F�B5k�)0=��I�DP�����e��4��,£�2��3��|��C�I/�H���{���kO*>�vO��yל��<�c/�$@U�!�4B_���	�L�D؟�Ҁ�_M��%�d%�D�d��3��,�BԀ�O=I�!�����)s��*�1YG�I�D������vh5���;��D@P��y��6wFڽPw��"0� �A�.ϗ�yr�N$�@Qj$���*N�83,�yr��?�x+�Ⓙ&�f��"H���y�\�OӈHc@o�,�����ã�y���=iĨ�
��"�P�B�/�yR�$OTD��==(�AJ$O
��yb"�c�I���ŋ6Ӝ�(�"S��y���e�e��.p�1�yBb,{�ISHR2�m:q��=�y�
�)��q��A�=��H�	K��yb��93��x0�� 	�(�!� �y���{��y�ĉ��5Ȏ��lϹ�y⌀�k��Y��\�_�u�'R��yҊ�
aJ����XG�c�M�
�yb57�4�U��I�>١��V��y�ϙ{���{#��F:���v(�1�yra�*��m3��]�J,�¡D��y�Í }���'P�Ak.�2Tn��yR'��Ib��7;8@2���/�y�4 ?Θ� �H�<508�	��y�`��*D*"�[�70(�Ά��y"K^
s���&)�&�2,qF�U�y�E��(*�N];5W���(���y�!�O�f]s"L�,U(X癁�yRŰ64�X���!�z�@�Z�<�@,����s�����[�{�N�#�D_��gf9D��ZW�ԗ]&�iKt遆m��=Z1�u�\�傞tx�dj�	�8˨��A�T�=d�@M!�Oz�aC��<�!�V�(�@T�Q)ڥ��]�r%RZ�<� Lk�"�{�/%/������P�'qj�S��'>��jWb�s��L�3�DLB�	�Oժ���>f�̌zD�S�@>`�ԭ[{�S��ybmݕ?�Ψ�!`X�)B2x�C	��yB�/2��A���)ƶ�a� ��y�g\�=�L!�TK+
a#���y'ѳC@N�I�hE�vB�f�!�y��^_��I3B9���� ��y���7>��0�6D?�4���@��yR�S�b��S��e2`���'�yb
��u���+�lЫE�������yB(�h`���t��
���5 2�y"��E�|=���C��mh�a_m�<���& ���b䗆O�R��2��F�<)���
��4�R
K�;U��"bc�A�<�wN�G_ ��g��;@�� K�~�<��-dh�6OD�"l��Q�)�}�<Q��7l<��L�UF ���y�<��L��b��#��H��
�M�<�Xh�abîZ��H�	2Z��ȓi]��t�M�����c��XI��5j�Lҥ��im}�&-�r��-��S�P�����'d+�ěD�Z���S�? ��rc�4C�]�cj�||t:q"O��xVK	�i{�����L�3�Z8�U"OF�8�mZ�l���S�G�H6&�i�"O6%�"NF[+TJ�i�0\#�h�"OQ��^?!��m��[�Tz��˰"Ox�	
9t�B�bmT���"O>��Z�`��@@�VVvna��"O
m���V:d�LU�E��+dj�8�U"O���v`Лr���z�IU$UPB��d"OP�o�2�&]QiD#1tis�"O�A{2��'XNpd)����<r�ap�"Oz|h�n��C�0q�/S"\1v�ǅR�)��I B� 9�DeA42P��'���E�������OU�� .���ME'>3�eR"O}���^�����&��9w���C�$��]�X��E ��@��G?9u���0�� =ij�٣"O�!���*�i��j�!<5y��I��m�d⁶�y��K�5��r~���E�4$f]b���1l����S3�|��&0��q6�	(َU0�oѥUg�m�ƕ �����/M���#G�@p�͑��E&	��y�/_� �̒��]i9.��� =����ͩ��!RW�!�$ڍ/��)��_0$����O�>��'6z��W�^
"��DLB��(�����.�#���#�@?T�t���"O���-����Jw�kK����G���.�f���E����L��{!	��X��"���~��ت�a24��x�l��:i&�K� I�
!�|z��ʥ7�(��j��$����'J����h�²�I��1�Z�����i kRB� dD�OLTB���.#����Õ8�Rpr�"O��(���Y�Y1?��U�'�>s�[��f��CT�|���D��퓉P�:=��H��}<�*�*S*�yRI"	xv�B4��.�@}�͕�&U!��kX?�ꚺf5�~�&�[}�Δ7F%�s`F!x��@u���x�I�A���;0�C�w����œ�8a��[���c��%xa�O��I�%ߐ��O�����;k� ��D,�9����s�'�`}!囬"�	-�vԁ��%
�����L��/X���oF�~�+7e� �)��$L��zä.��'l^1郗>�U�"CH�O'�3���$�&�r��!%b⁃�'�&�j�e�)dY���$"HZ� �{�@ �Vb����%�uF�;z-z�!��/�H��d"OlU��$�G�Ь��Mc��1�g"O-"�a��F�����[�7��i1"O��$�I^Q��Z%��B�"Oڱ�f�ٖLV�(�0� �+	B�Ӷ"O~������3��"b�8>���Hd"O�Q�F�&��<3A� BТ�Y�"O�����X�9��9�%��g�(��!"O� �17}�MJAk�7z�ڥZd"O���B�Q%� X"SK@	:��鲴"O���!n�D�	#!���j�"Oh����Jy�"��du�"O��1r�ťP4>s$�K��Ft��"O� ��,�*G%�g����"O��j2E�=~���ٶ�\�M�L�1�"O �P�U$����"bH���"O�Br��a4��D��)O'�p"Od	�Oço��X� �5"
i�d"Op��6B�%�jL� ߐ�,=�"OL�	��6����S� 3�"O�P��7Vip!S؁$��dp"OD#Bӫ5:��đb��ɒ"O육5�2Rv�zӎ�Q����"Ol��&)�+a�(LJ4-Ş>�4���"Ov]�PFԛ~�+s��;�e�"O0�����v3
�@��Z�D�ԃ"O� b�[GbsPXaF�ڣ{�6�"O��E#�x����P�V:k!f��"OvT�R-�Db̔�W����yK&"OF���/W�[#��3$dJ$I&��#"O�.�^e˃EBfq�//tX!�$�',ZAq��8]��!&c�,�!��?�X}��E�SSL���N�!���q\��� A'SA��8e	#>�!�D�9��ԙ���%���Е%K�m�!�T(?��]�3�*��d���ӄg5!�<j6��Q��:L$J�QRj@J!�M*/j@js D�>�J�	؂H�!��6��`���R.����T��!��Kb�@ڇD�*��[���V�!���R�	���5:�������
5!��2����u)o}t3�"h!��U��\H���v^�QH� �4!��y�z��6��s7��@E#�Z�!�$6^|ѓ�GDY������/y�!򄏸wR�����q&B�`�\�!�$Q�0b�3pI_3G1�\�A��B�!򤀚D>�84�.ˤcC�.M�!�䌢!X8������m���fƨ-�!��09m,\�1Kċ4*�LH"�Qhk!�dF�.O�X�G�I�@3J���EP4:f!�E�yA��3�͂��R 2ą S!�E�q ��rӌX�_P���¥Y@!�D�	 �h�ķ5��Pϙ�&)!��)3:5�	Y�j�!as�W"\!��9F������I�M j ��%Q�o�!��]���EHt�L�T�j��֪��!�D��E@ ���mDZ��QD@��!���%r�ؑ�\�� ɉsc�:|#!�$J!V��z'NF�U)��1S#��!�$&{u���a��;bLi#��F�!�$�4G&Ԑ�JZ*��=��� �!�d�n\V1�B�/*�"YJ��Z!��h�~M���?j�T;DDA/ �!�$�'g���G4oVnXK��f�!�$�.��h@vl�V���1���
!�d� �
k��.T� �CӵF�!�$�,$&h�6���9頍"pC�^!�d�I�~d���U�0��#���Z�!���@� tK
�P>�u��@�!�!�$��}Ϩ(��� f0�b���!��Vξ��as�$�j3��%6�!�d�DrsE�С6�!:4m�2c�!��U2`������Ѵia��s�!�$�3�F�8V���>��!R�*�0{�!��Y�r�@k����,����Ș1�!��S�{Ѐ8�莽C�b��K@�d�!�$�}B�I�ɥH(DQxg
;Id!��am�T���G�@*�� O!�$HT��\ّB��ctExA뎫�!��-T�,@�F�7� ��ꀕ1�!��qǌt0�oL��IS�*D�J�!��4 6>\����f�D�i3j<�!�A�>o<E�vD��u��2`	N��!������c�yy�G��sv!��n��9�E�d�-�U-ֳ_z!��ߥf�~D+��U"bȒ�
œr�!�āf�����D�((1��Caʅ�a�!�d�&,YD!Z�v$1�'�Gl!��z��a!���pvU�s��*L!�� $�Cj�+j��x�#*c�T�u"Oz�b)қM�č�c���ɲ�"OB1�뗝Q;�|���0�z��C"O���YW�
J��PwD����"O�]����_/���7�я@6�8�a"O�9�@ȥS""��lM�V
�u;�"O<���LK '����',?
�J�b�"O��*�e8N'>��F
�$t����Q"OԤKv! va�h�ȑz��!b"O:`�6�({dH���QÃ"OQ�@������� �ty"O�Ғ@�%&-�C�S�dZ}�P"O��qǢ�0�\3,�=9���$"O(�;�#@�uÀ�P��>�r	�&"O|��r�ɻ8}�qPH@'#�"�"Op����<��ƌ�ch��#�"O:��'��Itn#�رAl�A�"O2<����.D��u���2]�L��"O���t��`sF1��놡=R"5ٵ"OnT��m�>M�iPtK�5��G"OHa	w%~t,�T+��7�
,c"O,-a�7%|�I��ۜ���yr"O�4�vK�s��*@Iި�P��S"O�5
Џ3��u��(�1	!,I"g"O&l�ӒM�be�
Ǳ$� "O� ���u�^�׉(w'R��T"O^ ٱ�A�h�2� a�G�(p�3"Op��(Q�<��y�i�=X�$�@�"O8�*߹#~��9��;2�1ӂ"O0��Fn�+h��㗣��ta8�+"O� �R�($�P5��.8K^Q05"O��{��wI�bf��1�!��y" �,:w�mA�mR,z.,`��J��y2����yT`Ty'����y�D��u��@:tO�0vH@�J%����yr�/?����LP�s�F@@F���y2똎G�V�Б��-k^xJ�+Z��yR8#�:QX�㏅`�|�匎��y��O��К��z����ō��y�ŀRJ���I�Z�Aj��Ο�yrL\�6A�mR�ț/`u���Pŗ��y�bK�D�@%8� �0	�r�'/_?�yb����rAH� �'~➸q�O+�y�`N�>�( B1��q�|`WB^�y��'j�ɱiJ}�)aa	Z��yR���D�@�u�@!q#��y��G
[����t��ts����̼�y2CݏHi�-���B	m-p����y� �N�b�!ge��QC
�yB�J� ���J�:��=[�@ٿ�yr���J��q�,�8Ԉ�v���y2�O%f[�5k�6 8���iF#�y"P�/MZ]�V��%=���1�ܕ�y�J�.[N�i��4��Prb�%�y���&^�ѺG��*I;�oԞ�y�)ܞn�P1v��`��v&��y�B�n��}zA��1�Y8u$S��y�%���8�߲R�t\���J��y2#�)Q�(4��Ȩ6̰��J^:�yR�SZta2��ɴO��!e���y�-��u�(]3�ԋH��E*��yJQ�C����5(��&G���y�$\T;�lhP�3;ؽX%�ߊ�y"ĝ��6(@g�R�[���R���y
� L��[�oc�Hp��?tu���"O�Y����Sļ�򩝘;=�4�"O>��a,�M�D�t�C \��p"O�R hs����P�X��U"O�}�6
��Td��J��ADV�ؓ"O�\Vȗ�|Ai�X�vF2]J�"Or�j����W�}A@��-�Z�#�"ORC&������1�W�J*S"O&l�Q@Z�,��qp��ڶ�a�"O0A���L�g���ۅ�:.Ծ��"O\��� ֻdy�,c�ʒ�R�3�"O�pR���| ����<&�vD��"On8��ʛ\�����߯uV�"O�a ��˴`Jؔ�pm��#f��p�"OrY󵌗�=v�R���V_f�S�"O��[�KPu�D+���5_t9�"O�mr�k	�`����"O�6)KƳ^O���Qi�&�d9��'�>@[FD8j.Y�e	�4�ѡ�'����g8l�� 2��	 V��'�|�i�*�0��rB�5|tب1�'��z��\�z��h/��Z�'����w��)b�:}�2�֘e	v)�'&���Ti�!�yt�ȕ�>�y�`�8,�L�dSk�p����X;�yQ6���p�f��t@�c�،�yR,�H��Q�
�t&j�
1H��y�"�=@�h8�d��<��ym��&�"0�c�V�"<�m���y���=ƨ�fFR����b�ԇ�y∐�c���P0��Y:��A���yB��b}ؘ�&mC�b��0 �'�yr��[��[���
��qp �E��y������Q�̔(:;��T�;�yr��L=� �'�1ut@d�D��y�37�j<���t��	��͍�y��D��!��%Na�tLT��yrd�z�^52g$�)�6	�pf�<�y�
�/�B���3#0�g�ۜ�y�n]�
��w�C�q {'�[-�yR�Ǚl�032���H��k3�yҠC�G�V�bf�I>�=kE�&�y�	޻h�(a�w�K�x�<�� �y��8I0;�F�����$���y�)�n���#J�)3�����y�f�4FJ�!!�I>���]�y2.ѽ}�R|Z�I�v�a�AW*�yR$�1I\���H�NŌ	#�M�0�y">n��y9��ی5��-R4����y"nw�\���![�z8�R��y�o_�����U�RI:ĝ��yRak�p�\9"!��;���q��ȓb�.i���e�v���'���^1��rZA�#�^�*u�4e�77T&Ɇȓx1&\ S%vQ��Ⴡ.T�^��Q5��#�c��$f��@m�&@�!�ȓ5�2( 4��%bBp�a`�:<�ͅ�h���J�G��\v0���+`2�q��Sgl��t�T���1Y���&>f.x�ȓ0z�xc2&�3:��L�a�!'M�Ʌȓ)��v�,sH́Ѳ��d꼠�ȓ;�|�t�nK A"ȳQ����P+Pĉ��dP"s�V/m����]�<=�P僵PnB�i���.(,���S�? ���1� 8���Q��% ��u1�"O"LS��1��
P늝U��K�"O8EYa X�P P9��[�t�v��"O����o�8���#7WL@�7"O�qs��u�4B�Ad��&"O��.���FH�T �B]r���"O0P�bE8&"k�-GvD���"O��a�cޞ3�u`��P�6�<K�"O����(͚W�.�{,�M��"ON�!1��_��$���<�Բ0"O�i�e�8\V�Zu�V�	1^��d"O����Kا=	��d��_���c"O�]Zqh����t���T�=u"O�8�P��.<f���6%� !��Z�"O�Q%U�uSVu�fnӧ+F��"O�Q��Q/AD!�Ε�@�q�"O�Չ��F�F`�u�q��߰%y�"Oȹ����}��t�q��/N�.�C#"O�:���/0^I ��>,���r�"O�t���'!��.A&|u@(Ǵ�y2��^T�Q�A(}}�����yR���k�dɺ$JJ&i��T���^��y�͇�@Vɒ%�
N���Bݡ�yB`��¼a���:]dr�(��4�ybdU�Q���4�V��3��D��ybL��e�|4���ŀ$ppQ�H��y��G���B��9̲���I�=�y���-\M ���g?tR�Y"���y"�ݛJGlY���&C���2�.�y�g!bU*	��*�L��y�`]���`�T�y�ȍs1"��y��["Im8�P!�n�����*��y�o�.�X����`t(7O�yB�SQr�$
�m��^����K��y"�7�Te��b�&���1ʓ�y�E�?y���j�g*���n�(�y��V�G7�<���̒��9�ì��y�)[!���QF�� �d@3���yR'V8>LM��g���[`CL[�yFח#��  Up$�h���y"d�_pƀ�1�_ f��ȋ�O��yRE�?�� �*��|��i�!�,��R�
�J�MJ{�(�-FVD1��0N��[���gh$@�E� �f��ȓf!��a o���d]�#'�c5��&p I���4���-�
̄�Cf�e(vL�Q�xB��� �8X��|��xu����R���k�	p ��p����'��x~�W�O�=H�,�ȓ"��L�S���X�`�R�Y6>�!��zH�2���<�f�r�,��]�ȓ|�v�Р�n����D&�nE��%�yIW�L��[3`T�>����$_�2SG�0�n �"��"��	Y��Xq�X9!�.�1o݄X�� �ȓT�a�F�vN�M��Kٽ)�X���U����V,�#=� ��3�Q�S8���Qnv):V��,�N8��nS�����4&lD��D�6�E��+c����pK�iS�!�|�*T+t �(U�м�ȓaF$i�W
>h� ӕD�&���ȓzeX�ꀁ�$u��t�g�)u慄� ���h��K."՘2��nB�8��&���� �Q�`�|4�u-��+��]��S�? L�ԭ��_���U+W/�ʵz�"O�Xr�h��q��"�c�s��T@E"O��� ԕWL �ɧ#˷D�H�!a"O�l[w�&�4i�8 ~�Sc"O$�����YU�]�{f�  "O�R'��<E�@�*\�To4��"O�̹��^�
�.8YƩ�MFdD�v"Odl �䉝qr�u�4I�69Z����"OԐ[���&b��@#	M;~��%k""O�I�‥;J�92\/~��'"Opm�ʅ-����$n��_�I{A"OL�!`�<��Q���;�H��|���I�\bF���&2`Vy�G��Q!�D��9H�ef��nXfP��c��D�'�ўb?UH1��e~�V�̏`%6�S�=D�x��
F��zS�K�q��4q�;D�������ʉ{�b$;�D:D���#��Bp�!ǁ 	U��0�l9D��a�ՋD��\C�m��@b�:D���N�n)j(�ĳDPX!(�d:D����jM�g:�1ؤ��H}0��";D���c��>�n���k�"=9�}C�,<D��U�!pԸ�r���k��a�(<D�y�"��Μdk�3u��W�8D��c���F���X�_^т5C��4D�x3��6=lD���]�.�Ca6D�*�AX�q�$p�q�_�j%�G�5D�PZ�A�CL���A�`�
�O5D���>zd���#`̨� yH�3��d����Hi�ҍAQ'Ƭx����0D��3��D���� ϹU~M8.D��[U�@F�P<	����jFf1;��,D���c\�9�>�Y���'@�\�C�)D��P��D����%R���y�.4D�<�v��RS }R����L)��+1D�4iT���O�&�`�� ��2��-D�0X��_ -��kfT�%��D�%0�,�O�!Q�нXb�Ґ�X��'"O&��Dn��OM� @IAB��r�"O M��BB	J<�P���F:�i�"O<,	�:�*�k� �"&�L�v"O*(�#�R�"7v`[�nC!{��`CB"O��AJN�[F��GnC�v�q�"O)��&�4a�Tz�-�%����W"Ofq� �/�� (�L��#�ވ�r"O�l{�L��Z�9rퟃ;��L2�"OV��!��A�:L�@�F�(�Jb"O��y!��Q�P����Yq^��"O�=�B q H� �� ULhf"Oh8;�j�
n@� !ǎ��h��Au"O�}2r ԃIˤ�c4��w��e��"O4l�T	�,,�nl8��3��a"O$09`�Y����w��%c_�T�"O� I�&[Ҿ�z�i�'V��@�"O�y�nܹB4h�k*�(}�l�J�"O�I���6�4DsĉB�;�}p"O�����fe�l����D8��"O8�+�-�6n A�ʍ"8����"O8��̦TxV�CO�r��q�"O�\��k�M(���v���d"	B@"OXI"��)�+3�3LO&U���d)LO��q�iŧ]�,�-A�U�ꐉ"O����I֌F_(} `�L6B�8���"O��06bUI~L�'ȷt�*��"O� (��T���F�zt��@�&)�q�"Odi��ٞ����eE�@��<	1"Ox%���ʕ5�DԠ�E��q��`�"OPa;��	�{��� �kɾ�lH�"O���ʏ�F3��5`Y G7�""O@b@�]cN$9��C~Y�3"Ola�f���a��AQQ.зX*����"O�9;Bk�YH�q��M�!��"O�`׃DdZ��BL@(���"OhԉH��*p���&�O'4=�"OƝː��&��L���֧6�e(B"Od��c�P,I�\�éS�b�Zh�Q"O�|�eH�z��b���5��"O`���gc�D�L�����"O��r瞺#p~��!ӡ��ȩ�"O΄ ������`��M� "Od��5D�3 �l�D	Q5���C"O��*s⛤<d���ڭ*>+�"OL�A�"6H�2p:�[=d�j�7"O���qi�B����+�*|�d+f"OjTSq��B;�̒�f�؃�"O%h�i�9bPFP�vNU�3p���"O.m�.̈�B%�*67��ZQ"OvE�&o�"�h�)0	��2�̂v"O.��&^Y ���B�*����"On��#	 8R�Q
�G� �Ԁ@�"Ov�8sU�5�"��FH�]�\Ha"O��H$��(I�U�eKD�����"OjX��-Q"dӾ@�E���^��M�"O�8���4~��9��'��A�N��"OҼ蒯�|Z�Sf[�H���S"O�:Tp����� ;�8F"O0�V&�7i_6�� ��;p�^u���'a1O��2��@�e<�Xڒś�#D��"O6�:�	F<{\ C�7~[R��%"OFD��J�?3j��3��XTj��"O�2f@U�����εHj�Q�0"Ot��I�,�4��*��Wf`k"O(�+��j���!�$�1Y��a���<�S�i^=>��!�^+V0����kK�e�!��0}�(e2RF�r�Q�D�w�!�Q�?l�� :eB1*�Y�h!�䖳V�������
pL����$v`!�$Um��y5�^�54�(�L@�L�!����mz�������j�Z�!�d��t���ձ{�樳�T6{�!�G�.�
e@%��9e(��&҅M�!����uc��A�Ga�0��E�l�!򤅾X�h����jH5CɨW�!��2o��P��HէbD
��&D;{!�D$[c��G�͘C@X4�G#��"|!�"`��PVg�m9���cሇp_!�d݄KX*Л׀J-�A����m>!�$�#aZ:T�tDB�%0��t�Z�!򄍢m�Պ���{��@��D�!�D²sͮ���&�)4\���
��!�� TK�
r�d���NL~V]q�'���Ȥ�R)f<A��?M���X�'@��)GIQ�N~���A��(�'�x#���I)6���h[3�yc�'�љ��ŰsI(�'��
>=��'���8���#jΐ�W�E������'�8I�SD3e������=
���
�'c��c��*Y<�y�n�z�.�S��� X�[�)�6t�b���LV?��0�"O�dBt�E�V���u	����XW"O��
�����2GݲUϘ�g"O�������O�*�c�J�D(b"O���G
<4i��Չ2�fxQ"O�}i 揍0 1�%)W!0��a��"O���a��+};��%ȏ�{��,�"OV1"c��8rPC�|����"O�}8t��( �b)�3�	�T�����"O�qrW���S+Ƒs6��Ƶi�"O�DH�eʳv����t��1}��9�"O�M3��[� �]��ޗ�@��"O.����ƅP\�(a��V>;����"O��Ӂ��o.�����P�.��a"O�x�҆ �`-��@?u~���"O)��X�<�>���O1c���"O©�B�(1C�҇���HlH*�"O� R��Y�'E�!�./ T"O2!���?4R�����@�Q̙S�"O��y�N /fJ��b�C�#sFe��"O��gHS!���	٤XZ>�!�"OxU:7iċm8Ūn�O?��0s"O�LSGM�Q��u:���Vޒ�3 "O�q�3�_8�X��*�M�$��"O�e�I�5^lK��<:�& �v"O@�!wjDh�#B�Y�J!�W"O�M�U��$Y������n{��[1"O(���ŀ�,�� ���gv4!�5"O�	 �슙z�`�3�5N���"Ox\h�F�o)*���A�N�qPV"O,!3㈁&��l��TS0����"O�Q�Ԃ/P��qe��]��T0D"O�I���c#��R���0]�"O��!y|����$C<I&���"O�H"��ԧA�Ct��[^� "OP�8S�Ȓh�� %�X�n�p��"OB�c6΅�Y�%j���7gh��"O��(V!�z���a�փX�ԉ�"O��;̐�|_@4j �!z<��"O��dD�[�������A�i�!"O���e$\�O�c���+uZh�g"O�E�r᚜G�XK�g݁kל�"O��3�O
�w�t}�!�۞��$� "O@��M�2z������y`�e�Q"O|H��V��ʐ� I>Y��"O���a��Y�ł�f�#*/  �"O��N.
�:aB���p��г�"OPˤ�9�8��U���	�� "O!��m�& R`���\'�^��3"O�B1��O�:�
��+O[^�r�"OB�[���xN���-IV��5"O���O cBP��׆�RC���7"O|��EH��'�4:,�7��cA"O�Xba*����)��?���"O��`A�#4�䅂d�8��T"O��K`������'v����"OrE�A�>.��@H���W߄�s�"OX�@+֯X	@F�6�v$��"O��9#�P$@�}b��ˮulfL�W"O^�ZЀ��-$�	i���,@�.��p"O����Ʋ	�Ā��nݧ��@!"O���ea�plDH�3�V����[�"O��墋-[+� �"Ob���G%b�°�L� O��b�"O� "��挍�!f��7�
/N���"Om0n���l�K�O�*�b�#p"O�� �
�"^X�	�΀"OD�`��KZ����D�z�r܋0"O���G�,o<ܡ�R�T�~��d"O�AT��w=X�1��]�Ƅ��"O4��eF¡QX��;RC)HU�1"O����#��ItR��8�t�"O`�E��A��`;��A@^Y�E"Oʝ�T�F�P6���jI_��"O��;�̓����a! 4T���7"O���T��l�RY�	�&V�A�"O&a�)O-**.Dj�HZ7*����"O~yAu%86���@�Ĳ�"O:$s3bH�
�*�I�o�ff�;q"O��c!n�:��C$�\�)aK�"ON�����l|��򀝋B�,���"O�R�*��P�����r����'"O,��#뀉fA�K@뗶*�8<h"O�i���b�
�1�IV9LۖP�v"O�a��M�`�>1H��Kٶ���"O^d�6�M�8�jp���\�<8z���"OR8�edK=k?@)� �]_,�\�"O8�(�L[���H�/D�v�"O��:�Q�{t�)VN�
oʑS "O^l�'�����Y0�S'X�E"O�E��̙�IU��l��n�U��"O�<���*y����E	RBҽ��"O,����X;Oc.,;`,�<E��f"O�l"5嚩2fb�ktI�	*t �"OQ�G��#o��pD�X�g���j�"Olp��E^���%�B���rE"O�Pم��	I�mӲ%�W����"O�aY���A>�����$��Ic"OL��G�K� v�C6bV"6c�`�b"O����"@䨳@E�SV@��"O�@IÃ�4E3��DiϾ.ߒ�A "O�,����~�z�r�Ƣq�ޅ*3"O2|ZwmҸq1�-ci�)V�ht[g"O@��+��_��,�Z���%�V"O��(CO�6�[��]�I���F"O�� �%$Zx����">����e"O�`xV�\�Sf�RE��O����r"O�$�G�U3Q���%h��_�*��w"O< �F��1�$���Q�D�s"O&� ���	��}cD�\�8 ����"O�����׽'�t��G�{�J(I7"O���6M9����a�D{�0��"O�*Ξx#���0 �,X`�-J�"O�@d(�:�
M�@o�~����q"OZl���R�@9\,`Gc� EBp� e"Oz̢�j�b�>�!�ǚr�:�5"O2��e�9=N�ڦ���p`Г"O�|��C��o��٫��@&�b��"O���g%5@x��U�Ӡ�h��D"OZq"[!D�f�pI�0����V"O�]Ag�׭ic��'��s��Y"O� ��\�Q��ts`��5�0�7"On����\.��'ցlЁ�"O�hwH�c�&�qH?R�Z;E"O��s�r�(��`b�Z�r�˗"O>)����3�6|i��طRo�|#F"O�l��.�
fD��T� �nT<0k2"OP��%�/��[���@HY8T"O� %r ��7\�dh�ŊU��퉇"OD r�ΰ%f��#�N�T�j1"OnH�
��NZ�����M�-b�a��"O�j��+=��玗�'�����#D�x����Լ���˷�|J3m'D��Q$ˍ�c��p�a�Vj- �8D����M4g�y��,C2*qp���6D��@,�.vq���ߩ.� ��k"D��I��GZ��7m�>�Ɓ���>D��a�E�{�2��4�3}l�I�B*2D� ��MY-t�"i�M���)�1D�8�֯��p�����H�j��ԛ�N.D��f� 9EҐ�Ӏ�3N�<��,D�4Ȥ-�;c��0#dI
G��Di�C*D��ɑ/��4LJp��&qh�&D�8�PJ .}��L �E;� �ˆ�?D��RUDC	>\���c�Hlĸ*�o>D�L�1���`�"|�s�ůN-��Jr�;D����C�,:J�A�N�]�H��-9D�,��� 3B����#�f����f8D���e��"|���c(����4D��l� w�)A0ATJr�rUk6D��ڤ���a���i'>f���.D�t�c��������W,���`ă"D�x�'(��u����3����=)v�!D���ª�0&�D�&��f����S2D�h���5�R��G�>Nn�8�%D��pg�׈!Hx����E�����	!D��RK[�]��:Tł�>�a�`,D���W�X%��a��A�#��$.D�D�R�P�^	���$ߡQ>�S�A6D����H�](Rar��ړG�2�@�1D��9��r�t��.8i/Ҥ�5kj��D{��	Є���Q�(	bN�+�ھ
!�D����j��V]�6x�5`�C!�<%ڰ����@=���#���!�dT��r�H�r
����L �!�V�/�}Q䄆=Z�^a��G�V�!�Ɉ&4>�Q.�L�TIk��1DJ!�D���"Tr&��=@Zs��@!�ď&q��-���Q� �9HwFֿOR!�0$���1!a���V�H��:5�$'�O|S��Ad��<d�F'=�L=�$"O���V'��e�,!b�'u$��D"O�؉�@�Dx��a`�x���',�I1%Zp��Ç`kH%�� 9N�dB�	#Z�90���1�$�H�i+ldB�ɱ7��ًf�]�v3���O̊j"
B�ɸX��i���C�?�R�Ï�~�HB䉝'F�I '�?��:&���bC�� Z��&k
!��䀡"�6/��B��;�ҍr�$��l��|p����K(zB��*V �1@X�������Tf�DB�"Kq� �Ӈ�-��fV�4>b����Okj0A���Xd�������$�Ff��ѥn��5ti��χxrp��Ni*�kd�QF �Ѕҫ'�B1��HW������_q�`�C�#iA2���U) �/�>�����i�b���jD���&D�L��"�c�����	m�	36��=�c�кp�}��$F�:��B�0a�W#ؽ8&t� �MD��B�+����1�\�/٪(��KY����7�"��p�ƫE�0�	3%TC�!�� (u�2Hۗ.�Z�J�	O�\$\1�"O4�a
�B1��I�g�ș�"O YX��R
:�
A��g:<���Kr�'�	���kF�PǋIO6��m*��<!��5|��:����#�[l�<�c�}��dA�'T�%�0R�ŋ`̓��=�k!
�eq���	,)x<���Y�<��nf��h��b��V�Y�<y���!w�$�AÉW�c84�a�d�j�<1j ܘyh�iX�*��)�Hh~"�D*ڧ{�rP�u@��6,RpP劭o;�ńȓ>�8ЋA	LDJ��B'D*wE��ȓ<$x�`�Ŝ>pK�.�$}D^�͓��?aqdI�h�
�`��pT\�{�C\[�<�m+r ��:q�ST�l㡍YX�<9��W�ŋ���OC΄����W�<Y$	��N���"õd�E) P�<����&�`񫏜t8iQ.ZL�<���oQ,ʰ��Uu�a��K���?1v �7hg\�y�Y�/��Q� ��hO?�I�)_�9��W1��P���	�X�HC�I�*Ѳ���"������C
��C䉜¢Ѷ�[�}Cf@��BkJ�C��:r,;��V�:�@|�r�ŴC�ɢG�\q�sF|Iz ������l74�l��I�7����Re���� ��T�<��g��r�0
л��MT�<�1I�/��@t)� j�	���O�<Ɂ��)��%�� �|�x�5m�f�<ٲm�y�bu����	�XX2��}�<٤+IA����CP�K]��Ùv�<�`R�e�U��CvvdX6� r�<s��!�����:��%X���v�<!7��&v=����I)
�x�3�u~B�)�'m�@��#-Ԙ3�]�uA�qt���!z���sď�i�l,2!%��|����A�Ե��ϼt���##��$Q�ȓ_�$�{R���5a!I�#���'tў"|���78��D+1�P�p�X�<QV���#�"����#C4����U_~�'D,KR��0n��]�6�B�dЎyR�'���.Lg�0��C�Z�p��_�|�C��6 �:��O�='�Ҽ�a	%9ijC�I);l�E9e�	zc�ȃ$A�<�rC�I�;
��e�4}o��kpk��uKLC䉦} �[ħ�$<����(D#<�,O��}�׏�)M&	�0k�TjT���<�㇝�>(�Rc���xxby	�u�<����m
�i���	Z.yˣ��y�<����S�lL�MU,\�;tFw�<�JP�~��H��Ȍ?.N8	�&/�j�<	�)]�}��L�&��U�d�'|�?��Ã�<ddh�O��\�p+0�D���B�>���FC�N&�`� /� #>��	��/��aXA`�y���	`I�_�!�Dǖ;�fX�ԡ�/�M�q�]8h�!�s������%4 �
0	�K�!�d�*6Ⱦ`��N�:k�N쳶�I�n�!�$L<!��FE�A��ȓi(+���D��×'`��3��=D��SH�y��F�I
V$1��G�E޼�t%���yRH�yTM�#fG>zV ���`��yB/օb�2����k��A��Ă��yRm���N��cH�i�,��I� �y
� 2�A��X�Y=:PS4mH�X]3�"O�0�#d�F|P�bɶyҭb&"O,��CD=}�h4I�A���P"O����)�Tp�G[%t���p�D6�Iy��%�f8��jڕ���#u�\-G(��\�d��Ch�;�^(#�L��a
i�ȓS�|��&뜱'�Uj��*�����nV�h���^�c�,��|?V9�ȓZ��9�JH�X��D�a�#h~]��q�|8�6HO�q����s�^:2��<�
�b��D��k�E�ށV گm���<)����WI��RPΛ�@�R$p��� ���O�,G{2�فOV�wdϴ4��FOS?�y� ��`4��5�2*]�,��A^!�y�"M�@����(�4%�H���*&�yr��-Q=d���b��!$Ƅ�e��y"X2W�j���i��|�k��y��Ⱦ��it�;���Bu���y�`0'A����5z�����yB��5L������wlP�K�Y3�yRKW�(!��"Q���W"�~f�i�'b���BEB�a�\�_�f�X��	�'��{�$S�c��Ca�&q?������O\�}"�oV�+�t�g�ȇ|��=WM�~�<��ޝ%g��ɵ��(m3ftF�w�<)��M����_$VJ���&�G�<1b�ʲ 8j�h0��)t��d���o�<Af�12�*Y1fH�Y%�!�eGi�<�sM��j^8�����?�~�C�o�g��\�'���Ct�	�R bM��T�{	�'*�������*)���|YN�I	�'[������+��E�W�rR&�����8x���P�Ӊ	EV������;P2�ȓXP�� p��%U��a��) �\���A	��w#F ��b�E�ȓ���� �Zɑ �M�����":�2�B�(S�h�ÁO.x7n �
�'��	�ѩ�����A��?�F9c�'�<��w�ܨ`"�xѠ ��qr��5<OH5r��B6������4���q4O��$ڰd��\��cD��n5���!�d�$���(u��*b�(�g��}�!�ĕJ��n̺���i
(gp�Z�"O,B����(����	ϥw|hXTI3�S��yb�({��  4��9P��cģ	�y�&E'���㬜�KN�8#�ܐ�y��i�P��]'������yr	���S`꟡.<����y��81#nĀԡ�+�$ѴN���y��;�n���Q�*��i��� �y�ܔ��ѻA�Ց��I�mA=�0<y����'���rC"��[Ѭ�&r�\��'�fqkiY�<+���i��ƕ)���[�ÔlÞzn�� �nڰW}��c��$9�H!�[R��e``�ɯnܽ����=�s�X��vq@r�Y�c`D��=`��W(�X��Um ����Ex��):���77д$�a/-S�Dp�[�'���Ӡ3yB�
�o09�䧓�A��C�ɤ�2DJg��%*�2�Ã .�rC�ɴ\�	kŤ�(Z�ȩ���ʹZ�O܈��*I��@A�ԘP"Ot�@ǜW�BLWJ	=Nu��"Ob��&���MH�ɘ�Oـ��� "O� xeǊ �kL�c�͔(�J	�"O>YPժ ]���Z1g�"f�Z"O�a�bo"*�b$q�)�B�� "O��)��W�#���FC�渹��"O�y5D� wϊx`�����Mjv"O�a�`$/`�H� n;���3�"O�AA�c���
�,+�M`�"OdJ��ęS���b�A�����'HўD5Q�)�`	B���s�[�*D�0�%
��&�](x�Y�&�)D��!Pm�F^�ɘ���?iޑz0`)D��i�Er�����عf�]��%D�T#�m��h�BR�#��p��#D�h�uʆ�<q:(r�ďd�f�(�("D���
��Z�44a��q�&��M>ⓛ?و�I��鹤���)>��`�F�
.�!�d�#�2`�anS�<�Öc��5o!�Dֺ�HF�F�R�^)Ӣ��"x<!��J=G�-�CZ�� 4�Q"�L�!���H�D�X_�^���BA�+�!�DR$,��EKXj<��_�V�!�D�9���0bpE��$�!-�a��'��m��a�?��0f�N  ��A�
�'P�ֆ�鴵��!Y-�2�K
�'^�r��+T/~)�jϣ3:����'�
m23�8FS�a�Т&��ي�'	ڬP5�D1������#�p���'z@�Q�Dô@ͤ���-�$U�@�'���qπ�E��a�DcĜ��4A�yB�'��$�a��>;�:��]8~e8`s	�'������&D�Gn��nqH��'JTEJ�\$X*��S0�(iB^��'��"���_�bH@�o�#f��(
�'�xɀP��iq�X���Ҳ�Jlc	�'>�\���ȩQ��	q� +�,� ��)��<�P�Q�@�,m�`���0�.�#��^5�hO?�??( ���})�pAdەzTnC��L��� 6��s@�L�RŘ�Ĕ��)�dX+gCҥ��$��0I0 ÐI.;�H�=E��'�F��EK�c�x"ꎺG�����'e��;��ЛF�5!�I;�� C�'�%�Q��@� �3�f$cl����'�p����:M�d(�/\�@{eO����?jx���(�M�j��"O�#�:p�Ƅ��H�U�8ٳt"O�����[>na�C���}M��y�"O�PaW��pR�0�Ә-dVM�7"O8�ADߎ!7j���D��b��Rg"O}����vS|���#ӻM��i)%"OL��1oƚg�P8Q���*�P��"O���o�>Mk��cC��� (���"O�D#5LN�WMZ�PV�.@��1�"�S��yb��>+w0�#�$G�e h�(�&O&�y�Վ/#�Ĉc��#� �3m؟�y��<=x<i�w"���l�R�W5�y"��"U�����L��x�
�y�_�y��ؤ`���*ӏ@	v������y��H��(��
�g�h����y�eq�ar�F�~�C��P��O
�=�Os��*T�O4vWֹ!qLѤxD�Y�'�ў"~��Ҙ�=�	)�V�]�JŨ�"O��#4! )EL��3��aB�tV"O�ػ�u8&4٧g[-\�Лp"O��$F� �z�&h
�gJ����"O� �)��B�{G4��E���1�4�"OYK�F�8�T�1�B�x�q��'�O�je�ѝ�nM�$����ʔ"O��BQmGyHx�eЯQ��yE"O��9`l��
�����'����"O���v��8GR���C�=`��X���'4�O��S��ĘcL�с�bL�t�RD2A"O��I/J�\xy�B�2��@rT"O`Yp"J/�T�+o�<�>�b�"O������NU�}�m�*|ui�"O&Q3���vbL�F�#z��5�v"O��pG�,$��{�JT�}�Fl"O��BVLЛc���� D�A�""O��`@��10���r�֒p��t��"ON@1T��9.�0�Ŋpj�P�"O�m��`ݘ����]?P�Ak�"O�����'r�h�"ػW���0�9O�����E6����N�a"����I)j�!��K�|�B	!��ܿ�H�̅*D!��V]������4�KS�a~�R��R2�B6j�V8q2�6J�EIs�4D��R��"E	���-tΞ q�E6D��P�%)@lH@�c��"�\���C������G�	�hc�K�X9ҭ�%���!���K$�� !Sw+R�ɑd(�!��D~�hSp�Rč��"�(�!�D�u,H�Tn�/�d�4k��/ !�dR5@���`	.ŏ��*[�C!��]���jB��2�(Ӊ�Q!�Ă�_}�LP%�7Q�1C��N:���)�S�OE���G��(U�]B��%Cͳ�O��=E�T�Ɯ)j�X0��B^��YR-Î�y�
�dm�&%
��k�㈨�y�9�Ȕ�dcM�z֍)��ٔ�0=��(�~�Y9��9x�@�3�F���y��)>c����Ł�p�-��h_��y�&M�S
	�s(D=f��r�+� �y"�ݤ�p��3a�2�|驖���y2c�`���V*з#�&y�� ��y�"O�d���X���tC��߼�yB-��<4S��(OZ��O�:�Oڣ?���Т��V=/Kp���ª#)r��ȓ~�NAPd2&��
[�J�~Ԇȓ!��x2�Q�]��M��ዉb.4E|B��'ҀbP�@����ϕ�nƖB�ɀ�>ěE.ĥb����b�I�2TDB�#x��`�N�?��L�!�D);�DB�	);�l�i�A�[�>��UcA@~t����<I0�*aYB���+�6�s�If�<��O�'���ʕG�4B��Rg�<)�Z'U|9!VC��fAb���d�<	ʎ�e>4	���u�<��C!�^�'X�yM�Gh)��+�0���V<�y���s�|I���w� �� ��yҍ�o㠸�0�Lz�r�AVi�&�yҨ��@��-��k#t��En��y2 ��`��M��o�`��s-�yrΗo}H0��;m)xe�kS��yBlß?p8������*�B2�yB�ƴR=C�'1+nt	����yҭJ�BW4fB� ��5�'N/�yRl�o����2l��R�$8�
A�x"�'�E��ꉘFW$�H$��j�2��'k^-���G�4d֘ɒ)�`@��X	��� &l��٩h�&xK$
��s�H9��"O$%� �Q�&0�Gɒ�GG����"OH�"f�4h��a��O+� 	�"O��ծ��x�D�ztG��L�l���"O ���C0&��}0f	s�4�"O���w+�J����5Z���+T"O��JT�7��s�̋a�Xh"O�4�s�[�;K"|Q��ڡ-���e"O
H����b1��.\���M��"OZm�GϱX�jL��-�-qw,-Cb"O�h�(��AШ E��`E�8�"O��Z�R���r�=k#xS�'��g�Sp�xBE͔mt����lC�I�7�Թ�f�����u����G[6C�I /�0��@L_�8f����6x: ��&�O�
�(La�xD��/��X���t�B٢9�� (1*S�z�,�����Pv�� 7��P�Ďxh����u��a�+Ů})��g	L(�ȓlX`i�P
�T�L�� �+�\��'�ў"|�U*�U��p���t��m��$�i�<	��������K7�r���Ol�<!vfB>Xf��)��$�`�Xj�<���B9��H�0��pU��l�<�nL$:�Xu��%��sBI�k�<	�j��sߌ����e�\q{ /�i�<�H�/�P�XW�V�m?0����e�<Q�*6w�>-��P�Q�x`�2oBU�<i�-\f����+��F��k�<��f�O�Ɓ�e%ި0Jl�0Q�Ai�<aE�'-����ˆ����R*�g�<�6��N�2���@n2��I�d�<��l^Ȣ�kJW2e����c��,�?iaa�%{+>9X�^]��+5�]�<Q��5u��M� �Ɖ0 ��䫅X�<����0�
%�<8���`P�<�Gu�@����J#L�M�<�p���X`�G�8�<�gRb�<�$�ҡ6Gt�뇤{9v� s�<��!׼Yb��0@���>�x�
�Y��?���?y�MU�jE��}*�8�+?���?���TXҠ�0!Ünn\0C��O�<��"� J�I�g�
b�Pՠ�B�<i�F�")0,� �	K�4xs��}�<qR	Q�^��Xq5o�^Ĕ�����z�<iE�R�Q����e�#�18G�q�<i5�S�Ig��(�J
�Y"��p��b�<��#G0r `���0F}H8�a�^�<1 H�F���9pDð�f���e�<y3�@��B$
�m��I��! ��_�<!�,�0����@ކ8j��ctIQ�<�G
�]	�%��A�>Y��+1.BO�<a�j�?1s�۴�<u�(��N�P�<Ag�9>n�9ҧ$�X.t�E�QU�<��k��N|�%� 'R1:$�"c��L�<��^��Yɷ((��P��\�<q�j�6?�~x�'A*.��(#��Y�<�2.FAzLA2�(	i�X�<��o�`~���7��� ��qV�i�<��kN�	��ȹ�U�X�&�@cLHi�<7�ֵ�(�I#`H���`� �z�<I����i�"�fɜ�5�ep���r�<1��� E����3��5��j�u�<�c ��^(��fɕx��l �/�s�<� ��Zա�R��pp���6X�ƭ�"O����F�&h�hC���L!�"OP-�P�.��̹#�Mp�|ZP"O;p�S�C*�)tK(Hq��;!"O���r��a��Z )Y8{�xx�@"ONDv�9?�ndFH�D49����D{��)�OQ��a�٘5B�h#�Y5!�䅎n��P�U-�S.Д�f��(3�	Gx�ܚ`F�4]�td�B������9D��y�	��WZ	{sɟ�W��y�K7D���!ҋ3��{7��&�Q��O5D�H���љ2H����f���8D�,�Ƥ�,J��IV�ք%�~qRk6Ọ=�#DI��(� I*7[hmЁ�O�<�� ��jD&dP4��K��p'�O�<9��Ʀ%\�"�I��`?�U(�k�M�<AU-ڝ&�J���g�(KpP@P�F�<Q�KSP8����B�,�����G�<����U#�ec�������CNWy�<�fO�%B��t�])bD*�`rƎM�<I�
�d�~�����2�����KJ�<q��"O�t���R_d9XDn�<نkѿjZEy$��,.��� �^�<���.3���ʢ�X��.�sRaA@�<�b�ХlA�Œ��2H��i�y�<Q0⊜��Y�C�J�Ĥ`�Bt�<A� U�p�,P�4����c�V�<�¬B�*�87gʋ't��"�O�<1���MBn=f0|�Qa#I�'$�y2���8{A��E>��Z��yB���G��=��^Ej����I�y"�\�!\+�װL(�0�b�:>@C��y�L�	'/��u@>-�h�?J�:C��/(N5֖'�i��O�+�"c�pE{��4��./En�{�G�89��`��#��yB];IzN9a.g��h�Yȼh�'�x�v$�C)��\F�'[
���Oq~&lW+�_�DK�'l ��P	\�����W�a��L��'9�а����b���0 �_`zp��'��2ţߑz��P@g&�K`ɠ�'. Q���_b��a7e�I�r��ʓ P�Ʉ�/[Ȥ��^�;e��Gx��'P�����"xC��xfG�'(�4]`�'� %y�᝴�>$��LK�R��h�'�	A���"�H���D�
�����'�F�QG�N'U��d"��? S�y��'�|]�cBYN�F-UƖ����!�'8�5�[U:v��
*%�5�&&*D�P����p�b �uVl�y�*��A���r��n
(��� 7a�d�C�F#D��"����#\Hˡh�f[,���?D�HAtcЫ@)b��K�4�h�ʦ�;D�L1�f�U����{,Xر�4�OX�O���@�5|@����I�"�!�"Ol$3� ����wO��w"Ol 1�EQ�i�����]�E"O�,:�O�#�X��@CQ8���K�"O
�ơY�w��$��DD�Rc����"O�Zp)��4�<��e�r4"0�"O�M�Ҫ�4e�9���G�-����@74�0��ϋ�;���1��% �C��uh<�� �#�<Jfǽ#J��K�Ph�<���~�D
Q!	�*�a�c�<� �l���= �����%B��"Oʭ��#С9��A�0X{RAC�"OV�_��=k�AW�V��y�R"O��Cu&J9k�"X�e�QH� 1����D{��键+�5�c%�=�Z,;���y�!�d�#U�%����}�u�e�A5!��D6H�Bi	�D����F�~'!�C4��T�����@σ�Z#!���M1���.�
K�x𢧨Q8np!�$�/e�ΰx"���6���!��)Y!��,oY����	��ؚ���7L�d+�S�O�e��O��^�`���#b5Љy��'8�yc�bX�UF,0���_�e�!�	�'�h�2�D�~�9i��H�\�`�'�B�ŧ}�`�:ǂX,e�F]c�JT5�yr��"*B�0��S^A����҉�yBoM�/�py����L� iK "X��yB,�B������R�	+��y���|ṳ��v&y�Am����'o�{��J�U)�����L�ha'	:�y�'�7Eɚ���D�zInm��S��yȀ�zo�d�3L��z�F�I����yB߱5V=U�<nY:YӔ.���y�흛1��ݫ���azVe;��>�yr�)�m�J����b�*l���p�D �<�ߓaV�z5^�3��Q�n_$Q� ���w�ؤ�&A��T�����c��І�E�^8�b^�_\�h@��ְ6]V|�ȓ�(��%Ɠ<W:(�{a��!ƴ��I>�-Q4N�3)!�%�R�ɇ�u���b�H�0P!�`�&���ȓt�"�ҥ�c�H�`e[8�|��IBf�(F(ϻu�"��2*Ÿe댝ϓ��#|O�mH
�':���#�@�{�BH �"O$�����:�ɥ�%���v"O
I��$��Hz�t�D�\xa�"OB`q@F_��R`�Í��zD��"O�Y���#&�a�'HX'1�����"O�	@WGL	�ꅈi=BT��a�"O.���ŵ)2T̹�H��2Hl���%�O���+&����ĨJf��)ɱT�!��l�(-���=���DF��O�!��ًW�T�q�ʍ�2�v5#�D���!��?sB4�B��Е1�<��d�*�!�䜝K�!(�+�@��D����=E��'��z��5�R���$H!!_T�'2�E�Ë*��@��"BE�a�
�'%���"�I�:�U��AQ<,(]�	�'<\O��[���21�"6^^L2�'��5S����?�N�s3�<1�Bs�'���i�L�))����l��Z���'�D����	*��1�0oM�f�1`�'.<j���I�^`�!]$����'x&uR��äx7zԧ�R�2�`�'Ͳ�+LO�T��4E��I�'���H%g�2JЩ��O����
�'v6�폔0�: !�d
�J��
�'9��K���2
4@��X�6�J
�'P�X��r�>���MNl&��	�'�
�����9�"����D�G�r�S�'e�زVV���Pg��i[��C�'�LU��苴
�8ࢎ�_P I �OZ[�ߎ2B}�6 R�.����"O�嘄�)2l�FO�n;���"O� R|��@�*��2�Њ)N��"O`�Yc!���9���P���$�B"O��
��S @��������V����"O�D�х�?f�kC�ϑ��D�1"Op��&/F�Ǎ*����,�C�*D����ͣPER�Y%R�E;V���`4D�H���/EL���A���.d(��' D�C��!V3()&A�"�����?D�|s��R�5�e�Ę�D
�e���{��E{���7��e�����V��%�!���$5.8�eB��
!��Ȇ�:�!�d��jD�Pr���J�ҧ(O�o�!�$_>|��iH����>�ौ&,�!�d[����ǘe��L�R�J%X!�$�sYe1�툥~�� O��3i!�N��pɸq.�PtD����<m!��[3!ㄠ�Wk��1U\i�
A_g!�F�bV̹�X)&�jPA'G���ȓ�c�ҡ{�lA:��I;)g�X�ȓ �D11� ̂�,d�B���
:���ȓ��-:`��S�b�b�,\&C�����.�C�Ï?2���@��8c2���P�|�N�(���q�"S����ȓ:�d�! p���3�;D����ȓC^QQb ��>��p�ӯT�>݄�`Q^���K�~#�p���.w$�ȓ\����X�V�����C�E�x��ȓ) ���b��*p9sIG��1�ȓQD�l��B���,�$ ��`��ȓf}�\���f�0Q I�D� �ȓ��u���!Q��
�&2f��sV� TM4��%��	S/`�^U�ȓs%���̇ ,p�E�d�p8`��f:�e��o�lȵL�_���ȓ4���k1nĈE��Cܓc����ȓc�=����E�]K7o-� <��H`b��әz 3p�	Tp$��R�=J�,�<=����l����ȓJ�z��Y�&Z5�	%�ƕ�ȓ0�nxJPfG�)�4˖�!e��̅ȓP����=+��D)0�O#(< y�ȓQ캨�u��%�t�S��$Ćͅ�YL����׽c �#�/C��u�ȓ~"d�T!y��$�׶H\)����q�,M��d��7�lh������N"��X��@\�!dp ��2\��j�y.9�-� u۔݇ȓ�jp��g�
&�j%��'��$X���-  ���ŗYIz��ĂZ<J4�|��=�}���)E	xR$�$��|�ȓ�� ��\�t��TF˽N����l�X���dD��;���t����}x`���+O�6٧�"'� ��ȓ]zQ@p&�{f9!����'�0$�ȓx��u�֣�
	��%�-��	��9��Y����2Il�e�;X�-�ȓR+���$U�=� �3a��>������ d�D 0#o�2��B�/vQ��{I��9U�V�?�j�A)����ȓxE�=r)�==Y�p���~{B]�����Z�$צ :�q�$�Ռ)�^��ȓIk !�6�D�}܎UH���N{V��gf���;;��в��S����ȓu	$,�(��D(�}�'�@�Bx��S�? ��7Eۗu%z��w�B�jH`��"O�`�E�-F��T�%��}eD��#"O� ��03��8i�*[�8�Q(�"O�����!$��(֫�x�X��"O������-t���� ]F�0"O<PA��[�TTc�P�(���3'"O����EŒ���j�(�d`�"O^�bf�L� 8�`dJ&$���+�"O&���.��Ye�F/��"�)�Y�!���L
����/:��3I8�!��� ���SB�8l�RAJ4K|z!�ˣ��cc�G�D�n����?@]!��Y�Z�� �(v�����CF�i!�B� �����CX�t�H|)�%_U!�dH	u���I������\0IA!�S*z"M�4�L�FH���o��:!�dM�E�б�q�J��|����d)!�өx�|�	��0��%G��Z'!��8i�R2�����3}$!�䌃&Dԍ
�-ϭe||�s���f!��$%�N�F,�"(^�eچ_�>s!��9oȵ�w��h�S�
,�!��<�Z���EM�J�� ]�;�!�ʂ$GD$K�"r����� �!�䇎S������=��GΆc�!���	��ܻ�d��=��t����!��\�:��В�+^�)D�QǖAx!��F��p����l����u!�O�Ȉ�c��7�8��B�bj!�ϋB���y�"t��욣�ƌ9j!�<h� Y�'�{�*�I�� &~Q!�.w��a��Y }�̨Ǌ�W�!��ɟc7�]1��
�NE���N�!��%�1��V�� =��_�>�!���9��ȁBΗ�(�^0õ��pf!�d�N ��t�Bw�����RG!�D��D~R�e(��t1��P�@�!��P�h�%��P�}P� z�!��M���K�%99Դ�b@HP�!�$%F~����#�|�YC@�-q!��2<����*'j/A!���&8!�D�F'���s �1"�����f!�$	�d9�5�PЛPd���ۖ\�!�d͚L��t��K�&ML�\ ���T�!��S�>38�� �
)4����[/V�!��Rj������4�����KM�]!�D�ZB�
�)�@�z����C�ms!���L`\�*7D@n��c�랍=h!��B D�� .%�8�0�I5_U!��^<C��'� d�Z�[RF���!�28�nIr"�L;G/4�Z���!�dY�@�qK�ɛ�|..�c��P��!�?"�A�*@q�ub��n�!�D�ap�
%ұ
B�'��:!�ē;��K��"oxe�SlDa�!�D�j�h�jw���k�~Xm-4&�!�D� U̼�X��OV=�*W!T�!�߅4n��˒ bmq��̢E�!�d��4��<��@�N�#/�!�$Q�`!�����Ƭ9���J6s!�D�8��u!��J֒�H��K�)l!�dT�K�V(��2���S�jD*%;!�$��I1G`� G���# �j!�D¡;:D &M���*�bL_�A!�� FMjTl�H?b���EҎp��*D"O����!t�p���S�N���Q�"Opi �꘳3/��E�("�;p"O�Y0�=+#�J�O�Sޜ)�"OЉ�t�!@��ʶ�Ԕkz�S�"O��!��'�>P1�r+h�i"O�0�t�H�>� �w��.d�(�"O�1`Fi���o�u�@�7"O����O]�E!�!�w��;b[�{�"O��S�`�/��ec�O�TF��Z�"Oxt����Pw| ���+26r���"O�i�G�Y�1_�#�H?g�r�"�"O���ehQ��)pA_��c�"O��8 �K�Y2�QH���`�@|�"O@���w�0hy��6hp���"O���J����휻~��b"O����F�2us��R�(�Z���"O�Y��ɐ�H��}�%&��!׎u��"Ovu�2�����5�Z*��H�u"O�!� Q�=P���T1N�� �"O�8p�lI���5�d��tE.S"O� $��4����;����"O��t΀F��z��*&}��"O�A�g�
Z˞�Ё��+9�>(�e"O���Մ�IjeC�����7!�dJ�7���	�
���чY�)�!��)]c�4:��7i�J�ʇML;"&!�$�
T{Q� c�O�xQ0�#�!�+���2�f�$��iի^Hh!�Ĕ�Q<<�8T��L���O�,b!��ѨB��8���Y-N�<)�����!���Sҙ�n���!����Z�!��7Q�>����=n��;A�]��!򄜔s�% �`� ��a�D"�5�!򤕯[p�RRGY�^�B1�ASr�!�d��[�Э�!��V�5�>G�!�G�7~X��@C���h��&R)e�!�d�s���H��\�F���!��S<!�dB��*�[4��R��D��>9
!�d)1nX���'�*"��%K�-ӛr#!�V�Vƾq9��5Ts4-^�D8��'�Ġ(6�X2@����S���? �a�'�*�i!ыD*�(��z�*t��'uvdY�5a�Ty�Q�&����'���"��F�}_�i�Ç� "�Zr�'s�����;����N���#
�'�(���W�X��R��K���
�'�|�q#��ma��Ц�C�.���1
�'�ʜ�SK�`/��V�G0$6�s�'�v�)�DN9gE������[�'�Bl�N�	5X�Cv���#����'�J�J��$Q��yFJ4��P�'�<����ԙZ�t�h5Jȣ0?D|#�'�p�k�SU%���W&	!0d���'��A �P�_=���+��D�'�ruҥV$�jH�a��2�\��
�' yh��~�����4%����	�'��5�#�'�уS%P� ��k	�'�RY���W�4� �K��ڊA��'H�$�G_�N�.Ra��:>ے��'e� s��:+Ֆ�Q.׈0�`�a�'tx=�Ď�Pu�E�)����'[2�[��y�� ��!��(�ح
�'����G��BoJ3W!�'�ָ�y
�  ��WI��J��7/�n�9�b"O�J�:���e�E�^�6��'"O2�R�BN���#gS�'�}��"Oh��".�Q��9"�аM��<�"O��##�*m���a�l�5v���g"O:q���^�)[�mp��4bE{�"O��D� 7�v���~�D�0�"OJ���ȁ�%6��m�l*�p"O��k��s��q��N#g�8�	"O&�£�u��9���u�	�"O �	#*�9�U�W+N��̐�"Onys�ᗍ���#$�W�3��-؀"O�ȴ�A�-F��u�R�b�+�"O�h�6h����c��� ���"O}���̘G��Z Ǐ f��Հ�"Ot���]z��"F��'Ԭ�Jt"O1�E�Ս !����B�"Ӵ��@"O,�@⊶{�J@���A�h`�4"O����Q?,�\}�'�LB�5!B"O��È6]�I�A�S�aA�L٦"O>a;��#�$DV6rm"q"O@ܳ��dR��p��A&��"O��GS	-ح�ŊZ��"�U"O����i��%�T�Jt��5���yBNЯt��I��Y�<�xJ��L��y�&^y��3�..%	�aD�_��y�	�<X;��(5/�q��yb@׀=p-+���cY�a�B'2�yr�E����g�D�욗�y��r���XS3�(��F��y��C�v��yWEGO:V�a�� !�yR� �X[�g����a�$
��y2��$2$�:��"��4��̉�y"Ҫwf��W�Z�N������yr�Ճ*<(-���3
4�i��T��yR��F����b�4R'�d�^5�yh�A{Q"R���rR��6�y���sD@����8�����NA��y�,E�=����`�	k��j�EV��y�F� ���1FK�+�!��-0�y�o]F� �!+*�a[�&C��y��W;e)��Ц%�w�]��%°�y�	ms�8Kt�؟u
�� ��F��y2F$����0CBn�\��B�<�y��ïR��y�$�5�������y��E�Ȁ��2,D��; N.�y���p����OL+0ݘm���\!�y"@�H�����ֆ+:Z�����yR��-I��-�򡘥u	����A���y�S�T-h��b��m����y2�)
���j�X��#�.T$�y�H�;v�|a�L��]`V�+V�F��yB��!-��U��Wc��v��y�J�{��x�Q��V��$B� 8�yb$\�M��� l\Ht*�U�'�y�LE�n�|��u��BkdA�jٮ�y�n�dJ����
:��}�"��y�F�
r�4��eA�8^vAʑk7�y��x�rU3%�9��1����-�y�O�D�D(�ˑ6@c&�y2#)��\�UeǓ���	t%�*�y�+�r�٣� �>s��mA#!���y�(�vY�p�A]�x���e�R��y�aăn�Й����x�9�*�y
� (�4�<ǂ�"��� ����"O�A��_�I�R��4��l�5
q"On��C�Px%Xͻ�N�<U�B��"O�0��̌
%���PM�;���Q"O
��4lӯt�N=:�AE/�P�8�"O�X�0��:7|�`�J��`�~��D"Oz�h0�̷Xe�����6�X\(!"O�щ��As�@����Z���"Oȵȓ^Z�.�0��d��t"O�Yɠ�Ƨg�lU�Wfڏ�H�Qt"Oz ���(ܢ���E"�����"O 1�`F[W�N8[ň��n��T"Ohk���/h���:�f�=�,T��"O���ոV(���䈮�j�"O$=Kp�Ɩ0x�+0$�5$�d=qF"O��D�W�4���[�!q�p"O^+���*� -s̙.8���"O��pWL� `�0y�`�ւ'�"4"S"O���e&I�%^ݑ��ތ<z�$��"OBe���S�^�v�EO�7� c"O�)��M V����.]�F�mkE"OA;a#�5f8S�G�l��	�3"O�Ό�f�ᰣ�
��\	%"O����a�(*Ť"�H�����d"O���a 8+�h+7���W�b3�"O���M'tP��b:9U* �`"O�8���N�#�v��t�@�#E��"O"�i�J�B�RvMK�X:ҽ� "O4�d-3O���D�37���"O�M��#/�8�*&BE%r��"O�8�#(��^ �<�waM�g�FT��"O|X�ׯ �M��!���q0y!V"O���ߖ[u��H"MĶ3"Z|��"O� �B�kK�Eا�2;"d�A"Oؔ�vo���,��
�4<���b"O�Y�Ɔ�E�j���?k�)҆"O��� Ƒ&o���BQ�P�J�F��3"OTX�r�&2q��򫓢q)60�"O��p����:XBA�1K��>T���"O��q� �S���Z��!�"O���L)+���#!ɒ��]�"O4 1��Ŷsc0\�  �4�nA�Q"O����"	>��2@�F�8�{2"O���ՠ^!�\���˟!��l��"Onp"P�T�Fv<:�+G8<���"O�Hy2��-j~�`(�A	c#
�"OnRՠ��.l�	�UCG0E��I�$"O��b쟓9BM2h��C�洡�"O,��L/ggԉ����,T�,pqr"O�Ű�����"VƝ#Jܜ��"O��Ӧ��Vd��UV�8�!�"O�(�Q	6y�ph��ī#ֆ�"O��P��"�ti�R�  �X��"Ol	�㍓7�<�0�cƥ*�LM�"O쐩�H_(%� �%�(OJ9"OU��E(쨁��^�H"OHiq5eaG� �����[q<pr�"O>�co4Jx�-JoT�5"O�ebg���v�����kYD�j�"O�����+Y�&	�ցڛY�tK�"OH�c1K�c�.�kQ I�q�� ��"O�hx�`"u��僥�0�[�"O"!��G�R��Q������p��"O����Cܞ��GD��wC�Ih�"O� 6��`��� e�t��#O�,?�T"O��CH��}��A #���2��"O�=�$
�9,@�"ˠZ�\51P"O�� �"	6g(ȉP,p���b"O��#R+[�@��MP2��s�b�(6"O�p���{}���W�
�(8��t"O�Ĳ��=""����ݏ��A�"O*��L^8&v��FX�Z��÷"O.e�eI���B���^�8���"O��Ag��{�zA��d�Dy��p"O�l*�B�d$F!�Bݨ0v�us%"O.i�6��(ty�o��qH��v"O��`E��x{�O�*K�]"OR� `3_jЕ�(O.!�i�"O
�;���\ȃ0a01�"O��Q���k���y�R� �"Oԝx$���d���4�Js�<�J%"O֙�pCX]�N��'%�]�`�#�"O�1R�
�`�p�L�`?Zh��"O<Qc���>& �e�
;@+�BV"OZ`��,G�@�@���G�](���U"O��I��R�,��+�㒔*/60i�"O��rf냘E���ѳÁ6�(�d"O,z��N�G�P ;�d�$}b2=�"O��`�钱{�:�'� _.,H�"O���H
1㊁��*ѦR�"O�I������3I\Ki d9�"O�(q0�5\��#(�"%�:���"Ot9hՁ@�@[��Ai�z��F"O�!���ȓǜ�{����"O��w.I&� )xCdΆ�XQ��"O�]�7�F�@!�3��ʃ|�
�a�"O&o��J�H��A�}��a�"O�p����9[��qh�Ϛ���yrH�&�p �D
jf��bhЪ�y�m�7.< <�լH*i�*A��ƚ�y�a_w�0JP�LZ�D%$�ʓ�y��9��<�2/#(y^��DA��y�S;\��y�ѫ2<��Ѷ�=�yb\�q]�\;'	�/y��˵L���yBN�JV@����nE�p�����yR��A���s��5�Z�*���y�*@�A��倀��^�ya�����y��+���Y�+�<[�6������yrg������*ժG��jWd���y�˗�b��4���F��0�&/�<�yr��i>�9zr,EDQ$��l̘�y��N���	�ADk�2�[��P��y��
���ei\f���Ĕ�y���<��9*��^������"�y"bC�)֨��f`.h^v�X6�Q��y2-J�l�����s|�%K
�y���E���b�lѦ��K����yB�̫]�����*W�8���jŲ�y"�̒n�NQ�$�1|�f]c���yR�C{(tp�Ęo�����8�ye��|5�GHBz�S"h���yR��)測����R�r�`\%�y����	����Z�2�X���-�y��1�:�cՃè��%��oT�yR�zߘ���K ����s�J��yJ�M��m���$�l�HcE���y&Y���╧߱~�XPC�,Ư�yB�/���`��ֱE#6L�b��y
� R]!�FG�<�LEa�Q�F�q"O����!��3ȩ
�*wDFY��"O��PBS�fo(�I펢^���A"O��;D�	=�� ����#kD���Q"O�e	W�݅l����3����"O*A�v��� ���zwaDZ����"O�hňԩZ9"X�C�·l��})D"Oc0��
���9P�7Cv�H��"Oh�t��]ZN 	��?_�b$"O$�8D�E{pJ!��呍\^�TD"OX���0 U�wn��)n�ys�"O�\��C�N�xL��.Wԝ�C"O,�`b���{�ȓ�D�P�5�"O�-A��E�6I��f>.<(���"OnTn��I��P��h0JF�"O�1�ìYU����G� e�b"O~�"m!�(}��4����W"O~�!6�+�)ao�.M��=��"O<��ʹ,�H����> !��"O�邇��</����-Oj��"O��0f@̨ �h����`xI�R"O���lK&��I��E+a�Պ�Z���ɹe��R�6�oG�d��<��T>}�p`K
+伋 �F-dbly��8D����G�0T0�HR�A7VS0�P ���hO?���0R�����6N]<J����!���3|a֡��BX
lRg�$#0��V�������^gX �4n��]X��Rs�#D��e阥��Փ{6�H46�訟�Mh�����+�	��f���H�"O�����]f�xS�Z�~�]��V�0G{��O��dc�( �^D��6cg!�?�z�+��QlV�s�O�4[!��.kg���!��g�=2u���!���O�i�V͆ )M�ƅ��H��x{AO�j��ۗE�����eG�vN���n�<) K�O��(��u۱�W�?�t���ҩsD.���'�����Y�h�&�	¯{�x�aU.-�I8˰=YD���/o��:U&�zJ!H�e�W<��v��\9��ώ;_V�[�(�<+-�̓��?�W���a�f �}ռ��Pp�<�3D��{��E�dh�0;H�K�+�r�<�Cաk�@�� eM�g[�e���yyB�'8��� �=N (05�+YiR�ю�$2�l{P�:���'+��#�fM/s(��<�	��t��b��$Z�(�aL�+s&h�'�ў�>���9�N ���5E"z�N�G� B�	
5��pp �F7Sh0��̖rEB�	9f����]�VD���Ҿ1M�?A��o���}�"�,4	LU��K�
K49�BVN�<�$��D<@�G�0���C�r�<a�KΘ6��iSFO�5�Н	��NW�<y�gI�h�Cd�)5����#��T�<I��T��8���ݣlf���q�R�<Y��ӳ(0'��"-i���-]R�<1�Nݼ${^��hJ#|�]�!l�J<i��H�bM�p�F(8$�AI�+A%�)�ȓvI�`As�i]��⌅�-��Є�IG�'��X��fՆM5�=�tf�E ,dx	�'**��g�"K�4�-���%��'rў�}r���Q�tm��/Cݎ�cb"��<ɔ�џ&��`��e��]����QP�'��y�*N(0�4*�B�M�\� �!D�d	R��l~q�R�=�n�#V�>D�� �=1�,<4���#ь�3e�8��OV1�B��/w�Z�G^$.m��GV_�<)�4��ؓT!Ѡl��{"GR`�wܓ��<��K>9�<�Qf	�B�P�ԭMR؟��+4d���&0��)䋄�a�T��'@8Dy�D.�1O�P��N@��y�ֆ�Zl4I0��;���� ��/wrz��2 �^o)Jb�$3|O^����?N6��D�@�{~����'p�6MD^(�-Ȓ�� \S*U�L?Ul �	M��h�(e�U�'zL�$@цL(8$�ű"�'
�#=��Lq�Ȭ	t,���^Ѻ&�у��x����ho �˃ ��7�ڐb�K���	\�'s���P�F�y�j�� ��G�F�js"O�Ԉ3�Wnf}�T�@�]a��z`��@� �'b��e�3%�h���J,� ��2g��I���a����:pQ�A��j��B�	�}���rLNM>x���-��">ю�)���A�D�n��Y3!֩\Z!�d �2tn�ؓƇ~ݺ2&![c>�O��=���1�%	S�U��yд-E�Yl��"�I~�OY�a�.T��0��M�+����	�''� �C�2n�ޙ�c��{���z
�'��|�G*I�{�&���kHB�Ri�FOj� ��'Q��E��F�����'�ў�k@AƻfعHc%�uTq�:D�H��`�{�f�IA�%V�� ��7?�����0_,yc6L�:GeLA�f<'�C䉿�n�p��GL���1J���C�	-6uN��H��i�����\�t��d?��@2�3Q

q"fu��†e�C�	�"��L0(H,�7��v��C�	$5���x�EVn,A��jY�]�nC�	"S�&	rƆ=�Jݪ�DݳNC:!j����O� ��NG+!
�iӧHG�Z�J
�'>0�U�	N����#^ 4���'g��Pc		k$���OհM��%1�'�$��ā۷O��]j�ɮq�@u`�'��qA� �
l�P�`0	�/e�~��'ڂ�jd'ơt��U9P/�V��P��'�}0�kM��:�bOF�	�ON�=E��LW<T�l����e)�u1$/U(�y�/h�x����2b��`sf�y��V�HfN᪦‐NStPC�a�
�y�B��	�6�⠦J">� p���5�y!A�G�Tu��K8g��;w�A��ybF� �5�� Ybg��Wܓ�?1�'QΈ��WK�VF(p�̊H�G{Zw�1O�z�ꄣ��c� ޼0r���V"O��P��==���d�Q Y�ıh@"O��rd��8!=Z �ؠ&��( Q"O>�Kq	�c�X�p'���)Z"Od0��>Kb����X/&��"O^%�򂐥`� ��qDˌx�S"O6qx��\5i`F�b�0
���:�'s�OJ ��n_�6�Ƅ�� ��p\94"O��2@*���L����;{$��t�D2�S�(��� GƂ�#00DF��o�C�ɊA�6E�"�ٗ�Ī���$W̪C�	4�ZɋuE�)i��^BZ�C�I�`Q�!P�ƍD���K�C۵k�B�ɋ<]��{���ԃ�^���c���'��'��O�5��n]�A�B�JB%M�h�\ ���?�}r��@���B_r}t艄+�~��)ڧ cLY�͓jc��s�!�4)�V0�=!���?ym:� ��R����~������m���Ӗ�>��/� 8b��� S������^�E� �������<&�<)a��j�I8A���y�� )#=F1HA)�-�\ ����y��xi���U&#�����IG<��m��)��LVn�ӧE� 8d����
���d������'��E:\y��0_�\ZB��-�*�7�VL�lu(<�Ղܬi�P��R�D�MY��b��$�Ob#=�{��ӢJ��y؄�"f������y��,J4]b�S�X��dH����yrY��4[��"OJ�<��S��yr���9�\䨑�xxx�bU'�yr재Z�8�;���vCjn�>!�!��#���B`*Q8����JKN*!��ޝ!$���2���H�ޔ)�!��͐a���S!"n�J��J΃I�!��۵0�ZH�G`�Ra���A	#`!�P�x���t�[/ �@�Hz*!�$�%��� ������'3!��2X�j�����0�j��p��<e*!���lXd��e�$,rW��*ݠ$�ȓx��
��=t�͠C��z<`q�ȓm����e%��<)��@��P��2h���,�Y��Y/#��%��G�rPq���*$�4E�Z�4py7�� w��ȓeS��r�Q"�V�S��ߔ6�U�ȓR��h��	�a憼��I�r|���ȓ^�4�[�	)J�b���Ê{��Ɇȓk���+b(\�}���[�G�<�*܅� p�}x&��9�H�#���E����ȓS�l!�/_�:y��D��f��Ņ�t|�0mV��8Ӥ!Ѡ03 ]��C n��'o�D�m
�/Ě]�Xم�1u|a���,�F�� _yБ�ȓuX����ζjm��)fk��xɇȓpzՁGi��
���=3�j$�ȓJ�9"����d��$0��OL̕��3�J�8���=@୻wI���ŅȓYId�ه��J.�Hc��<,恅�{PD[-�	~$m�G
@�1
p̈́ȓ4��4�;BM8T��'[q��|��N�Q���\�{>�"�����X�ȓ��ŋ1G�(5���	X0q����fn"�����.<�j`���p�͆�r�ԥ�B �1Zȍba��6M�����?�����X>��4�U*~ �ȓ@� �!@�uZ�����b���Av`qaQ��%t_��S��Z���ȓi����!�S++�������FEx�ȓ:]�g�f^)���ƀ
9�)��P� q D/9���;#�:e� ��H�x�&"F8%m���C�6O,I��SS��I6xu#�ŇSư��ȓ�`����O&dҜ����V�̆ȓ}�2��&���6j�P�W��0r���*9���VBѷ|#����l�!�$�>�u��eP�B�žij!�d�(��i�g�@$C:�zJ��Z!��	 ��6 AҤ��&<�|p��"Oؑ�͚6G�x�E�ۅA��k�"O��� Y2=�J�����\u�d�W"O�*ǯ_V�&����+Vۦ���"O�P�@��=��P0�%��$�a�"O� ���w뎌}m(�����?��t(�"O���$J*��jad�$H��у�"O��-8�وQ�19� ;6"O�骦�6m���-V�@ ąp�"O&l��=.��3NN�!Z��Z3"O����OtSG�>0��3a"O��P�3��u�%�aX�"Ol�f��)wV=J�/�D��u"O �an�����"��i8��y&"O"`�w�W�G!�&������z�"O�\�«��O̐���U��D�"O6uH�ʂ�dj̘C�2��͉&"O�X�����V��x��ȹB"O8{�lQ�6g�=�C� �x�bEX�"O���Be_�#^Ъs(�mu�Q�"O �҈> ��j���:
b8�s"O������lz|Yq�S�~����"O|lhTMW2��ي�@�6;+za�"O� �$k��p�*�����&c�"Oܝ�.<Drp�ٙ&��\Z%�TS�<yЯ��<m��0S�P�k,

�Ek�<����2�������H�i`�c�<�d�	A����dD�eE�6nF]�<����r:Zu�TFݠj��A�b��X�<a5���h�\���G!z乘�g�U�<�T�
�Iv�p�5�&>a��,P_�<iF��L�A��ڃ(��!�b��]�<! 	��^�JA��a0 �S���b�<����*~>�Eŀ8o�R�ÓcTZ�<ɤ�\�8c&��=�~M�(l�<dV)<vnͻ`d8�z L�R�<��噁|j�0���C+�Pf�<��	�rW����
��@�$��n�<Ѥ'^�~0*�i�)\ h�n��Ŏa�<	���
j�h�V�� �)�{�<���kW�#���jR-��
�t�<��TTZ�f,�^1�l��1�HB�ɖ	jiP�I�i�p,2�$�0$. B�&{����+^&�BXA�%d�B�(}��K�ǝ�+�DXłЪ[��B䉦	�α�nx�B�čWIvB�I7�2�ڑN!In ����x	�'��!�k�$Aθ��H.
�:,��'^���P#'���i��xRDD��'{z��Q��'S8�AE�����'j��y���)���+_<	���'Y�3��ϷDy��	�T��'Txd@��|k�,���ÉԠT �'^P�*'@ڽ	�DZ���?t;v���'#�����N1P��53�.��'�j�p�(��) �ϣFd<D��'x"�#�-�oȽ���4�n��
�'%�uq��R��0`���5�X��'6 �ᘏ]�2];�E�,�>��'��$���(�>ٙ -
Lo�t�'���+�� t-eKA��+��-
�'��xJE����a��#&6�t2�'�D܂E��Q�N�*�9a�����'���"�ON\�ͨg&�	d&
%R�'����C�C���(�g"@���=��'���W�2���7	�p�<�x	�'�,0��X�$����G?Y�v�'��r#�.�tó�	5M�4���'���3P;�VVK�GT��!	��� �A��c�+.jz�C#��L�@�1���R��/��zr&�H<�����AO*�'�[9��>	h�+b����,K �n��sh�=$�,�F��y��)[�2��L� ӲŻb��;����C�m�W�L�w�t$��C���'����+�k�7z}��0�O�>S>��I�?W4E@J+W��p�	[2�$�@�Z&dSX�Z�JK�-��� J#��$��(�rF�X�L�/`�6�ⷠ���HOÁʅ/s(��/����@��˱�
=V�:���Jܻ4žd�ɤ�[�*�
n�ʩ[ϓ,z��&�8�ȓG��y�8mڏ���q��|��X��O�O��X��o�� ?L�Pa��y"�%��h�/}�^������D� l"�q�����0��m@#̖�H����H ��.g��E�g�5��p�T��"gI~���.�3xHhd������0�=�O.l���y��y!c%��آ��хt��{��[j�$�.Eh�Z����`{��<�S�9i\ȕ��&�1� ����f�':��4N�7+�RY:cf��u�'l��h�7�0jB�d�2wf���F�)S`���9G< {ϓ(�t�b@�
z������C�4^��l��R���\�P�i��FK9��O�i�5�J�W ���kN�1JP�FK�]_����/�y�D��t�6��S.����:�Fp(�
l�$�����?�T�cK���t�O���17�M���C�L'�&Jܢw��E�'����(|���D�.~�hҁ��#@|�lB�L�HO���ߴ��:�����o�\��X���:�ε��S/~Z�a�C$�+Q��Jg��8U��D�e��<���OBPS�CT�,��Q�nL~+�Ɋ�Vl� �'�:����_g ����ʡu	L�+K<��a��E�
���6��Q̦ �bK"�����T7p]�Ȇ���N�LjtԛFg��M�������I�[��S��L<�#�H��!]_��З&�jH<!��-c�.0��ߙA�Iw`�3���b��jM����ÅP�Be(P�֋#<��@u/.>�OR՛�ˏ��~B�ެ@vAѪ|��
?�"q��̣���1��M��y�n�c\1���p�"�ȀC�,�*Ơ�\�w$�CF�t$��<y�KD��-1�Y^���9�%SF�<�E��7@� fʁ (�Y�oY\�Ià�%b���"~�6���N�jAщZ8{R����%$}6��d�<*�!R��~��֧~&Ţ�G�d f�A���y�`''���R�E�o���j���Ș'���:+�ML(E��:v�0�+�m a�T�bK���y"'�	��2P'B�V�VY� �]~,��`A^o}��B�I�D�$I��y���-O~-�4Wr<���6=�>C�I�W&IeɃO����@��$Z
��0e�6\� Ф;O�eP���)
P2yc���
;F�s�e܋ff�]�׍�\fazn�27�:ի�E�����㘊s��q��1k���!E	5"��W!�U�,�v�'�
�UcT�B�	#`ӳ6b�H�y2 ��5e�x�逎Y7B�21��2<)Cc&��%��d#�u��p��oHD�X�hé��y���8O@�pg��(�t-(R��=�@L��$�u�,�W!⶙��/��9N1����w>���Q�9J��Qr�,e�Mp�'[-;�@�D^���#ĔS��ȉ2�0q�C�EI�;EB� ek���u��8�}Y�}�ę�JJ!2N��6����T�B;�0?9a �(tb�eU���X�Ϋf4����uSD�x��@
v��A�'��җ*��e`(���Ʀ:+�L�D��Z�J��M|s����gğJ�&���oߺB�f%��*�+�j0�FV0RK!�dN6L��UhDdտ
|������\1�dENN��`ϝlTt!��CO4O��Y`��Ɇ�g���jr�P=�:��k�=\!���	5�:#S�z�!�j��e<�����X"0g<���!h�R%9�?i"$��ɁZ��(oʠ�bu�N�;!a~b'A�D�zdjZ�5��2Əybn�h��Y����+��Fk씸g��H����Ԃ�h�xdC�K߇w\xk�*��PH�s��i�f݋ .@	j%�T9��9~�!�HÂMd��ҩ\t�u��ɲy�B��~����ةr%����2\��k��Y��V�K1G�`߶T9��S�;.��/7ll��IvL.xB�	�D2���`+rm��kvA҄7�X��C�����1׆Y8d*m0�$�-�Qg\�;��۞\}V-�š�$��BSbP�F��#P� !�u5�%a�d��a�
2�	�+f�99�Ε�Z������obj�G�;Uf(��Ja�����ٺ;�D�]p^�م�¼3��0q�e�R�<� lqR0ڜsVR��CM�������`B�xKc��,L�DG��I�7�2�9TEYI�=�'��*�y�+�$({jP�@�J�b�YG�R;�Y��ǆ @�nFt0$ᙋ��yb% w�@x�LБ9�����<�Px�# ;
)�\�b�>l����.S2~����bʄ.�x���
[�: N�������y�d-��i;<O���5��x�`%��O���ƪ9n�y;Uɀ.L�nlR�"O4�K�&ϙhU�� pF	���$D�8�}sço{\�q	�|]6x��E7l\�܄�p�*�e
 ;?8 ��
�{=ؤ�ȓgc̱�M�@jidG�k���ȓD��0[��� �&��0� �-d����{��\����:�*����PrLf�ȓ[�VI��ǔh�W��1e�͆�S��4BdN�$A�X�l��d�<��J�b���"���@�i�[r
��ȓ$C*i���Y� =BH�%�%E�0�ȓ6A�U+ġ
����`��az0��%�=@v�\�6>�@�4�^�?�L��ȓRC��R�*=�Y�G�N��!�ȓ��h*�An贮�7�v"OzD�`MP# �a�@C�)b��	r"OS��۰@�����B�>x$<��'H��)�9�"��P  2�<��'`�+�	K��)!+�/,X�'��u-.>�1ar��A��'e�	�$�1h��� E�^����'l��JVm� \&T�̒;�9��'�J4I�j�4L�di�m�9�NEH�'�lZ�9cњ�" �:9 ,3�'<�ae.�{ь�����>q�T��'`���VHպq��򋃙D�hl��'ҥs�g� ;�����E�pȃ�'}^u
u4a,+�V	�0��'�4z���.�������&UۆY�'Y~��e���&��y�Ń�B�X�	�'E&,�v'��:d4(�AN�����'���[d������I�%��EA�'���C�#ƅSq~����^�|��Ey�'F��c�l���P�� ��-�ZH�
�'QH�;Ƭ��|Bm�!$��'��z�'r<��a��"N�b�b�.��x��'���a�/ck���ѣӪ��H�
�'�Xc��EB�V����
�
I�
�'A��ӡ��l����AĘ����X
�'g�Xp���.ԥ٠���z�RU�'�J���*x���s#��r	l\H	�'��M��j�dq�Ga� �PM�'��L3rI^�Z0��@߯,���	�'�x-�2O�r����v��8,����'���*s�� �D{�C�Ai�$��'g��s6��	\mae�L,��H�'�I[wgZ�|��%iE��HD`�J�']����\ع�T�
�3j���'�z�:�	�T8E�#�!����'n����	�,8̰Yn�)�ܠq�'�"�U+wS0b�\���E��'>�x�5��=��r,�{����'pN(���ig�|���.���'�`xR���Y��Q'��	���'���i�W�k ��3�IН~M���'��=S2��BY�$2����{c̜��'�^a�&�ː~ dk��T�h�<h��'�MX�K���Zݒ$�ك��Ġ��� N�Y��W�H���)0�ǒnQ��"O�U��G]���"EFɲ7	��y`"OlLsD "F�÷֍QH�0�C"O� ��@�c��K3n�?#*!�"O¥y��N�.����m�0\y�"O8H8p�^�f]r���H&���w"O,X�5i��lL�W�ޏq�E�"O�A�p��K;�u�g�$l25p�"O����� *@�l�!M�v�� �A"OYND$2��B�G�b�Ua�"O
�e�9g�\er#L]�]��\jc"O.�Juh����+�0�2���"O~��u���f����/�<�U��"O1;� ��3�`���HI"Ox��dO�:�8�@M�!S�u�U"O�P��׹
+�	�G�ֺS��#�"O� J��R!��C2��^�(-��'$j���b�	aԴ�'N K9��"�'��=�n�N�BE�l��E[�0��'��|�&[�u�F[Pŵ8;�t3�'�F��#�W���cAG��2Y^��'��ܒ��&S���B�;�*���'�$�'*��	���k��9/F���'p�Q@pO\�h��(.M3!ڪ)��'�N�9���(�����NAI��
�'T���AD�m�X��NI&[�����'rz<bE&���(�b�ϰ_zz���'vZ� ���<H���̃M�u��'�bar���?�~��pC���B1��'���-�4TAzm���/b )��'�xHDoG�0_�ɺ`~����'Ԫ�ÄE�G�J((%�A.&� ��'v�e¦[<$θ!ڄ2}ȡ�	�'f�]S����<5e�v��n�	B	�'��|K��*v�Aڳ%H;m����'��xD ������+�a�@q��'�"5ɅǛ�x�5I%ZFP�
�'���f�R=V|$�"PK�#
��
�'���
׼b5�=�MϷ群�
�'B0ˇ������B�����
�'�$�8EcH�ː��gE�}���1�'=.z�j	�-�!b�`T%m$d
�'����ʁ8V٨1���X����
�'SH8a���C0�r��E� ��	�'t��1E.U^�� $��B<��';���&|�x8jū�@()i�'R��B3늾&��d�� �43�����'�V���e�R\�������'&��0���[\�t��j�6�&��
�'پeyuC*e��)EE���'x�����g��P@*��~*�b�'���$@F:B&)Je��
=�ث�'�.��D�!%t�P�K5!�R��'L�I\����I��bKP���HW�<6k�����y����Di��JS�<Ʌ��B88t�5�_5�����%L�<�@���{m@d�V�m5V]zQ��I�<qQ�VFQV�­�9N��y`A�<�/�$]0�f�&��i�ǖB�<����\��� ���`!5NV�<�'d�@�\:���Tf���Y�<1!�1C�"��1��Z�x\,4.��0)���,ȩp8�VF�<` x�ȓ":�MG`պ @�u�>L����S�? �x���s��j�)�+�0��q"OB|3�ǀ�&ʡ0䯐�D�V�S#"O�$����M�Xq�v��";��I"O���A���d��g���)���9&"O88a��6X��t��2��������a���d7�z�M��BX Y�@�.$*���R��>�7%�j��� d�+(7t�	`����ɠ�%�?�y2$E'H	8�Gof�IJ�������^.!�1���+����tɁ�%���'?��M%)"E[��Tp���Ҕ�N�L��}��NN��D��B�)e/&@1��G���0��̳-��R��f�hD��`,?��%�矜�Q�T�e�b�Y�cЊ1>�)�+"�\DŐ3�X�j6�4�H%��ˀ�l��/D�l��p�E�!B�DK�Y�L,�V��Xq����CV\!'Y�0��9"F�=�VH
* I�����?5A���S�=3A��1q��� ���@Eʄ�iPqID��b���!P�Hh<Y�*�̸$+����Z7BJ��~��$\}��@�hV9RD0UR fH�'�RTA�w]��g�/c۾ZR�Q�`؈���yľ9�!� R�U�A �H��.�QĲ|����>m�`�"���B_j����'� ��q�ՠfb�`{� �X�����X�L
v��B�Q07e�)P �;�$�dT�� � G}8���`�͡�yb��Gjt��c�*W�y�HߕG�JU�%\6kZx�q�,�.�M��HW�O�p���
8�ȕ�	8�-����*����ɢ���c''F�Z�T"O�m�rC�5|l���Ò ��@
�o]+5VY��f�>412�q��q��5��IK����
#��@�e�U�D���`��:|����:~����<g�(q�dIJ:u�A�CAn��;�K�4H��V�|b,�'k� Yى���<��U	�$(�P���I 3G�0�E|���+C���re�v�"H�X>��eN20�V�QIׇm�bT��>a�"��K�<���W�Bʘ2�q	@/�����jR�x2 �5B7�=��o�OxR����z=,�� Oҟ~uJ��	�'L��߰d��1C �E�G9�]�b� J��	�|`����x���	��T!`��ki�a .�(��x��B���*6E��0���S}�l��NH�fU���ɥo��ݙ����D� ����<{�b��P�nO#��ɇQ��]ڧ�������R0�Ƭ'/�x��d�<$��%@�'",�Ia��C� �
�g�� 3Z��sbN�	�=���bV_�O,b�͓ N:�	D�_�+W�����|�rȅ�;��x�K;WT�P��-�;Ivx�c��T�J�[e%���Y���
|Q�����?M��3w	�("	����%LOԉ��.��O�}��'v�YXeժz@�	����3��'��P��eĊ�!VE�7O�Thj�yr�D6J�LX:�/�U�υ�K�����)>F�*�yr�V�^Yp<�Dd�n$�R�"#�v���GC��P�FL>�tzL�4�N�v �iǋ�f{�L��T}�`�ğ�dc��AU�Q����E�qf� �O��V�OIT
��2Ϛ?c64��G�'�T�Ǎ3r���Ql�`��ד
jD�� �|�
�ȓ,<@G�:U�t�&M+����<领ͪ���!a�B� v0����T'��=1�)]��\Pw�ˀ�y�$ĩ,J=J��ȴZ�$�"�k@�$NH���Q�V��X��i�O,j��Y���PK��S:8+�EP�$R��E/*D�耱�G"d|ذ�C %np�`kk���X����h�r@D�ln���l�=ڐ���N��C�S�:a~�)Lg4�#3Ŧw�%�� �\U�T8�ةF�Xd�Z�\�j�N��o�`9���+�`�G|r+X�Ya�9!�m�lܧZj�P��.cU�����,v��ȓsʘ�s$&R� ��9b�C�]6�i�Fg,h��]4ҧ���y���2Q�4�����#�Ѥ"O ��b'�D��ԡS�Y&k�X����L�3�U�J�>ؙ�'z�0�OR�v��D��OO: 1�j��^��3��3+��1p4�F:Y�*E�¦Åy=�h��=�(��O�ɾ�6�8D#*�|9���d��|l@\���_��O�Lpaթ��Og�|�� FH�%��'��kq�2/�
)y�-T�2m���'��i9��l�ɧh��I��h��[�P���bY")��"O���b%�;Be�Q�sB�8v�g�xҧ9t��)� BQ��]^��у�"(.l�u"O���V�	�%_�pJ�j^��6���"O���ɏH�|(	B�V;.�\��"O"�{3�
@!4#e�H�ưzW"Or�ʇ�G�q���A-��iqT"O�I#���!>�@ G��U���s�"O`D��JV�!a@��+C��t`�"O ��5�0��CG�G*��9�"Ov�#PJ�	2l��)��b�̨ �"Oh�F��<Gdh6dԞGh
�R"Op��f�)!-�e(��֜@{���"OȌ����׃׽8m��ӕ"O�:�o��0HF`�w��5L\8��!"O&�p+ؓ-������؜!,�m"�"O��A��@:L�J�xcI��v X��G"O�<1a�4KL>}�7*Ļ�� d"OD��K�P�x�ؔ�O�h�&ق�"O-���0//<A��Ѓ<��0��"O0���l�YD�D;
��5�д��"O~	�KE
z0N�Ä�!<f��P"Oh���ڋ&���!R"C5�̳�"O�l����rSr��k�0 QJ 8�"O"@��C7-�$�еo[ BBP��"OI���wx����L.9��+�"O�L:dIU�t	R�S&��zT"Oԭ�χ�	u,��~�v�"O��E�	8�i%"��w��� �"O��%��˼������t�����"O�Y2 �7��[�+VJ���8"Of9���m�T�����S�`H �"O�d���D�a��ɓ�+�ƕ�"Otl�ܗtY�!Aiܖg_�( �"OdU �
	_��Ђ!(=3$"���"OĄs��	7~�@�Ԛv� Y(a"O�|j�N�
^93&޵f�j<�T"O�THf-�-*�XH��8��l�"OΉ��g[	1`dh1�E�t|�0QW"O};�F��q��$A5dWz���"O<p�������5Q�	>!_����"OΝ)�`�;;��ѻ��*C>��"O�a�i f�y�a	�W�+%"Oެذ�!��(ʰir!��"O�9�&%"����!�>l*0"O<)3�^���QDO�J
l�g"O��9�LG�Wh`x'�A�:S"�"t"O��w"/����/˳nF�p�"Onx�c�U�*.�����dsH���"O*���ț�"�f{FH��$g*�He"O4�#BG�N�0��G�,Sn�#�"Oh�qG&�of�Ud ��>�`I�P"O�u�toهެ�d�� _מq�w"O�� Qi��cت-�q�ӯq�Bd�A"OX=jń
f���3�����( ��"O��JS�$J'�����;"�5P�"O��!v��x�`)�U��o��("O��Z��
�US��ۣ�P�$����"O@���ȫ$����K�޴�7"O�(������
Nh���"O�r��`�T�E���k�]��"O��d�ىx��L:���$��4�r"O �͖1��$���1܈4y�"O�b�V�@EZ $+H		 9�"O�� !��5�vxY��+��JE"OV��Q��=V"x	���D�Vi���*����� ���5�W��u蒄(K�A "O��X�%��q	��{6�pU"O2�0��S�r��`Z%b��&Q,��"O���$/@�^܁��+�5T(f)ۂ"O��x� ȺWp��E��C"2<�"O�-��M��f��h�ao�/4��c"O"E����>O�1 �ͅ3K��I%"O�iT�S5QH�5�͟HR̼q2"O:��IC�=��S7d�3M4����"O��5K� g���Mڕ,� �$"OPq��	;��k��(b�=	2"OvHi��s��8��`ldD�3"O��شB׾L ؉U	�k����"O|)iO�&�.�5��"�0��"O�\c���?�ICK���L@�U"O ��� Nj���$�8���'
ʢ<�[wH0-D����h4�����%��́c#�P/�M��=���0|b�*��u�%r®_�B5�\.d�1Obug\o>��%͈6g�܂�Ȥx��	�3�D�K�&L��{���	�&��`�� �44�4/� ˓�Gx��i��+�dI�m @��`���\�5��Ėu؟l���@
�
��$���M�:D����.+��-q�������V$5D�4M�.�ӯތD���jf�1D�$��$R:�H���c�/]�>�;-D���
0�m���=+�a1m+D�DR2�Z4�6��UE֡	����*D� x��?l?�HK�bP2A��Ż�k(D�{Bт+�QH��M����4�(D��@Wi��$�˃�M�t���,D��"V���M���;׈̠$>��+4D����*/�V��Ŕ&< H;�o%D���&D��r-���"V&�H��7D�T�tC��Lb�H�PjL?���1`�(D�܋��P0Ukv��f�IQ��8���%D�\�b�s�T��	۹x
�LSv�$D�t2���$>Mzѩ���!}"T@�w6D�H0�N�<���	t2+}����3D���`��7��ݳ�(�w,B��WO3D�(����m(a��T�!1�i	�K3D�@ �^�P�R��o~�R�!'D���%�7#�ب�6(Ŀh�,���n*D���V���,�:y#���5*��D��c5D��ʷ���(����� QĦ�$7D��@��o�r����+h� 1�3D��i�g"@xxf�[�F5L��3D�@��b�f����WJߺ�>| ��/D��QE)�^M��26��`� h;�/D�t1�@fD�s��W�H�$� �#D���B�H<�^B�ĕy��i��!D��s��.\A���4n�CM����	%D�$ �h֟O����)I-��C�8D�����R
N���GmNeF�Չ��6D�8 ��\$��࣐�
I���c�(6D���f�
n�(Ӆ�;�P�Ȱ3D�Ppi���U����ZK�� /D�T��5_2<� ��*E
ܜ�W�+D�H�c��>�1q���~v��V+D�9fہa=h�sa��j�+ԔaO!�#�����C����l��<�!��^?�t�mֹ��L
�J�%!�!�$߭u�P�	�^�f��@qS�� J�!�d��G�A�Ql(ra����*�!�D��	������%gc���C�`!�� <`���,?h��f~tDxA"O*tS����8�k�C�cx��%"OR	��K��
P(�!�#�8/�� �"O.upħY��EG$�.%�n)s@"O0�+�ć�oU�=��#�51��e�%"OKM �ȝ��c����Xk�'��y��'b�ظ
�X6}� ���F�y��&=t9�`�݈pV�2����y���Q4���
3�(`�hK��y��D:d0a�� �ʌ0q�
��yRHO��"�n�|��(�̘�y�Xu��ci[v��+�璷�yRd��M�.�V��b�j�#-M�y2��9�|�&i�.e�xZ�����yB�S���HV�=�:I�c�Y��yb�Y;l�DAb�ʕB�hS LS,�y�k�"=�<�#��B�=��'���yrN;�Z�k�/��I���!�yb�ˣ	�<Mb0J��{�0����C��y��	�� �+��{:�Qr7b�y��g�C�#G�g�p܁ �yR�<�:Q8���`�f��,�yRL�'mH퉱?cc�d�U�_�yb�HI�ڇ�٥)�~m�e]��y-�b��ٰ�ኌ��+O�y"(�E�.��o��!�Z��cŉ�y�τ�
�D�[rj=f~r J��yFK��8�֮�6
����ܶ�y-ȤL��h�B@'�"h9gL���y��A�[�*�pBhG�(���X7�y"�O�9�.�I�A������y"bJ$zvI
�LB$b�;d��&�yB��)b�  �~�zy�C���y��E�m�t�
�B�cBN���y�!L��\0A��l�ң�.�y�'�'a� ��&&&y7�,�QΘ��y�IR�W���!��	?}�]k��&�yR�[ݔ� 1 ޴1���{`��%�y���G�$�8S�X�(�,���&��y��W[�j� �
��us�I��y�F���-k�䅘
����#C*�y��_n*ػt��E�ak�E��y+C�.j�C0%�?FؤH�# ��y�D��(�R�-2J&L��aH0�yǕ�L�$EXF��>E�d8�A��yb��c�lH�"L���h�*�+�yr��O���р�X4|6��to��y�Yvj��3Op��IKԊ��y2^e.�\��d��g����B	ɪ�y�§P��]�whĈt@}��b���y�%M4@�T\z�fK�~88�ו�yR��X�Ѐ�W�	L���ŭ�y�OL�7�D�6��{6��KƂ��yp�>��\�}X�L�C�y�F�7z��p ��E�`EǠ��y���]J��5�P��Jܐ���y2hS&0�8�1F(͵���b��y�)�)\8��Cp@�)7�v��aaU��y��K�̹""*	Z)x�*ц\��yb�ϟPP���W4d�~@��J��y��l�I6e�*`���v��(�y2��S��p�(�kK13��y��W��Z��A��i�DՉ��^>�y��+=^�a���VƵ�h���y
� ���f�B�v�k�
���,(
@"O�i��ס=-�Y!�D�@�����"O�uctl	�I��YP�(ح_X1�4"O��3U`İ�
tɣt�^�h�"OXq9�CO�}�lP �y-����"O~�[v�Q�,%���1���8)��"O,�0�k�t�IAv�S�`}:]��"O8`��Ύ_:�!���?Z����W"O�D�dOO�8?z�֩�-�ܽ t"O>�BO�]Hk׮S��A�"O�$�l�y��m�5���@�S"Ox�!!���4~xh��@�8�v�K�"Ox=�BI��dT0��P�K{�����"O&� V�ަlmB)1�HbiL�(�"OT��Q�`�>�s@�ɴtUR4��"O�y��2M�����FO�oG�t��"O����|�"��$J?b �k�"OИғʃ&X\@�N�C����"O@�2D"����Y�J	Cd"O���T���1�M�����BV"O���Cʥq>Je�P�A��x(`"O��R DO�@~��9k��S\�,!�"O�]���M�C�^���I�E�i4"ON}c���x6��ҷ�_��U��"O��P��)�fl����W��` "O���O��zs�!���!u��"O
�H�
�4�Q	Lx�܂"O��"fK3f+dI��D��:o��S"O����� OIX��'E�~	�'�H`��^�\?:��1��Wv}i�'Լ�q�
	jRȬ�Vș�"&&Pi�'V����֕iD��6 �l.�9c�'� )����K�1�VBY$jL41��'$ clwaD��4W2X��E�<�yBf�z���9A�U/g��0𔠀�y�	ӹ[�t�(�Ĵhp��X�!�yR��;-j"�wCV\X��Se���y2@�2ː�0#�X"!�H�Ys��*�y��J0&`��Yz�Z���y� ��RH ��g�? �4"0�ʶ�y,��|8��ʀ	j�,qk�yr�N�$Mh�&߶eM�rc���y�Dh���"�4aͼ$�R�R�yB �2_Mj��f#�]G�=�"�M��y�c�Pl9I������@�ř�yb� �yI�С�`��zp&�"��N��y��9w����ՠ)aL����O��yB�B^��i�m]%�d�rc�L�y2H��H�Js���'!iv�	��P6�y%N�2�4x���6�V�W��y�����$�ЩJ1CO>���g��y�MD�!q&,����4�d��Unܬ�y�*ŕ=R�1�cA�&\�b݁���y��P�m�3I��|k.|��hް�y�è����S�t��)P�ȕ�y򫟷f���'g!�趠١�y�_�t�
�!�	K�<��Z��yR��<h��8e�Φc�m2�ɏ��y��;o⅋p�Q���L`dP+�y���?�1Ąz�@5ɤE��y�3_:L<��	�
oh�Yt���y��� Z�.q� dq���0�F��y�MԤZp�d�r
ʼ(����'���yr�\-<��<�u�[��6�Ӏ�y
� � ba����xK�G��'4����"O�h��F�&�����7R�N4q'"O6h�� \0�&큒F 2�tA�"O�щ���-W�I4١\��-��"OƐ��+Ў�Q��;.�`Y"O�\Iddk�.,zui�9#=�-�5"O=�ς"q(�Q�,W-��K�"OT�Y�,֦o��l�ł�X��q�"O.Db��3f��X�4f�-B��"ORH��
G���$ ƒ.Y@92R"Ozq҃���REУ���r�h��"O���������0q�j�\�'"O�3����4��*	�FT��"O��Mq��hS�
�9iTtYb"O~�y%b�,'W:]���~`H�IP"OVx�Ad�"%5P�{��i�"O�9pA�Y�ibry�t�ӹ����"O��a �D�A�
!h�b�,K,=�"O�$�"����0�E��%�0�yro�l4�"��V::���a��$�y�"�j$pCT�V;�B x�'��y�HL	f� �$r`�Q�X��y�/���b�S��%��}�!B�'�y�L,>���M������bW��y"��2),��Aqf�6A��e���y� S�\
����5����!���y"��+I�P2�Jܞ/��	����"�y�yh��
WJ�T��1B$�Z��yb�ě�T=� M�Q���-mN꓅?y��W�xi���?I���Pl�����rj�c��ЀzW�L��?YC��:_�����:{B�E�Rt8s� �{U.9³�84*��d���ij2��$��d�NP��F���a��5R�	C�P�nԐ�/a���'V�C5�'�J?��?�ߴP��1{D"��z>�Ԫ�ɋM�U����?iBK�I� ٻЌ��� ���}�L�I��h޴�?���i#��?��O�ޝ�w��xTn�A8�����]_tP���i�"�'��|�O���F�g�����*DfVek�`K.,\1k�`�ڰ?��͌4E�l��c���#� LE� 5���>9���ͰAήF/h��P���'ސ,�2���?)O>���?IO>	�����s�Z�
�����(UO� AT"Oh]�P�*;�U�k-Hn�ĳ@�>��i�R\���Δ���d�>� aڼC��D	d�ڲ���j� �'���'.I�n�H���O�l��t��ڇǰ-:`�5��,��Ojmb��'l|D�ЃGU$~"&Ye���F*��4�Q�JƢ��TP�$,"G�<�r�4A�����ݴ�?Zw#�%�jJ��ebqfR�ߚ ��'��_�<��h��p�f�9S�`����Y�������'P�Dd�(6�'9��8i`�N
6
^��To������)�M�d�Y0R���'��J�t�'��&N�P%ܬ�ug�!{� �b'lA�:����*kܓO���/��ON�y�J� ���c��u�2W����X�L��$����0|rcgPx���ǀ6NlT�C�c}��կ�?1����O|��v���_f���{2
UǺ�c�>����hOHO8� �O�$;d�$�4o��/O*�1��ɶ�M�����OPy��*��v�I��<d������Onʓ�i�ǿi�b�'�r�x��ǫGA��׍�*<B�p#�(�~"�'=�e�!�'�F���	B�He��*�0.���IX� ��Dm�P�rKf�3�I52��Z�E��<F�y��b��Tt[���G�O�a�J|�IΟ�ڦ�S0E�d�c(�:n�Fa� �,D�h��!��(UV�0V�=��x�N���r�4���|�O���T�X[�ǃ�U�l��'wvL�E��HF<d�ٴ�?	���?AJ>�'�?�"��M�b��!h�\�:��T!gp���TJ؟�C�b�t��j���uF���,Z�dՋ�,�7\�Y�n6��?X��eυ/	0QCޝ*y�9��6���?������MIw��p�úd��0�k.�!�dچU��r3��6�YZ�.�?]W�!*�vqӔ�O����O��(���  @�?   �  �  �    @$   ލp�F˸���b��P5f��p�>I2�P�?)����S�$�F�8u"�7��+�6-!lB�ɖ6:|�(DE����t��C�	"&�2́a��z~h�eϧ@ӌC�A+,ɘ�I'\	~�`%Ϲ>tC�;zh�x@���4e
����gˎs���,"���^2.�9 ��}9����ƪt�2��b���9���O>˓Ol�Z�Cړ6�4�7�_�j(��ȓc�x"��
�ZH*�LT=ovV��ȓDٙC�Q��~��gR�>��ȓ�~%� �%�E� �B��=�@�7b[C�H�qnBn�~H��G;��HHG�i�㨑�6i��}�L`M�e�����O����/�L��@)�v����"�!�$�z�0`�j��`璺r�!�D$r��(����ʄRu�9|!�DN=w���#�6��E��&*��x��'�w��Z��ު[vĭ�
�,��z
� Ex�Ow�'�ɔ\:�����-��)�	�?
8C䉩r���ч���A�����?@JC�ɷ?n�yB�R�ѡC�&�հ�)Tt�E��E�R��B�C���r���Tu����F��M���'V#=�5hA�n�VM�P������@��P_`���'4r�'d�|J?�fJ��	� ��fgU� ����^��s4#�9&�$����~8�(YE.��C��K&)���$I���|��`�kT��CG�k�(rUn׮�y��DEϟ8�	���	Fy��'��O�mZ%.��
�ʙ"��1�"O��Qt-�Nyt�ЇD ����������I\y�%�&�RZ?���J��,�20��0���hP	P��?qH>a�S7�X�gI`�ObԠ��/=<����1�򌒗�'8��4��o���ލ�p,�;l�H@�D�!7'����؊%��'\�I�v�J|�2hٙ	�ܠ34$Ӏg��I֟d�	c�S���1�����4�#�;a���?��ہ�7K��������9�?��B삸���ӝ4��`ug��`���G�n�8�$�O�����-v<������J�*��σ#!���:��)(R)�c�B%(�,B�!�D�1� X�s-T+�&��ː�2�!򤖙�\�dDɥ&kvHද˛`��x�C,ʓ4��ɨ�k��P�d�)��K�^b\���'��'P�5��
�D�O��0�d�2�L-S�6�	���/i���>�0��XX�p1��ة+�a�ֆJ�t��.��+v4���D��0h�}8�$�䦂Wr�a����ɳMo*P�)�<�S8�0��v+O�g�V�b�3Q��$!�'b�d@Aʃ���`��cM��Њ�4���D�>aE���^�L�$F.A�W��(V]��0�'E��'�Ҕ|J?� ��7U�������@ڶ�;���C�I�b��U�7�A�-8.X:�Ʌ"l� YC m2�H��	�t��P��ŕ0�T�R%K��U�*�������_�*Z�lq���!�DE�l�B�K��I�CN�(�aBqO�inZH�'�����R�Ȥ����"�p�Fh؆ Ӷ#5�'O�'���Y����$׎�Tx���uB T�6d6T�(腣T�+H$L*�T�P0Yc$"Ohu	��,6�풆��nb�7�:D��s�V9g�#D�0ypp2&L7�(BCKI�z��Y��\*0� �Qc��7�Q�HQ��"ڧF�V(��f��(=��	>�Tj�'��'O�K���~]��X���#�'�&�Zu�Mw�v�h&¢}���i�'R9���-2���*
v-�p�'ov����G��ȴ�2k�(�Ǔ8�Q�8#���?����.�5�TH橡� ��)(��|���?ɮO� �Pr�:n�>5�jބK?�]�F"O�B҆�3xh�̡�� ~:ּ �"ORR�g��$�`� X�(jlA�"ORM�Be�G�0� #a�.1n9��"O�P0�aD�\�A���z����>y��)� �t��U�
�CΑ��.�91��'�xa���'��|J~zaŏ�n+�4�תE;����z�<Y%"ѐjl��1���'��-{Ыa�<!�%��	4q�̅NE��J�T�<AFսe4�Ŋ� R)1�h���R�<16̜�����ĊZ9NX�	3(UܓXS���*�OTȲ�M�,����oZ#!���eJ����&���)�gy⢎�M�)`��}� H�$B��yR�ԋ$|
A��L�n=���c��*�y����A���:d�iT��x�)_��yMRH�`4��͖�Q< �BCF6�Px��$[��Bs.G�^��
�ZVd��D}B���h�*���lУe�9Q�H86j(�2p�BΟ���WX���M����Oqc��#�B�I�$�X׊�g�`���5
TB�	����s$75v��j���	�B�	�Z>���'
�~���$�^$i����`�'��Ic�
H���5Ѳ�U�xƌ!;�'���ۈ�4�����O��=xv� kօ6#��0��)�伆�L��j`��Եx�A�`�\i�ȓY$R�k-�M�9�0a�7}|u�ȓ���hю1���#�	�[�jɅȓ-3fq+2LO��.A��GJ��OԠEz�����Gz M���̎ZoxԛB"�>��&bJ ��I�t$�����B��>���b�9+K�k"O�� D�1�t�hu"�$69�u�"O�DK�H8	'�d���U���"O�U(4+�D�Z���\�u��"O-Yr�B�<�r<��A0XVNQ`���S�'�f����9|$���"@*����7r4Ț��'��'s��Y���r����\��Y�!EN�`e4D�z6��E։����5,�z��W!>D�Hx��O;#|x�����Rٔ��;D���
=��5��
�X	�5l%�8q�Lևo�tڐ���w 1"q�ϸ#Q���i0ڧB��\"f��.�6�������l(D�'���'~��ѵ�\�?�8� � e�8��'�Ȁ���)<���R�ǎ0ĂDz�'�v`��X �����*��lI�'U���׫lD����=�RH�Ǔ!PQ����lQ:�:�wG9
<r|c��, .8��|��?��O&�0�A�,Z:p��K�.1RP��"O��y��V�}�Hd��I��h���"O�TO�>Z"@���4P�)�*Ol$xr兡���t�ܺWl�D:
�'Ux��B@U�W$,�y�oX1J���I�����)T�/yFf��s&`��3��t$�Z�=Q��?�L>%?a��ҏ�\ts �Y� ��	��#D�H##S�Z��p�4
�U'z��ed"D���e�>'0��%�#�DL��D>D�S���}8�	B�T�
�#ǎ)D��s�c�9/�ɢ�e]�.< @G(�(��O.l��'���⥣Ւ0W����+`Q��,�Oz�Ob��<�
J��H�L�e������h�<�)ͩz���	���w�xeBn�<��ݙq�h�q���4/v�<1��W?v
�|ʀ�=oЎTz�Pt(<)#�߹|�8�p��g���)���4j�>1 g�p�O0��`I�
�y�%�*;�d���OD��>�O� �l�1,�Z�" ��[�\X�"O8zC(�2	ج�1�ݸ^�@���"O���%��.3If�
V�E���8ڃ"O��"�"	]4Xx���i��%���'ے�<Qr��=:D4���@�y�ƴ��.E?�U�Py�����'��_�`*c�É��!�	J">/�pjr""D��c��1l��`C#lǱlJƈ&D�c瀀�*�ؼR�c��*�R �GK/D��/A�6��AևP�l\�!#:D�2G�LNJ����#q�Vt:��%}rn>�S�'��a�1�&��P���4��O��bV��O��D=����dP#Z5�h) ���GC��J��y��;�(�B�6D$�5Ê$�yBkC*OX`�:��X1���D���yB�Q�?�~��=�����T1�y�N.V�"9SQk� R�!��и',�"?���ğ܈���6N�| E�])Q����hЍ�?�K>��S���d�)QĄ�;�
�.Ls��&�ʄ[H!��M |�c$,���Pt��ˊQ/!���$ &Hl�A^�J\Kٌq�!��ݝF�J(�C		�@��������On���0&P�W�]���Ǳ^:�J��V�p��>E�78	8U�eC�� ��U�0�L��?���а>1Pnߺ}�1h���n���S,�X�<�f�;B-�#��%��+�'�V�<�3�H&W`ģ��׀:L��31�w�<Y�
	�)"v���� 5uT�c�CL8�t#��׈6��azb�׽`�\�q��)G����TC�������m}b�D
G��y�(B71�e� D�yR��pЂ0:7)!��4R���y�C�7k4	�O�zt �e,� �y���;���A�dɖ+��0DZ2�y¤�
]HvH�@�0%���rc� ��	��HO���Kq�Y�}0��7IT��cw�>��J��?!����S�ӷk�>M��o���*�s`�F�X/�C䉦	;ҥp'�����@�V:SP�C�I�J�PŊd��r�t��#0�fC�	8s�t1Rj7u�L��-+dC�$p�B���N(V��"&��!p{�������mB,���l@�J��n%ˆE�i���D(�d�O>˓&f�D[���,X�#�P����ȓx3^p@&͜`9V(��%z<��Hi^����H	F*i�z�N�ȓw�*M!��˿Q����E�#PD�=� j��K��W�f�j$��E̠����&�kLE��k�9c�� Βd�q��O������O���I2m�R6�J� D�"!!��)x��Xp)۝5��x�4Ñ�!�$��z|�\���BP!����2�!��ـl����đX�R�ꖭ$��xҥ)ʓ=C6���5/�}�7o��>�~4��'��QFx�O.2�'����y�y��i�Q��jS��U��B�R��PӇ��!ø�r�fO�R��B�I�[��Pe�L�h��
����B��kG
�� հ@KnH��%�-d'�B�	4z7m�VN��M4F`�R��/d�|�'d�#=���e�M7j�'*
?�4y{�G�d�������$�O��O�O��1zT뚺xf!��gȧh�.@��'�x��A��_MD}�Ǥ�-��0"�'`�3�K�*z�d@��(H6q>���'Є���^��bx�P���_T ��'����vkM#(*=*��E�L�"U�{�;�7*x���4O�Ԓ���+]�p�f���hH3����?E�,OhH�1H�"`�M�c�X�
��5Y�"O� "�S��N�Y�~1�e�T,[�p��b"O�|pԧ�rzt$�*͒r����"O��:�(��[�ܤ��)�8\���3
O�`@$�;(�BL���-]��,Jŉ��O Ex5�Ӷj����T�^�~e���z��l����?��Sle8&�+�������=u�݄ȓ'|���IO�K����Mڴ��ȓ{5J���B�>I�f��tlڹ*$���`��Tہ�MP~\=:׮֝yV����ɭ�(O�Șu)0ˮ�c5G�>%T�c1�O�|���i>������' ��jr�(U�4�x��#RE����'���tFi��t�F
!F�8�3�'����U=�DCVϘ�8�jT��'��ٳꏼ8�J�ضCZ*F�0��'5pt� #ס,P�r̄
DiZ8�I�ԑ���	�#�J�h���-	=�d�c����$�����?1K>%?� %�Z>�����q�10e("D�8ӂɆ@����˓�	E01%G2D��!�H��Z�d`�� ����-D�����_(֨;֍�*x�2e�6L*D���a-? ����%K/l���a)�ɉ��O�%��'�@YC�ʂ]�2�+����D���O�OF��<��O�nA<(s��o�b���"L�<�2	͓-���2�ɀVn��CI�<�S2fv�}��o�"h ����A�<�遁=;�y96�͇[�)���|(<9πH!"��Q�M/cM�%�Ħ[�[��>y��t�O�8;g��2-�J񘱇ћ_��ݰ���O���6�O��aG��R"]-4���kP"O�E��cϮAP����B���SU"O�$��i�|�Z�&
��e�`"O�l��KW�5�F�P�dA2��9�3�'�(�<�BD��Mj�p�"Pdk�M�"�X?��Yl�����'S��ae��b��
Rcǣ����'+D���&OU$6������˦��m)D����-/<Iʱ�q��- �B�J�''D����O��~��KaA�#AHL��#D��e�G�lMdE0W��<~��D!}�A5�S�'N�)9�*Ԫa
�瞤R��OV�8��O��D5������	)®���f�,������(�y�L!pVB(2�	X�F�����3�!�D�1Z![3-�8�� SI!�d��3  }��a�8~�TQB與+�!�D̵m�|��&l��dׂ���I�M�qO��E~���?y��C*T��E�4�5 �č���ɜw�|�����ɩE�Ƚ8t�+/����e׀pc�B�ɀ}*��ӖD�N|eE
'VB�Ig�P�s�,	4�������� D�H�W��2
|ECЄ�n��b�i �4PvOĝ,� D�,�Xe$���{MQ� 25�?�'Z��pj! @Zv����
W�Še�'bb�'�z��+
,�l�b�OYi.p��'�L�{&&L<N������'a�l��'3V���I�O��8�ц Z�NMy
�'�|�#��	lh�많�eZ�`!
��Q�B�I 7	L���P��4UvI
�`�����"9��|���?��O�iR�M���|8bLO6J�*��"O��a�$�
/�e�ā 9�}*�"O1!�OQ"<@M�����}�e"O<�ZqJ*S7z���W;t����f"O�R%ԀI�a��N��T�,� ��>9��)��(w���QB�;�:��G	ЭW�|�'������'��|J~�W��5U�Υ�a���[�By���l�<�)��b��sg 6*Gf1����p�<� �1���!q�h�d�W+QL�5"O\@�-Sa��a��kùc�Hy��"O��(�@ `ܪY3�	��6�x�{����d�'����A�����}U�y���5fR���'�'g��Y�xȔk�Yz�;V[o�4� �1D�財��6]�+\�u��3CL�qg!�$G>�*-p�%��9l�M{ƪ��2]!�d�H3]��#[Z	��_2PY��ӛP�u:r�� m\���.o�����$�\��>���h�Y�\�ar�[&��Q�p��?����>QNB
^T!��L�潠��W�<��b�Lhma��)`ϔ,r��FN�<���߾�����`T�z�:�A�f�^�<ye�4i��kƥfi!�l�p8�,���N�(���pDN183T,"փ�b�x"<٧';�D�'��^�8��W0(a��! -��v�HD�@K��x)0%��C5��kI9;ۨc?O�1ht���..�ip,U�Q���ؘug���!�R
�?A�#W_ѱ��'�z9�V�E�\+��� I�U��0���O>�w(� �i>�DzҨ��~�T�rp��v�2���y2I�O̾�i� ͎5�i`�S���%�HO���O
�m�T���ʀsA���e�r�G�ֶ�*�'��'7ɧ��/}�:Is���4I>(!��g�4KP  85�^/ l�Ւe'^�	zԆ�I�Fٙ�$L�b0����E�At���#C\�>n\[����M��(��?��M�c�U�AYb0�r�'�m��o�O:� ړ��'ފ5)e��N�PX�#؇ ����'����"\>5��)�g'ݳ��i�{bf��D<�ɼJ�^�I��viV�ڵ�J @N�q����L��8��k��˟"|�'Ɖ#���O4��y1�U�O�|�	�'��m���Й j��P6���M6d�2�'�b�H�e��	3 �JGIX�Lm1�'��-q���#x��.Ǧ=
���h(<�@ˍ�	��I�_�X�l�[���Eր�>a��d�O�X�sD�j��FU%6�tAʖ��O��D/�O<]��(P�3�+vjC%�tj5"O�	;D,�6
�H^b\�I'�֎�y"�DOt�����U
&��΂�yH&gfx�2�B�O:Z�����p<�剞fMZ�F�:>��2��F�0�n�	K52#<ͧ�?1����$̉O���͞Y�*L�ȕ5WS!�r�H��&�9� 1�4-ƴ?�!�D[�>^t�$�ىG��`9 �7'�!�D�v��m���ra�쒥	=[�!�$�)�^���*Ɛ2�$�@�I�'�^����?QhV��Xp��7��)����?}B�ٟpR"�'�ɧ�'���oS�T�)��B�<]�ȇ��L���
ҘX���O����܅ȓ%KR@��aO#�V,�� �.\j���H� ��V�rV��V)�	x�����VK�4�K�%Φa �	��R���=9s�ɇ<O��ğ���y4$�p d��Ԍ@-v�@|��\�	�"|�'
|��A��jڜ����-|ȍ:�'�8����j�����<Q�^���'���A�f���|#�� Qt��:�'�f!���ɏH�� ��:>rL���'LnDj�2��ӆ� \�L�9��C�'�����^�m�Ġ� �֋WC�\�������	����ɍ(��@��G�$'���ѿ4�>B�I~	(`�(Z#`�����!+�C�	�FEr ��\�P��J�)��%C�	^3 �С��At@���ɔo"��x�'ϖ�qLZ�`HԈA�n�%$����'��-�  ���   �  ;  �    	)  4  ?  �I  �T  �_  Yk  v  �|  ��  �  Z�  ��  �  0�  t�  �  a�  �  K�  ��  	�  p�  ��  �  X�  ��  ��    x + �  �$ a, �3  ލp�F˸��%�R(O5f��p"O��QD>]*Q�U
*��2�"O	��3!\�88�Gǚ:¼iU"O���@�/0��Y�R�l �\��"OtEC�/�9A���ӷ�ͬ!O����"O�0� AF�=����^4~XA�"O�%���D<��#o��0<d3�"OHR����g�LQKԋQ�0�V,�"O0)�2�)?��#7@�p�'�@9�DO�F�n�9��,~B q
�'�ֵȑN�Nݪ�a��
~9���	�'?��*q��X�`.&q0�(	�'�8��A�X��KQ�Y�a r�y	�'q���`��0�b7GK�/�jL��'��)`2�Z7r�Ұ��$��3�����'�X�8T��x���mC.��I��'r����\�lQQ��#.NI��'c>��ňBd �ٕ�R5o��q�	�'�p�çĒ�}U8`������
�'<|2"b_�2h���ˉ�
މ+�'�(��`ݜw�0	�CU�*h�k	�'��1I++��ʦi����J�'f:l8����$� ��et=����'�I��J�F����0#bE(�'����&���|�@�	��'h\&���'�:� WN\F�ѩ��δ�t%@�'�D܋�,C�;�
��4�T�&�J�'u���=~�ɢ��e	�,��'h�P�Q�ѕk,ژ�!☛��	�'��U�������M��	 ��
�'U�<�%�k@�̑PdD(x(K
�'Hp�re��#��Ţ7�Aw�N@�	�'�*]�Qn��C���vX�*	�'U��z2F�F=����� ;l�^(�	�'kL���xVԁ�F�c�qK	�'�p��Y�*� 5gI݄):�z�'��]Ȕ���5���`��Rr�z���'n�ţ��M�~��v�ܽl|�C�'���Lۓ9:��+��a��`��'-����Mٌd`(�r��p]�t;�'���Xe@�?TD���%� 2�h$i�'V��'g�gRh��+�>+��T�'̬�7��" X��@�:5�P�'��!s��/����#��1t�t�	�'U
髑��F�h���Xa��DB�'�Y�gOM�I��q��ǸQ� �*	�'|$XӐ@#l��بFBB3�\uY�'P�0�QS,y�4mJ�@S�*Y�j	�'�
-�䥋�+��к���)�t4 �'�UR6c��t<��Qg�,x�'Z � @�G6=z,+�Ʋ��@9�'�V1�Da6=$��b�DE	�`d3�'�>c��5w�ʁ�B	#����'T�%�d �P�Tm*`&D�o����'���íHF؈�'N�
u�zS
�'`�9��"З�
<X���e�݃	�'�����N���ĹȀH�gg��"�'q�t�I��"pۗ/�g��,��'U���D	[�Gy��(��$�����'t@�NP.n�ع�������r�'!���D�r����L�!u��r�';����<mv�a D�Q<z����'\�\�g(\lT�YЅ\�[z�0�'���+V�ׯw�xh���|x�J��� l�0ALӰh)�9Sv��/h��s�"Op�eC��>�=`�cƀ�"�g"O`�#�Tq��L��R#`��Ub�"O�mZ0U����q$�P"O��Z[��Uq a�_p蕫�"O��A�C��"Rִr�c�&�l�ȓ+�9����%"T<	{�%Z���ȓ`��+�$�!�*Ѣt&M7�|!��oi��#�LU�J�H����h<e�ȓ#Y�����z2���q�`�ȓa��CS��EV�A��фC�&,�ȓ�q�0ҕ�Pp���a��ȓ^&��1
Y�A&��!'��E�L��ȓn��jp�H�
#B��j̩bU�!D���֢W�80�.�b��]@u�?D���f鏺ͺisc�ͨ1����?D�����>[>-��	�N��a%=D�����1nX���@F��F�ٱ�9D��qdV�U���H�A�0LQ��1D��i�O.:�Q��ÉV� ��#D�p�Î1Nz�5�2(�9n���@.!D�, C���R�(YcW�~8Y@P� D�xP�F��!1W � �����o=D��X�LA���/J*\jf=D�d���Ĭ8��$�AJ1xs>��s�5D���m�{�8R�)ԿO
p�aM2D��9�ӄAZ���1.*��5�����N���s� A�����S�2�.��$=�I�wGj�*����_���!�ް)�B�IjE"yv��e�A���0S��B�ɚ~e��1�F��K�V=��CV]� C�Y
�C'#qP�KT�d�B�Ʉ�r���::O�)c�P�"�B� !�F]��*�dͰ��g�A���B䉯3���u��TeA��T�3��B�ɤI
�|9��T[+\����v��C�I-om��t,ރ]$: �0��3;��C䉹t�F�ࡄ=z, 3(��)�<C�� 8���[*}���j�՜l��C�	/�@�7A�.^N����*5��C��2r�h�v�^9F��S�й�����>�Ҧ9ⶈ(��*{)�Y��%T� �@o���z%9b�d��J(D���	�wp<q�gձ#u��c'#�hO��K����m� 3GP=���\^�HB�t&�c�'	�`�x5�Y���"O0�PA�A&}xDD�;%p�z�"O�!"��ԙ$��Ӱ���^V�� "O�����K$�<|�f�z��۠"O������hwN�Ą�;i��@P"Oah!�C%:�̱��� }M4u�V"Or9 ѩW������O$B�XB�*Oʰ��)cb�Q'�_�G��9��'� �iGHD1Q�9	�oK�R���'�8�)���$G+�P�w�8v)(��'��)"�A���:���l��T(�'�&�p�C�?zq"l���b|�0S�'�Lٷ#�Js&]��hC���(�'=��j ��+f���ccNL^�5��u���{�wwH�b�Y�$Y6T�	R�����A�b� �0���	��^�F�(��9D��
���.PP�&�+Y�Հ��#D��p&@:���Ap���c
�Z�-!D�́&�(qX*����$�k8C�)� ��kS��>���eW#?n�1U"O �p�ե@�譲��Z���v"O��FW��6MX���
�x�v�'Bў"~#K	*a�FY`׹]����T�S�y�%���h������q]��>��G*|��Ir%B� D��U����D�<�j�1F !ed��%�����A@�<���l����j�� ����}�<�i?k�^��5��9VyPͪ0��z�<ɰ��2��Y��Z3T
���ō�v�<�d�ۀB���T�LwB`Y�]v�<飦@�#���u �y�@�qd�q�<Y3���4���)ҭ`3:LQ,�&�y�Cޫz4�6F��0�š!��3�yfP3O��1
�"���K���y��D";��b�ρ���jP*_��y�
�?X�x ���)!8�,8�i�/�y2�z�|9�6N���!�v����ybjY������1"�U6��<�y":r$���&:10f���y¡A
p��� ��M�4���y���f����v�D0{I��y�g���y���Yi���ઁuk�
S���yl�7I���FMתf�H��㜌�y�S1I� ��_u@�¬ث�yB�������E��Q?��X���yĐy�U�gρJ)x!�p���yRi���&�xF�7=g���Fe[.�y�O�0^�����_;�������y�%"�����	9�5�EF��yR���R���0oM*.��c�#N.�y��A7�z峖�	�!� p�/\��yJZ�u��q��0'�`0�
ٝ�y�a2Q��qj��O&�1I����yҋ��~O��E�+��m)Wa��yRgE�{�X1p��A,-a�Y2�]��y�+і@�U�u����&؋f�ã�y�M��6�9���~���0f���y��&�j0��H�.w~ �1A8�y�b��P�X���@��x�@i��y�	Qu�(��,ս��!X0h�
�yB�ȱRa���!��>_���B ��/�yb�ï�&���Z3�ǝ9m�BC�	i1hB��W;B�aǘYoC�	q4��k���� TnE$XB�I�v3X���f�_'�8�%�þs\B�	�1xL��dFX ~�z[Ԏ�%Qv�C�I+V�>��U�U)	�!�P�VN��C��:� `R$�K�C�^=����9,�C��<o�����%��͙#C��1ͬB�I;j�4]pv����� yu
")�lB�I
y����e�27*U��j��s��C�	�I�����V5+������'� p��lg>(�w`��$�}k�'��	9R)B�M"�wC��۪���'K����'��%�����l�@,��'�n����<��A',E0w���+�'.L`�2�O$� �DI��mAB��'3,���P8r�M�3U%`�����'�qI�WδIf@�9:Ի�'l����ޭgv�*�F��Ҍ4��'P`��틠(��`ŉA�:�+�'}�I��^�����%b��Y��'4�	�qDE���t���H��ē��� B�R�l�#y����]�b'��@�"O�@��,�,
\``c�<C2|�"O�9�%_1<�$M����!K[�)�"O��b�	�<d	��C�(zVX�*"OuaCB�ff�sIԞ2鐈��'W�'���'=�S؟`������I�dP� ��)-�8�j!/�6�����Ο��	럔�I͟���쟄�����IF�|�R�sI�KѵO&�9���O��Ob���O`���O����O����Oy�#�v&}���ԾI[�0� �O,���Ox���O��d�O.�$�O��d�O0E�Q`����P�a�Շ���v��Oh���O���O �$�O|�d�O����Ot(X�I���;�u�ɷG�:���'�B�'���'R�'��'�rA1K�	��oۉ�BdX���+T�'��'�2�'���'�B�'^�
�2T'Z�pthԡo�ē��U�<�"�'���'���'P��'"�'�bCY�5LVe($NHU"��=1?2�'��'g��'�B�'���'5�K�t4���B��1��,'B�'�B�'%�'b�'���'-��@'� \�"���@�pcȀ=�����ߴ�?����?a��?1���?a��s;n���C�0��J��
� �������?i��?!���?1��?����?����X
�᎘q��<���S�T	��?���?���?����?A��i>�'^�bL?#�NP���E�
B����<1�����xXܴX-TiӁi��I�E�,O�`<�͓��D��)�?q�\���	����*��Z��ųr�7ܬ��I韸J������'���?٥�B�#�',o(��3�9��
S���O��h�*�#�-C�2��x���.q[2|�p��r}�P�$��g��~]��w�R�+r�ՐQ���կ�]CV�Ӂ�''B=O��ŞJ��E�4�y��4N7<�#B%/E �}�ŀհ�y�3O ����^ў���ەc�7(�B��Z!�X�*�3-�Ļ<YL>y�)�O��q@#��Dņ�)7��2U�V��p@-�ɓ��$�O�dk��']ߜ,�Ŏ؎lqX1k�K�V��'����!��������W񟬠��'���8����2&>$৫�% 舨Z���'��9O�UE_6@�E�b�~=>����O���'7�I��M[��w�(�suc� ������,��4�'wR�'-"),ƛF����'#L�T�U�澅��Y��(1'�E�0&�,���D�'��'&��'���A��%�((Yg�S�|v��9P��"�O��d�O(��0�I�OL%���U�S,`C��t@!�H�r}��'��|���a@4&��I�E6=���x����k���Tm\�9��:��J2�'C�x%�Ԗ'�J-�A BG@ސ�!�%7k�S�1��I�����/K�dTr��Ei![��"oo�DX�4��'����?����?)���D@��ҳ��6I�������G���xܴ���^/Dnbe��O2�O��,�$�����%_$���	�yR�'S��+�T�#����ڙd��@�rU���	3���?��4��kf$p{�o�Y9H@ �0�*1�N>I��?ͧ~szE��4����pkSIʫ(��$��F-��"��A�>���J��䓼�D�O��$�O����	����L2k���ZbKX�`����O*ʓy�	ҟP����$�Oo2��#�M)n�p���)�=�T���O���'���'@ɧ�I�Q��ۂ	Y
C�ݺR��(��8e�13��i�H��|����'� ����<J��łΌ�����CN����	�D��Ɵb>%�'��7�� _Vф�K�Z@�g�P�`���O��F��9�?�6P��	<�H٪�M�մ������k��a�	�؁��ĦY�u'H�	����vybH� k��� LY�lm���p��y�V�����"!�>$���ݕ1鈑+��]�h��钫O�ʓ�?q��Toz��.�%]@��q��("��hH�}�B�$�Ol�O1� ���n���I�;^\4�V �I�4D�u�扵@�ؐhE�O&�O@��򤐉/����(�@��q�l�%xax2�>	(O����Y5���r��b�"a���,
�㟈��O����O&�Oh� "��W�az��2)�p���X��$[�%{Z�m�>��'9J��I�ts0k�*<m����5�pI3����p�	�����ߟ�G���'����CU�s�N��N-��$��'4등?!�v���4��Z�▊LEx� �,��bM)y'7O����O��d$"H�7M>?��k]CK����r�XƠD�/�8@+$J����'�L�����'/r�'-B�'�<l;��H�\z�K\>xe I9UZ�䱫O����O��)���O*��hIth@#�B�*D�b�C�O�$�OD�O1�@]�q�I�o�4�6e�+�b�RmB��6'?�1�L4<B��@�	Gy�|���!����\bg��z�b�'J��'�O+�ɞ����O&���BU�{�ֱkR�>u��D�G�O��oZ{�S�����h�	ğ��D/^'�n|#�Ϗ	�@��1
J93��mZ{~�O�8(�6�������� �t�)
1]^�X�,�6�&�I�6O`���O\�$�O��D�O�?��E��Cd�<9ebٚ!�" j�؟��	џD��O�)�OV�n�V�	l~P�x�J�d� pJ2��8�lb�p��`y�F?(훦��$���>B��		3f�}����g��
@=H�3��'f6�%���'f�'<��'�J��/�3IR�����A� !ks�'��U���O����On�$�|�S�ށF4Ý� ��iG�_Y~R&�>i�����i�?r�RT�3eZ�U:����X1d$��&,%\=�us�<ͧc�z�d8��C"
ui�$�"Q�"���D*w7�a����?���?��Ş���Ħ�HL
8k�f�P@ɖ)*Ia��m����͟8�ڴ��'����?��E�?ƀ�ѠЦ]��a�i��?�����Kݴ���φ�^0�O��I�C��ё�ܕ}��$CgC�Z�2�	_y��'r��'5��'�bP>�;A��I��ҳ�w<�Q4"�����O��D�OΓ������?I��X�q�=x������s��������'�b>������3�v�PbAɿX�.貓�ێ2X��͓%�������%������'�@���ғj��,!5瘽����'6��'drR�8�O����OZ�䒄|�j�� �[��ˑB	�x�<㟸R�O����O�O&@��Ļʒ(rq(D1R(n�"D�� Q���+0ތn����TVh��ğ�"�2���@# ����ύ�x�Iџ �I���G��wl)�B�B b�t�c`@�rY`q�R�'�L�����?�;.���C�8r) O�|�����?���?IC��M+�O�S��#���cO�<$-�V�U�>�� I��L�~s��O���|����?)��?Q�� 2,�ZO)c�Tͫ�o��s}��(O���'�b�'����M��\���R?C�����	�Q�M�'U���)��H��Ӈ��h�dI&��� �)�BH�"�ʓ"^ `R�O� I>Q*O�Y㲧�a^���T)���SQ'�O>�d�O����O�<i�R�8�ɴN0��:6]4�� O�E��D�ɚ�M��(�>9���?���]�ڬ�ԈbB2��TjN)���+�M�Ob�ӵ��������wN�`
8Xw1@���L�Na��'G��'���'&��'O�@�R��l6����Ź}�%��D�O����O*\�' �I�M�H>�.��R'O�2���{���gv$���	����!t[H�o�F~@]��ŚhG����T��d�OW<$�b��ɍ:��'��i>����p��B�ya3�ߔ^]�`;�lOE.����ܟl�'dt듻?����?�*���rc�,E��a�!�vby��0O��$�f}�'��O��O�(�BI�=���K.M!eAڥ�p�I�i.PhHᎊ9;Bʓ�:���O�@K>y��e&�(e@ь]���@�ڢ�?)���?����?�|�,O�eo��\�lL	1���XgB¼<�>�ITy�F|���4�O<�$ϒ&����&y%vͰ3j�2���O��� t���w�Jd۲�����O�� $k�M���� �ܟM�*쁘'������I�����p��w�TLD���H�19P�	�T��$�����O���v����4.J�3�.�%6�@Da��V�+���	H�ŞS�����4�y���=䴔jS�h�S IH��yRNˤ6~D)��:��'�	����ɶ^���"֥^h�yP"�!O��	��`�	ɟl�'����?���?)�*˄M�P �w���R�
5�͌��'���?�����L�f\��K��W���oІI "��'5��*dOC�=� lJ��t�ٟDJ��'���{�o�g���f�B?4�+/�?)���?Y���?�����O��c����\��"��Әmǀ�S
�O�Y�'��	$�M��w$���֯�X�@��'�	~�'���'~���9�����I�C_��
8}vtx�v�KE'�1ss!&~t�'�$���d�'{�'���'Kb�{@��(��Z5�V�f�,��QU�T�O<��?	��D��JV���O˯M¼#7휶@���?Y����Şs�]�cҌH�ԙ�Sg�)] L0[���0v02��'�@�a���ğLJ�|�S�x9JM<L�����Ν@�n-��lVşx�I����˟��oy� �>���{�=���^A𥹂c��JM���{���dBB}r�'��'�&��`�I�W���(���R�ҥف��ٛV��TJwdG%I�Q>y�ݳ\��t���=p	y�?e�>�	�����֟l������	R��p�(��s�ͳDI��A����L�#���?)��/Y�i>��I��M�J>	��L�\㲙b�3T�$,��Eߵ���?���|!�M��O �9�Kϑ_�84S����´_����'��'n�	�����͟|�	]�x���֣^>.��b�j�~u�	֟��'~�듭?a��?a*�*4��$ւsI�Hi�Ƙ�D��1e��D��Od���Or�O�Ӻt�B�b���0
0�h 1c��9��UA�93H�����S?W��?�$��Yz5#7#��b�y�*�LT���O����O���I�<���i�dP- g���*D��1��y�'��	?�M����>	�+L�ҩ��	�
�!D(�=�2 ���?����M��O�t�e�C��J?� �`j"�V�m���;aGKP��� 1Ob˓�?���?���?������=t��H��C�X ��ǌCl�'��'2����'�b6=�r�S�cP3���"��1�)�g,�O�$,��i׬L>�7�c���q�P#>��(rf�2Y]Z�D�c�0���
"cr�H�Jy�ObC˙��Yĩ.���@��Y��'���'��I���$�O���O*���G�0xp��U�֠M���D*#�I����Op��6�Ę4�B�����({*@d�+K��_��rU
"\"9&?�b%�'V"�	1�@ X�ΏS�ܡ�fQ<����ן��Iȟ<��J�O~B�0J�v�Ȱ��e	��t��7�rh�>a(O@�m�a�Ӽ��S�NI�����-o>lՂ6�D�<����?��_�p�9ش����{��	�O����b*��c
�A9��[���T�ty"�'���'���'{b�Vj3���t�D�"�9b���$�O����O�����Ef?$��1C�r��&�<�M�',��'Pɧ�O�lc"/b�U `H��q@
]��e_ "�O��C���?ADh,��<�'#M/��j3o؞E�Lbd!�<�?����?���?�'���m}"�'����p�܂HJ�(v	��.p���'H�7 �	�����O �?R��8�C�;�d�����s��a2���M;�O��R�����'�I���̛�n����F�F?M\��F1O����OD���O����O��?1�R�ܹ<r��ś�iv���Bҟ��I؟��O�)�O�n�}�	�x�y�!B-L��!7 7D���&�h�	��aQ�tnD~kA�x}	��k�v��e	�w�:��E��V?�M>�/O`�d�O���Oh�J�/~���F�f�j!���O.��<!�_�T���p��m��O�>V�L��-ĺ6�@E�FD����$�H}B�'\"�|ʟ�)Kʔ6t���"�$�H��Ā�����z��i>);r�'���'�<��O�Y[>�`����aq���V�[�����ޟ����b>9�'��6٫(b��烄qf۶$N���O:������?�Q\���I�1�e��c��/��1�hͻzm�T�'w	�d�i��	
f��r�O�֜�'�
��w�G�������(�5+�'R�	ן��	� �I��	R�t
H�m���7���V�E�1�D> ����?����?!M~Γ;$��w��-+���c�z,Zժ	$A��|�w�'k��|���Ƭ���2Ot2�Ь3�d���,%v�B>O
ͺ�n���?a�!�Ĥ<ͧ�?Ib��:h��07j)�FJ�dձ�?��?9���$V}R�'_2�'@�r� � �����=FL����Di}�'��|�'��Bo�ĸ֎ʴ/�В,�����A@����\.T1�l���T��H�"y�YŃS�:FmP�L oI�D�O����OP��+��S�(�Z����3�?+�
�H�H���?	�Z�H�'n7�0�i�9c6�Õp���!`�JC��Hp�dj�\�	~y�!�%�V�� 0��N�d�C�%��I��I�����}�, %��'AR�'\r�'X��'�z�w��?��б��Vv���_�У�O����O���8�9Or���Ͳe#���5�M�4-n#�{}��'2�|����C%1�^�!ĉX��//D�x���U���_>v�J�*��1>��ON�F��؈��]�a|5kp�՚3ˎ�$�I���I՟�~yb�>A��A�4���B�g��}p�20$Y�v^���W}��'���;P���2�P:F���[�K�ZL '+��q�'0.MkрN�?�2ԕ�$�w������eʖ\�T�e��Eڟ'�B�'�r�'�B�'��|5�'a^8"�n ( �S��ŮQ�p�b�';���>�-O�)l�k�ɰ2PR�!����蓷�T�G�'���I���S*2k�m�i~��� ܻ��ÈL���C��Jw� ��/�����t�|�_����������z!��eM-{�*H�vkZ��P�����IuyB��>����?����)[�M�V�f�����XYv�>a��I����O��d4��?�hv#^� 0�r����e��f�	*r*�妵��Ĉi?YH>a�J�@��݀R1|�T\�P����?����?���?�|�.O�4n�b�������nR~ٛ!kY9b=�	��d�ɇ�M#��o�>q��`���P�ʈ��IQ$�M��i	��?1rA��M#�O�������i���Tb$�q��[��ܹ��B�s���<y��?���?���?Q(����S�,C2	 ���Q&`�g}2�'��'��(mzޙ���5Z���Ȑ�hUΥ��+����Ij�)�-��io��<y����	�N=z0o��A��u�VH	�<����#���f��Fy��'�re 2?ڶ R�,+��5�&�J�F��'�B�'\剮����O���O���A�N��ay�%D�^ш���!�	�����O��$��˚<�\H��		H`��C�+F��:*B���͋�W<8c>����'68q��)g���&B:)�VL��b�0��	ß���ݟ���`�O�R�!O��3͏�P��{�/�+Y>BG�>���?���i~�O�.
[ȐĨ�K�.���s�C���O��d�O`A�s�$�}��p[��?� ����EA<,D<��G�W<��)�(���<�'�?i��?���?�5J7c����P��*\���B�ď��Ea}��'���'�O��m�Q`jIb�מE[&@�U�>���?�����ŞS�F5;�N�Z�MJ�
�p��U�"��M{�O�zW��~|�R��k�'P'n<U��((� �JԧD����ߟ��	���syr�>q�PTI�4/T�T��J߄�
 ��<�����|}��'���'~� 0��b���
u�^�H�a6���d�����#u��<Q>i���蝙�� -�:-J6���X�ٟ\�����������T�'O9�)Ib�W�6����ˇ3D�����?1��&���gy��fӔ�Oj���N��ؚ�&2t�h�z�O����O�L	c��6-6?���Hΰ��g�U	K���1*7�����l��L$�|�����'F��'��<�4`b͐��Ŭ�6~�� +��'&bX�R�OJ�$�O��d�|�cg<.	$$VM�y���{�iu~b�>y���?�J>�O�)�u�[#@ `ugӧqW��[�.�/XZf�R�B���4��Ȓ� v�O�m����*7x>��#��7o��P%�Oh���O��D�O1�<�qk����(nd�A���9yx�h��A��ģ<���i�O��'����1M���Ԍ&|8�Y���4
��'�jc�i1��7��%��?�����
�
�@�e� 㕂9H�Hs�4OJ��?���?Y��?�����W�����	��D>dt��#D'm,���'Jb�'-2���'�>7=���2H4��A̂�	���0���OT�d1�󉚛��6ml���CְY^����f�(Z�=�Als��倈�omŞC�	My�O��N�*Ju���U�(D4\s�DH.D��'���'|�I���d�O����O�D�4.�$�p��=������(�I���$�O���*��� 4���r�ڄ Jؓ��/p����	@�R�S^�b>��'༰�I�Dr60��lX��򂋓�jZ�t�Iퟠ��⟘�	~��y��<3н�*�.�̸z$L��&b �>�-O��m�@�Ӽ��ýdޡ���ƐJ�=)f���<I���?���P*�0ݴ����8vO��C��
�4��A��vcr��!3dL0��d#���<ͧ�?q��?����?����E�����d�|h0HA�J���d�_}�^��	f�'5�:��&�T- �	�t/,ȁr�Y� �����$�b>��#��9�,�f���H�aE5,$�l����D�,+�e�'J�'�剺O���Is��c��4��88�t��ן������i>	�'�d��?�@��}����JJ�)���R���?���i��O�9�'3��'b�Ǳ*>(-9�d� ~���%,�->4���i�ɰx����1ܟ��`��/vT�k�[���[Dʖ	6x�d�O6�$�O����O���=���>��6e]�2g��:���	۟��	/��4������&���T�ܔS��ś��MN�^��Qj�Y�I˟��i>���	W���'n0E2'Y�漪���96��N4O���I�z��'M�i>	�I��I�h?Ҙ�CU1"evH���n�t�Iڟ��'a�듶?����?�*�|��q	�4<
�KL���s#���z�Or��/�)R� RH���:! ��yz�Mj�Oŏ
Ne��)/3:P�-O�&�?�@I�O$��O����N��pq��R�|nD��ai�O����O��$�O1�F�~��&���_��v#��^�@�͂!�y��'4�aqӴ�Ol�D�b}"�'^��dN�+'���@x> �1��'��g 1K��2O���0ZWP���'��	w�X��PY�� {�eI5���	}y��'`��'���'��P>�&%խ(0Ąx��G�H\��������O��Ob����Ǧ�]4E-� ��ܼ.N| [�o�#:�0D�	q�S�'Œ�`�4�y�/Am��u����I�.��sd�%�y��ߚ[)�m�	�>�'+��ß ��<s�0q�����X$��wcO-}։�Iٟ��I����'T@��?9���?��o�z�~Pb�-�	��Y�gK�����?-����OX�����/���� #Mi���"�c�0�ɨ"dY�)�,,�ɗ'��d%I�H ��'M�҂H�'�09�)i�zT2f�'��'��'-�>%�	*'� #��&Mc�˰�C�kz��I����<aB�i�O��� ����$�O+{0��c��@A�$�Oz���Or��Ae���O�R,����V�u��0Ck��
�XR#E�R��%�T���4�'J2�'r�'v�k4�X�E�\- �a�
vG<-��R� �O��d�O0�d?�)�O�K���,��/D�b��0KVq}��'���|��T�N��H�z���)w��Z��þ.V���i��	��b�P��O��OBʓ@�l� ��)b�X��'ǀ1� �s.O�$�OX�4���DI����tP"�/<ZyJd�H'B`@`Ox�D�۴��'��꓎?����?���٠��Ȁ`ȴ%�.�&��6�L�۴��d�Q��mz����R����c�F���lE�f���;O����O ���O���O0�?E0U%ІU�,0��X���qy�MIşd�Iß��O��8�M#O>�u�Q�ZfM��O�kO�5��(K̓�?�+O��V7m(?�uEW~�? <(�gB��S�BD�B��b�$"��?�-���<I���?���y��δ��� �ۮ%l��a���?����d�A}��'#r�'&��~Ԉ���T�	�J��B�CZ�n��I����	Z�)�ҌI<����p��Q��!�	�(-�8ģ� �(7,���4F]��p�w�|"�\��|i��B�%���#��Å y2�'�B�'���[�L��4@c�)f�\ _6Xʕƕp�̓�?��+k���DVZ}�'���rl�g��"�m�j@4��'���ה`�����8�g�u�q�`� �@@V>�C�	_"/1v���7Oʓ�?���?i��?�����	\1�dM�S-�	�
tZ��A���':2�'$��'�86=��`3��[8e�P�-�;N���b�O:��,�󩏈u�6�~��!F�3YfQE)Z 1�(X`"e�09�fƓU�r��E�Ry�O1"+�3s�<V8���A`[�Vs�	�I� ��̟��'�\ꓘ?I��?A𢆝!iz���
[�K���:c�G���'�hꓑ?�����9N���6�D����2�۾,���'3L��U�W5KEX4{��D���{%�'���A�Mļ���/�"1��X3E�';��'�B�'��>���7g6�k�n�2�(�����,TW�H�I����<���i��O��b�	k��&x�T)PY� f�$�OX���O��#S&fӰ�+U������	`!��x�cjE�~�	�h؊�䓇�4�J�$�O<��Oz��nLn�I�cQKL,r���2J��|�IIy��'2�5�3��6�H���*��Q��c}R�'-�|��$!ʎAK�|��G��\�fL�F�ܚi�Z�
S�iN�I1rE�b1�O�O˓I내��8%�*�1����DѺ���?!���?9��|)O�(�'����͢�&gޯ ʴ�p K��yBbj��� ��O����O���B���YE�'J��3�/ҰS:���u��I��L����EN~��;>J|\:⦚�"��`z7D `�,t��?i���?A��?q+O1��8Ŧ�$��)�t�\�N�Н tf�O����O��ק���'�7�:�D�
"`k��[*t��t��:N`4�O"��O�ɏ�3�7�(?��CG�p�ڐ��B����TH0p�:ǫ�&������'��'h�qh�-R2N�hQkwgϱ6~��t�'�[�x�O�˓�?�)�h��bF�	8�e����15��#���<بO����On�O�S38���B�Y>o���ՀI9�T<����}q�Sf2?�'_�0��ͤ��yN�Q�(̽E���__�R���?����?��S�'��D�ߦ����u�x�CЦ8qY �ir����ǟ̙۴��'����?�pd�/PR��R#��v�i�B�"�?�����۴��$ �t`��(�O%��"���1��%Lc��X#ȇ2h��IOyR�'�B�'��'R]>51W_�?7��Rԩ�:jX(�c�
��D�O����O�����ܦ���Ċ1�ď&�*̠�'׷+\��I���$�b>]� B��ϓ=�]@�D�.�k��J�5+�Y̓dA�t	񢾟�$���'#��'ݔ��e�B0}?���	�S�����'c2�'��Y�H9�O~�d�O��č�T��4 *a��wFG�6���x��O��>��'hl�q���8N$�8P��\�/n��q�$P�1`տv_֜�N~���Oܜ���P���7"%U�L���H�i^�����?����?!���h�J�䊯q[��� �d�ڱQ�B4Ѵ�D�v}��'2�w����+x�I��A�$U��ǅ^�$�ğd���8:����a�u7�ǀ_���O�1O�`C�mV�@� �R�dD_R<&�Ė'���'d�'��'<��{d�� ����F))y��a��W�XZ�OP�d�O��5�S�l�MZea�	���qD���J6�tۮO����O�O1���觌߽C��h¡��>Qm�ə&�Ua�T7�BMy�M�$Q�x�����DY�,8h��'K'H9�4�©��3(4���O6���O��4��˓}���̳��8-��E����.s I�f���4��4��'���?�,O�5�2N�rQĹ��!�U�r�щ�`�j7m1?���B'eO��	\����)ضe���#)v!�#��
���?���?A��?����O� \ѷ@��3l�}{��Q���{��'r�'���|R�D��ƞ|r��w�h����-&z%+F�O�'f����� <����A��ݔ^�&ݛ5$ѕ+����3N&d���O��O���|j���?i�)��͊'�U�<UK�CŶsd�)��?�-O���'���'�2^>�@�G���܁��Muj���K.?�$_���I��$��''������}�5X�
K���-�p"�*u��y5k�u~�O�J]�I�k
�'�ɺ�xd�Y�{�|���'��'����O=�		�M���Ȍ}J�ja��.+�(8��H�<����?�e�ia�O���'_B@�a�7�Q�@�x���J�E��	�$w��o�H~����q�q�S|��7@}�+7�HnA�9�k^�3���Ipy��'[��'�b�''"S>iB�o	�<4�	��_�^k����*����<Q��䧣?6��yG�F�h��9K+[p��7Ě�,��'�ɧ�O���ه�i��� |��@�l��lF�a�3O$i7�^��?! 1���<ͧ�?i�f	�T� {��)
u�C ��?���?�����dK}R�'���' U@�)�%Ֆ�Z�̚i�BA[f�$�h}��'U�Op�SA��I�����F�O�� �`1ń͜R�P$�Q�|�ӟS��X��"��tX�d���X�*������������Iޟ�F���'�B���	N� C~I��6�E��'�����$�Ȧ��?�;_-�<2T�-(�E)v�P����?����?�tnP��M��O����fD�����h
�e��LϟNJ���\�T��OF��|r��?I���?���_�zP��їs"�i���*2����,O�I�'g�	ß�'?}�	�dZX3'��j����)�9M*���OL��OޓO1�
���/E2G�D�A��8DZ�=sf����$#4��X{�ϔ�!�h�B��byR�H"r_��Y� ��(���B�e*�2�'T�'�OI�	(����Obx�kֶY}���1c�#/��HzC7O�do���_�����I͟� �\#E#�+p 	2� ��勌sIo�O~�C�;2<
��SJ�'��3�g߰Wt���N�6OT,��	��<q���?���?��?9����ߐ_�>��͝
dnz��2�D����'����>�'�?���i_�'� TR��ߢ(��U���!����yR�'o��d��m�Y~2�(E�Qz%V�}2���0+!GX���\�pڷ�|�T�����X��۟��w��4:���b����TZ$�ɟ���[yBj�>����?i���)J�LS�Lq�_+5�q
󯂟 �Ɇ����Ob��'�p��BE�#4�(���<l�ށz��Q�s�lT3A�	���4�إ���%��O>�r���h�y8���: �0s�'�Ot�$�OZ�$�O1�n�W���O=T����m! �DdWO���y�Z��4��'�Dꓼ?y��J�q����%,R:B�kW���?	�}���۴����~�#��+-OB$�U�3�Ź�Å�'��� 6OR˓�?9��?����?������s_�#��"f`�H3��(Dla�'�"�'�����'t�6=��C'���|1��o��Vj���(�OZ�D7��)�`W�6Mj�� �%�2T�J
g�\�7�����d� C��%ps��I�Iey�Os"�S�S0T�6+N!A@9t�ҚB�'���'�I��D�O���OJ�G��	��ϰ'��xuJ$�� ���O��D/�d�jJd�c�.�3.;r�8�g\�PP��gv��v�ˡ~�M$?ݳ�'�i�I&d����&ݦP$��y�	#���	ן��	ԟ���[�OHR�f�2��Ds���Q/4���VJ}W����4���y�fW�]��8`Ai��J�A�����yR�'T��'	0���ia�i�)ҳ���?��E�R=w�Lع��]E��i��I��'��	�Iȟ\�	����	�o(�x��� @KB�^aZ���'J��?y���?�K~j�ð������	G&V �z� \��I���$�b>����"p& 9"(V�0�l�T�Hi�.�o�r~�aҎ"T�Y������=a&&1�lO*��͙⥔2J�$�Ov�D�O��4�˓uC��Ο��L�%Yb�M��l�-f�<�Z��_�����4��'�d듛?�)O�L ��W$C�4�F)߸h�p� �n�7-.?�aQ-��i�*��'��{���-&:,@Z�I�V���1K��<i��?��?	��?)��4g߳ a�2�@�V(~m��Kʗow�' ��>�O�6-#���*6+<(a�נp�:�ZAn i1O:�d�<��Q4�MS�OX�Ҳ�ˊNf0ˀ��Jwp��2�P�b����X�O�ʓ�?���?���8�T��#&˅K�R�%-ǞO��#��?	,O\��'12�'�2Y>ݩ�)2A��:뗪I.U�Q/?IRZ����ş('��W}�
b��6��j4��%�\mq�'��|w��+ڴ.��i>��3�O�O`L������ C���p���g��O��D�O���O1��ʓ c�F ޳9�8�P�C�2Zx�s���y��'���e�f��h�O�����B1��Ѩ�Hk���<�<˓-.P�)�4��T����'��˓J��0�c�b9��&hW
^�@����d�O����O����O:���|Z�K�l �([AoE�$RE�&G�6-��	ʟ������%?��I�Mϻ)��i���
��q���G� %�@k���?�H>�|���MS�'�kTlR����f�˞@ʹ9�'�&-I��o?	J>�.O�	�O�!�amT g��Q�쉧
(&ԋE.�O`���O��Ĩ<	[�`�Iџ(�I2A�XZp+k�TL��F$��1�?�CS���	S���*��W*M�����	��7�±�'����|�����D�X֟���'�d}��e�;t@)���b�@I��'u��'C��'��>U�	'��㔺�:��e�Д�` �'�X듩?A�<�6�4�Xq����Lȶ��ġۛl��u#�0O�d�O���G�7m.?��&S'd���ӣB�j!в��.?LS�B�:��'��'��'���'���'0�!s�D�78���G�!*^�p��Q�$ȯO��$�O��D&�i�O��� �9O�V�2��J!N܄h��x}��'6b�|������� j��v.T�B��B7���kp���m{�z�V����涟�&�ܔ'iҥ�lJ�]恢QO�-"`Af�'���'����^��S�O�����N�|�[VD$NezZ��,�u�'Q�7-?�I-����O ʓ9|�勘��b��_�L�ڑ"D��Mc�O~���*τ�
f�.����ErŠ��n3�@Ч��#;5|�A<O����O�$�O�d�O�?%��Q	?)�p)a.E� �m`��	ӟ��	ԟ��O��\'�F�|X y~�㮚�A"ؽH���C�'b����dEU6����� L�
QRl��fM�2�����eob�e�O(�O|ʓ�?��?��G���pT&�x+�m��@��?)Ox4�'>�'��P>��QII1!tԍ�dY��X�҂8?9W�h��C�S��	Oy:=��,ܗ4����0�0^��l�',�*��i�5]�擲!f�e�f�I13���P,J{[������r)��ڟ���̟ �)��HyB�j�X���,��Ku���Ժ@��02v:O*�d�O��o�X��V��	۟\�V��C���*��26*�4C���Uy�oU��۴���աKMz����E
�U��ea��u8���	*��+��E�d��@�|�1�$O�z��u����Ukd�hV�^ؤ
��]��[Elļr� �b�B�>�0�$!u�84�6n�cX��0� V+�""��w7B�Pt`�
�Z����(|=z��7�AS+h �/BVYb� ��k2$��c��
�8��U@�-���'9p:��˓����E��%B��!���UV��� �Ah���u�)h��%�Ι�ƌs�d�?	J�$[�%"_�6=a�g�'zR�j���D�O��D�OZX�'��ɞ59�Q��H,#�ryW%\5wN�	�41HBd��r�i�O�� �"D�F+t�Չ�9�Z���K��m������I˟�'��'��O˕ �j�k�'�k �!"�O5�M3L>�#�n؉O�r�'�2Ȁ)��ÖN�>�M�5`�H�6��O���t}�P����@�i��k��	ܕJe�ՙp�&к3H�>a�l�;���?���?N?-CRӬd\H���d��Px4�l�m�'��ܟ�&�x��ܟX0�"B6���H7k�'\��H��γ&D`'�4����L�IK��	����['��} C��NĄ�#�M#*O~��,���O|�D�,�ɳ=��C �U��Tt�'g¼�,��?���?Yd���%�~z��`ZH0��"D��,�!�5�XUc�i���|��'�ҭW�`��>�-U�9�(�s�'B?I�I���¦�����@�'�ĸ~���?1��D�*@2#
�
?�΁��U�+�����x2�'V�C�wa�O���~T*d��vM��@�њl�t7��<��� ����'Q����شD��i����HԒ5��@3�'�� jE�3�s��d�OZ����-��^ܧj�j}���5�hś�mɜZ�� nZ៌8۴�?y��?)��ud��RyB��\� ��^��	�to��@K���i�� 6�'��'���D @�P�*�"� &p�r#ET�H���nZϟ���ן���-���<��~R��<}�D���
�7o�aG].��'��}�|B�'�"�'��p��U h쩒c��c������w�<��O\4�'��Iڟ4$��ؘS���B�,u���'D-�L�@���H>���?�����S�cI8�h"���0��}S�.'P� 7-�G}�[����h��������f{���#�9N��&n��Xf�B�OC@���h�Iǟd&?aY�O�< �$-��{�耹�O��C�}�޴��$�OҒO���OVd�R-�������1r�q��㍗o��t@s��>����?��{��O�����J�Ǒ:4��l��c�����Ӧ�Ѧ9�	P�	y�O��~�6,T/�		fHȔ kE�_ΦM�	��'���#���Or����pyqJ�c���
g��9g���d�x^�t�����'?�iݍ�5�ۮ�
��ŀ3tv5{"�l�d��?���i��'�?��(��ɷ:��)q�'$��@®��+�P7�<!��?1���D���4���bfmB+cC:)��B�Pe�4�'D2�'XR�')RT��'4�ȥ ��0t7R�c��Lx}�	#Q�\@fM"�S�ORP`��IM>��	���'$�.���~�V���O
���O8�S�D�>iBG[�LH|�GM�X���p�K�>Y���)��d�'E��9C��!	T��e�!�f����'}�Q�\���x� � B4��AǄ�R�nJ���v����<���������8|F1*���j&���h�@˓�?y���'n�O��8vd
Z�Ȩ��R/V�|͚0�i8pѹ�y��'�	Ey"џ�����6U;���J����r��iJ"�'��OF�ĳ<�f��æ�8�@�<Fk�p*�ӇQ����M!�$�OL˓���|*��b,�h��B�Ș�'�x=���i��O&��<	u��n�	�k��Dx"cXc�dC�kU%��7M�O��D�<���"u�O����5v��U�F����؍3Bxis!!���M,Ol�d�O���O���� 뱃,
�>�3���c��@@_�T�'���''b�'��_�֝�/�r|4���=�>�7�A#�z7��O�V��GxJ|WO
��꤅	����H���I��MS���?9��?鄛x��� 6��BÙ\�$��޼u  �$�i�r�'���|ʟ��Ov����b�4��Ԧ�~��[�d�����p�	ǟLcN<�O���) W�%��-O�n`9�l̛��'��'���<!��?��� WT��"�Q��{RN6tɠ���iT2�'��7-�O����OD��y���O��g�0y����̟�[�t���iF2"���y�[����ş���p�i�v������*�?CL����fӞYm��d�Iğ<��7��ɴ<q��D����N

�f����;r�)�%� �<����?���?!����+��f�i�T���XB��!ѥ/�`���n�<�I៤��ڟ�'������4��)��jp�Tc�b�Y�A�dȔ��?Y��?I��?��82��'��+@�gL �r���3)�`����Y:��6��O����O���?�wȞ�|N�<����K�8*!��4/�j}�D�a�<���O&���O��H����4�I۟�2�O� B\԰��C^�F��Iee�M����d�O(�>����<��Ab��� ��80�(�UV8u'�r��˓�?���i��'�2�'8�Ӻ�� R��S�4����aHȦU�IԟX� hx�	����8B�6�[��5�]+�`P${A�7��O��o�ş�	П�	.���<)��?v�@Xё�� ~� �Ѩ)Z�v�C���$�<y����'��yA2B!
�@	�S8Ѡ4
n�|�D�O���O���'�Iğ ��X�t�F�Y\("A*U��-X嘜mZO�%%�z�)B���?����Y�#LZ�ln�����(�N@�i~��''V����Ohʓ�?��Y_��G�y:�z�jˋ	1�'��`�'Z�	͟d��aܧqZ�(Q�R�hr.YF�W�*��lZ����<Y����O~�D�O�d`U�g|�ap!���y;�/W�1O����O��$<�)��|:���&{�N�h c]}������Ʀ1�'�W�4���,�ɳ
7��i�i����{�H��7☟^bѨ"�u���d�O(���O&��?YF\?m�i�=��d͕?6�p�v'S.8�2�pr�P���<i���?I�iu��Γ��iĚ:��� eN�"'�J)ʂ�'U��\m�ٟ��	iyZ�M˕R?����,�I\v��5gڇV���3��J��O<���O��$�P4�D�O������ΓP��=Hfi�'��Ԫ �M��Ms*O���Ŧ���џ8�Iڟt��O�n��.�&���Q#G�<Z2����'���Ҍ�y���~Γ��O�hU��B�WQ|)r���,�޴�?�źi���'J��'E^�����38rDаb���-Г�Ky:��nZ�D�b��D'������$��$H�� zq �鑌��M{���?	���?�Z��'`��O:E�E\�"��sO�,i�$��Y���'9�L�O���OX�d�Ov��B�����y�6�7*�v�"B�̦u�I���O��?Y/O��Ʋ��E�B!٬���3F<h�P�t���e���	۟0��\��LyZw�
u��[��X y�@\))Ƥ�aݴ2���Py"�'v�П���ğ �d�χbRޝ��E�c�t�sc�#���?����?����4�Hͧ{����ħ:F�9�RO��;���lCy�'!�Iß��	�� ar�( ���	���'�: �i�(K	����O����OH8%>	��X��΄|e����C�_4T�(��P"XnZƟ�'��'�+[���D���r�8k���'Ik7�� R�oӌ���OFʓ�?��S?���͟����Ҁ8Eʟ>��X�᭑>�y�O����O���W�fw��uy�֟��k�&��]�^Aj�"֧)���S�i��	ݟ0ܴ�?!��?��:��i��s����*� $�%7�ts�rӌ���O��Ô3O.���<��ć[�1�:DҢ(��Axq;����M�'Y��'���'�bK�>�.OD���d� ��B1I��U8�� ���@U�9���OAH��A��Ii�`
��B̀�O|��$�O���O��'q�I��|�/�$�n݊>$�uJto�I���'��ɄRt��|���?����֩P�M ?��� �:�ȃp�i�b�'��듍���O��'�N�:V��is�Y�*�&�����Ʋ ����L�Iß���qyZw�5�g%d,�(��s�2t�ߴZ���Oy��'��ϟh�I��p9dc�")��L�0�O=2����<*���Idy��'���'��O��S�A���'�؎Q"ʍ�#&�<V�7��<�����O��D�O,)�c2O.��|�!��ۋ$�������}�I��h��ş<���D��~:�/|v�2a�ߗMHl4��ř�:����iG�X���	��I� #��'�~��W+�ց�t��%6Y�0	a"���M����?�,O��$SU���'M2�'a��8�NYJ�P�4�G#
����>Y��?q�P��͓��9O��8uw�1�  :�f�7a:a806ͮ<A��_���'~�'�rd�>�;�4�#�4�>t�"���K�X<l������,��I���9O8�>����M��]�֡B��	Gb�R������I����I�"O<��TݲI����t&���oM�b��M��i{ܴ���'U�'��*��T2�:3�r8B,C�7j�mn���	ȟ`�I��'yB�OF��%��(�T��tN
��2`���H:lX1O>���O��d�L�$���N1;.��pc�+!ԉo��T�ɛ��'t�|Z� .�ڣ�ݾt 0P��1��\�xj�eq���'~��'�b�~b����JD��F	5pU�xB兛��)I<Q���?iK>Y��?Q`���s�H
�I�[dh����&\�jt̓��D�OJ�D�OD����ΧZ;.��6�/|=<U�%��g��4�'���' �� ����dBB�۟DB���Ui�<%AϴY�0��7%4��D�O��D�O�	&>�M|��j��'ofD�fl�>���ڀ�d~���'��'���'$�M�W�'�cvF�1A�a�2��ڇi�um���P�IvyR�'˄�����Of �@�H{tm�asj�A1�U���	?�0��^�	Q�A_�L��#?��|a�%�Ϧ�'��k�^��O���'w��n�uR��W�S��I�Eo��P�I�Ǜӟ0&� �}JaM��6H{e*ñl��H���V��	��M#��?����?!"�xR�'l*���`�QX|�����5yph�Fm�̽Pr<O<�O�?��I�����B��H(:Qy��%���ڴ�?9���?���_P�O.�ĵ�������F5�� �S�rA�Q'hӞ�O�3��NP�ß���ӟ$mZ�*I�<�ҫ�� *����A�qW�F�'5�� �	՟�'���x>�hS���9=���aۢ@���/��������O����O��O�T�qc͘�dK~%H&'d�p�P�4Am�O��d2�$�O���D7<]���
H[G��*aD&�O�ʓ�?���?�J~Js4�H��a�!jwԜ+BF�1�UU�D���t&�@���(:al?�gG�
��!J�͆(?܆��!i�T}"�' �'b����&>,@�ݚd+�-,�Ơ�e�[�^ �4�hO�˓�?aJ���T�G _-��3猕�b�`��	N�t�U�v�B��A	Թb`�@��ĆR1������(M+ᅁZ�$T�cQ �x�F0-���C�N
E��2'�YK��rQ�ë����e\.g:19uM&�Vl*��Km�i"%��#Q368�F/��U(�,a��?`����v�*]�ڙ9������&��7yc�xrD*��}xl ���1|���U���}p�y�򄏩Y%��rAe1`�zā�[��:��'&L��ց��Q(``p���M����By	�Y4�ſZ� �R�A(�*�W&T>{�r���8ea��0n{8��ߴ�?���?�+O��gH@'�0�^�oVy�b��(o�Ɯy�O��a.kz1��'0݀�Y�n��(#w�ٍ6)��9w�߅�B��'��d Rb�q�g�ɘ+�fH�J�]��9��!��E�	M~��C.�?�'�hO6���l
/J,���؝R��誃"O�X(�	�"Q��1�_�������L���I�<ф�R���-	&��D���c� �d��2Q�i�2�'0�]� ���@ͧPc�� �K��]�æ��lC��*��W�w�����)� H��ϓ_�t�)�8J�IhE�ߣ-���Cw��z�"5���f�,��	�y�"�3cbI&R�P����
UH��`dJ�����IY�'f�OR��L��i�ԛ#��]e���E"O"��qJ�>ٮe@D�Z!\Nt8��d�^}�X�Tࡖ
���O� �r,-�h�aM��[JvA�'%�O�˓�?Y����nHu��+���e�>��1)g�D[�,>+ȹ���G>Q����d�J�r�!$'8�����O*q�ӕF���%@� �����I�MWT�$�O��`~�\���[#o��d�5N_%xr��<��1�$�4d "�b끆3a�����N	���K�|g�����P
H��$G��y�W�H��V�����OZ����$�.[TP]� �G�aP`co��B�B��O\� R�����(����T>i�O�!ȒK��4��HM#l��9AM��7"\�q��)rS�����- W�Ԃ�F�˕D�3b��q�E�>٧+I����u�O��)֜(�&<��:BٔKA�yB�\'����F��}��X�a��0<�V�C��@��8 ��4n�6��|a�O���OP�00�t�$�O���<�S8,0���*	�V\58�͓3��ʁ'�>1,�#[����|&�0�B��4���g��T.�� ׸$���[��;3&�1�q��'^lJ��#;��IcG�.� �p��'��	&]H�4�V�=9W�  ʓaݐ;�p��]�<�f˝B0�q��i�3F�v)!0dC~� ,�S��Q�<�0D[A@���W&;�B�fi@�^�By�ٴ�?i��?i-O&��O����;}�؀�Q��	�کU�Ήk�)� �������6��J!��#��A��T�PeP�b�?&���8�+<K����_Q����uK��b��tU�1{��'QZ�M�������O�ʓ��$�k����Xm+U��	y�!�D�6T�x�('*�M@<�(JW�`�0c� o�
�M�/O�I��[Ҧ��	���A����P$J�{�6��B�ԟ�'�2�'32��!@��p����d�;i��g��6e=�xp���n�xR�h}{�΍�xr&�ɷ��M��m"2B��C�J=���\u�|�(߿M>����^�ROr�'�7��OV+��e�q���4T~��֠�<I������ (�1RȚ�'��Ʉ�M�9נD SO�MmZ�<�H���6m8���JX�o�V���\��\y�ɠ�H�d�N�Hs����,SNC�ɂ)�L��U���-����锖(:"C�	6fEĕ��쎵R��4����aWC�ɝ0<]���K�_"N�� �C+��B�I�)� ���O_L�Ty���`=�B�	�u�:t3ӈșy��@7l���C��7d]~%��斲" N�I'ěC�\C�I:e��2R���mo��؏%EJC�	� � ��6q��8��(�C�ɄR��	����6���5&ZT�C�	�q�z��$��)�>�7�W�wFC�����A����|[`ǖ�`��B�ɶ]$<�:�k@2�1��$K2�B�I�OT ����ІP��(�耝�lB�]�f��Fl�;AN(�f:B�Iy~�剭h�LyÔB݌9{B�	S��3b�Y�j�#��� ��C�I�M;f�*���=D�j@ᓇ�.l5�C�I�4%�,2�՘ �d����/D�C�8�v�#ǑP6����N8&l�C�I�l�~,����++��o&b|�B䉃�`B�@('� c�-T'h�BB�ɾ2�,�b�ӇR~4�{���5R�B䉦0+(2�~<�AF��:t�C䉥�e`�I�p���x2�B#��B�	�&�(�HA�L�[�JD;c@��J�>C��,e�:U��L�.l�6�ɲ���|��C�ɸ
��qAA� %,x�W-_4�0C�ɝghT������E&wVjp��'X*I+V͛Dⅸ�� =U��'��d��X)�2��bR�1A�|�	�'D �cëx�L��Ro�x:>��	�'+�T0�����D��r�B4y�'�N`����&��}���)o֚���'��!F�s��\(�똊jkr%i�'?"eZub�:����U\����'�9�#�+��Y�֭�)G&X��'|�QD=�։�EΙ3�$�x�''.DHï��|~`E%M��Ja�
�'�h-���g6&��̇)~�`��'^,u̓"\rI	�ʘ�
�`��'|T8�ѩY�OK���QM�3��)c�'��uq�X�d�j ~��'Fp(rA�_Vօ�#/�M(i��'i`��c�
後��*[Kl�p�'Ҏ��f��=2l���=>��ى	�'�&��*G�6���1b�=�ѩ�'dX�X7e^7�꜒"�C�hl��s
�'g��X��˗1�&m�R�hͺT��'W���i:�O��fR�p�x�v*�+,��UA��'�������<�ǃ��l��ykg��"�q��@�<!�g�ru����\�;��Qc��y�'�c�<����;F�U�d���&��P$� +�"O��򭚠zA��:Ħ�!M��� p�I�*׺)����O�kv��'1����.��6��w"Oȭ�����#���]"b�4ݳp^�<1lN'�0>�!c�#e+d����/x��t90�\m�<��@�8~�;�BQ�dX�P����B�<i��s.P��ьDi�y��i�<is�Ϗ	= �:����,�LA�i�<��Љt��1h���3U�����c�<)Bi��=�y�� �
7=�AiY]�<� ����6V���d�5sT2-{S"O��u+)*�d�K���1�X�*!"O6!���H@G
13h©
�R�1"O��"ԍ�>m;�R#Q��s"O�6%uN *B �|�H��"O���/�:�иTa� W8i�d"O~�)�@C%nˠp���O�"	]��"OnŒԃ��EA�xZS�D4v��L��"O�\z�Lن4���Iql�9NF�|x�"Oʽ+��܇#��$̟Z6���"O��0!��o)�,Ib�Ʒ��R��O�|I�"�qb��A	D�H�wş��t����5?�!�']*	�fغ)c>���N5��r�'ڎ����,i��\��_�F��Ë�d�>������P���@J���0ySVsq�6u!򄌃q�T���GB,�A��-�:/��9D��^�|�	4zZ��6��|���28�L��ˆva��N5�x���x�Phb%���Ay��U��U�_�(5���_�9Z��Pp�'�`葅L��@Qr@�MZ���$ �򀂃�@��i�����ɒ�
8N<���ب-J
���E{�<��'E�UTƅ���Ф0!�I��BC~��]��RM���,F򥊰��X�O���W�ed�� j�'�(���'P� �nQ�#X-��D�-*�+ M+0m�4�'�J��&�ȓ��� 1O`��F*W6[Q�*OP$
Z<|2��'�<}0��),��x� ����q
��2�����	�S��x���`��+��'�y��n�H���VC��hE*%����F�;^d�Y�$��$˨Ԓ�$J�
����13h�� ܒJ��ptL� ��B�	��T�f*(z�n���)12�$]�(&"����8k~�8�+�U��)�S�o�xE����'β0����$9�Շ�=6�ٓ�Uit^�	��1m�$�7i��}Y\dϓ@ђQB�$���'���Ѥ�1B\ �M��X��9, ����([>%"׃�%�J})sG)_�&���C2��X�բķr���	�?�%{�&D<��WK�\%�G|�OB�$��A�� SrjaK���>�y�띾*��t�Q�]S�ؾ8���?sn��R.�k0 ae&!f)��Fmer��	2�R`��3�������k�*�i�W�lLB�ɾ��}���	!�4�K��Ŵ<&�i�Aɇn_�ΓD�ZM��k"�$����pY40�H�� ���	¥K�,��	|�d�h��gE&���A�N�t$q��52�F9yRl���dq� DW2g�Y!Ǔ#��yР�)`L�@���|�,�G~2�ޣF�N 1dBOH�)`��1�MC@�6-@�%LӾN��qS�/^$D4�CተZ��hIǬ!�~�	P#Y���ʓR�U�E/P�$1R-�'�F���0�)���`���*zF�����*P�B�	�YA�e�/V8*d8��ģZx�Q��J�+pb��FN�O@=��o,擃(��<�L]zGL�/�J�#� 	%'l��ɱ|HL\`J	�@bT�P��ѝxDT ƮV ��	 N�+U܋CL! l��$F�6x��m�Q� ؁͐Gax��(��8T�.,�9`��"[!Ġ�����h��'��'^Ơ�J<$���3!\2
���Q��nFa�/<?	#�4o�܍� #N�v�&�IBi��c?�I�\�
8�愚�Z% a�-D���$i�pÈ�@�K�$�D��cЯ�!	3�H>A��7ʠ(Qt�|*��xQ=6J\{2��(5m2���	�xA/}����7HG t��;��½]�b�K��ڪ:t�E�^�#9.���#&,O�D��͆�D���ᓅ=�}�'�'�>��/����}��%�zQ��A�%LkS�H;�,
�O�lP�Ml�<�gƫU2`�9Ю|9���cLd�'�b�� �l�O�t@[5��~Y�l�,"�(��'�������1y2`
�aԛJV�gfP�/j�'�$�)��<9�E��'"0�rR�h�/�I�<�A���G4� �*Ȋ*�F\$�[�<y0IC+ (����oէ��<a'�I9-�ja����GO����<x��WH����a���\�\.$�֙�!Q��3$�����@�Cײa�%I�y2B@[G��4K�MDx�nY�I�d�� Z�v{d����T�M�Ob�P��4E2�a�D�'9�b����� �]�O(^<�ڦ�@p���	�`�������)�� ���H���9�m�2�Obw�$� č8,f,� �"O�Q�n�^�4H�` ѲM��9*
ya��C�&I�!X����B��6�HO��a@�l `��IC?I*�5�t�'��HP5�A�C���2�M�
S�ѰEb�pk�h�� �uҔ��e���DT$��H��P�qe&�!S`=y��L�#g���(e���c�M�G��D�D�^2hZ�D�_��"I�g��yr#��n�8�?\�0��*�0�r�I�#Q�����S}��$�E�!��..���IVOA�:li���܈x�!�DTZ�~-��F�}��#ܒ^x�Γ석�S��x��,��~~,D|r蕰	��	ؠK��s�Н#��Ʌ��<�I�<%g��9C�K��2IY)V(��ς�����i[&yO�Ôj��|a~rۅ5r�$$�5 �qe�M��P� �sa�]!e��\Z'/́���|�ڇ1���Iĥn;x�r��T�(HxqOƭ��j��Jk,��!*q�r��Pj̺O+�����R?�B��O%�4j��Nc�ןh�:�'���*�ild-����E��2�O@���bA��@�2��� 5i\��`h��%���G :,��U�Jּ�' tBPa�z�	�w�*�
Tʚ,�
d��c�E���d]6�2��5럂K����PA�h6�3���<9��w'�bZT�b[��vkݟp0ay�S�E�v����t%�Tc�����'ժ0�>yM?Y�TfЪU�w
O�%�
u��R*o�Ԍ:�'�8���)ŏN�4��c/8>(�*��$$O���
ֶ���J PR�-2v���y��	!?b�%�Q�-Y�vm���*�y"��9)L�x�,Q�Z,>=�4�5�y�k�j�&��JB>Y5D<��.��y��n����0�^�J&�A)�y���e����Ċ>����d�2�y�%� m#��A�H(�D�z�1�yr��87 ��3 �T�R�~��F�8�y"e�s����2`ԩ\ ع27.��yD҃x���4��l�ʍ�V
���y�C_�ap�-S�`�ֹ���Y��y"�ZL⦬p��S��A&G^1�y�ܯU�h�%���[+�!�4ɑ�y��Q�kC�PѠdN�R�3d�
�y����v�vسĢQ%Pح�R����yǝ<�\Ah�JبH�6p�ݮ�yrCɊ?�h�x'��+=�bP����y�@�+*
uh����U��D���yb�C��Y�%�N(�!$�y��]�i`A� ���i�7�P� "O�u���˓ r}Е�57x�`��"O�hYfH��|���ܱJ�Ȍ�"O�Ժr�y����׊R#.c M�$"O
�����Y�����qV�,i�"OҸb�eU B�Jt9d�K�{4�x�v"Oq��
��g(�;)P#R"Oz��c"@��a�GU�aw^!�F"O�$���]<\�@!��D. I�\��"OZ\p��ڀy�A `�]����"OҐ��c�-��)\�ȩ�W"O�����4��#����#x�%+C"O� *`f�J�(D��S�M���U"O�51 ���"\�"�c�|Jp`c0"O����"I�nE��p8
��"Oޭ�鞋7����kB�<�l))g"O�}���ove��*²c�D�6"Ol��� �H3T7�(��̸""O�E�qM^66�ӓ�7r�0�Cb"O\V
T;3X�y�`6,���"O�Ԁ������ِ<̼� "O�թ%#^���`���J=;��aA"Or���K�+��c�g�|�8� �"O� v���|M����!� ��sS"O�,��O!���`̡,�0E!#"O5�eƂ���]r��փ����"O"�R�@�7*V��� S8\p�R0"O���q�I�a\ | .`!"OڐC�+&pĜ��K&G5�p��"Ot��h��ne�23�1J7�H6"O<���H� ��P)�G4A��-�T"O8�pÏ�f��9�F��,�b�a�"O<����u��e0"#ΣE�}A�"O�Q7`\<R��M"#޳嶨�5"O�	c��8	� \��KO�WB��y�"O>D	E��|p�q5��y(�jQ"O�M#��H
]�������!�"O�lk��:M����+V�J��(�4"O�d��E3<w
�o��c�����"O���A��4a8 ۓǪ/n���"OP�$�v(`���IټnN�x"O"AKBB�����ïPR(!C"OV�rR�584M[��6��\��"On��q��7��@3�\�[��"d"O�C��)uLq�я��y��� "O�� �Mĉ&Ex��22^(x"O 0��'�B�4��g�]��#C"O�q+v�K1T�8�b�Nv˰A�"O�ّ�ɞ�rF��J7l
�+'పt"O��ٗ,�*�n�J�
S&S�e9�"O��#e�\1�eZ�.�-K�"O�,sA�d�*i:b��Ar"O6���,�.w�b�p���8�� t"OD��J�#E�d�5@Y�a�(��"O,��e�Y<̬Hi��3-��s"O,(�ύ<=�h��G�V��8�w"OB��4�]:���a��R��i0�"O���$�5�L��R�n�&혢"O�<�7��(�nlP&�ʉx��y�"O��`�K�w\��C��A�~���"OP�u��XL���ǯ!C "O���D�J��Xz`$��t���' �I& ! C�E2!�ڑh�c�'�0@�K�(6�2�� �[�+,�iy�'�^���C�.G&�s�u�>`�	�'�p�!q��p���qė$q#����'��P�W�R����D�Gg"��'9��iG*�8x�����_}$�I�'�ZP	����*���*��-[�'g�(S��\�pa��� s*`1�'13&	0++��N�h��3i2D�ęF���6���pf_�2{
��@�0D�����Ӹ���@eڰP��#D��2�f��f���@$ �$��,D��E���BU#1�]�P��)j�m+D�li4g�yo���oN8�"Ā b*D�Tbql�"i���B��Sk�z�#5D���Y48��u����U�a@Q�����x�W�b��8q�eB�
��&���p?�O��@�7��<�@�̔(�!��"O����O���(���?
|8�v"O�n�4-� ��ږ�*E��M�v�<�[�(8f%��n-N�p�M�-|Ň�4���Ȑ�ϟo�v(�Tc�SA
0��4����c ma�Ç��N�Fфȓf�$l�m�K2�J`mЏ"rFu�ȓC�,��*�3e�1Z4c��pԇ�S�? `�z2%Y�D�Έq�	l5X��"OV����؁�0�� �	?f���9�"Oة��)P�,��l��!I�q��hRr"Ox�����W>RD�P��5M�`"O.Q�6cL�P���q�"ߞCƅ��"O����d�5�
�����*��"O4�I�뜎[8]�PwN�y�cM���OV�~�T��>f�B�F�D���Z�<��J��|���PgΝݬ���Z�<ad�J)�f �g����Q�e�`�<���S/���'8Kj�14g`�<���+���g�B0i� �zci`�<����%��50 ��,J�AYaQb�<����K� )aRa��GWh�1�v�<iG/^�S>�}:�B��W��0J)�n�'�ўʧ_x>Y��H|���z��J�w���ȓ`�b��w�ieĝ��a�
�b�ȓ>f:ECf���y�2l���)e��ȅ�q"�,Y���Ń^�,-�c�+D����-F�Y7�t���#��a+� )D�8�AYYO�� �A�`�TdDF#D�ܐ��"��	6�A�|ț��"D�P�QI5}Nh�@G�;e�@�@�>D��p���`�|U[Ʀ[")��d�!D�rGD���f�B����TY�(	C�?D�0{��H�Z�e�"Sи��@>D�`A��&s�8`��]���3� D��
u힡|la֬�o�1G�>D���'�� iPg� �^ �//D��铧�b	���*��X�@!$2D�v7��ѧ�|�F��	 z�@C䉞C�bt����2���W��.}�PB�	�!x��&��$���OJ;UTC����)�J�d|� ���C:n�ZB�	"�v�z��[��(���lC�	<`$�X:d�",���أi�H�VC�ii�E'R`@ۏ�:�1"OE�A2#G
u9�HƊwP�E�f"O$��a*��:�­c���;������O�O�V4rS���\@����E��'\�:$�ȄN�򌓅l���]k�'
n����Ts��[eK\P��Y�	�'vf�`r*�j�L�P��%G)�i�'������G��Y@���s�2�`�'�v4S"�P���`oC�"(]�
�'\4��g�,%�ܠї��3"�
<�'Q6%��BQ kND��F쟛�~u�'�d<QF���4nQ��ȶ��\B��-����6�4����+qr�q
�'�Q�-8[�F-�r�$  l:
�'ԐA[� "SԬ�r�H�n��P��'�~4��,�QrD<��j��8.M2�'��Z����K܂(Jg�
,*J�Ɉ
�'��Q�5���`L�I�㊐u�	�'T9�'`Ջh
Ζk�\��vF0��b ϡ"��S�e��0l��9J�Esw��
d^��殞�V$���`�0�W�I��!�q��%��цȓ�R)Q"��o�t R��;W,X�ȓU��(�CK-@|T��OJ�#���ȓ{�d���	�;����:+�H���	1. �ǞD�J�K��M��t��G�X��G�/S@�h�ү��p9����)?|-!�J�&W�
e�t'�6z`��S�? x�Bᔦl�ʙ`�E�!X�E:�"O��&鈮=��֣7AG���"O Q��Z�Y�9xd�֛X# ���"O��@h^� q��P���Ѥ"O525�F�s�20�F�$"لexD"O�p�6,��&ۘ�ҡ�ޥ&ц9`�"Ol�"��	����q.�a�'"O\����;�Ɛ�F$�w/l�JE"O���R-%b8�%Z���2+.�"O$4X��!`�d#�#�R1��"O� Y2��}�ą+va�\�B���"O�y�#��#1�T$�dӪ���$9\OR��@�P�:�~a��	 _U(�ڗ"O�K� fw�����iO��s"O��*�}(:%�-?��"O8 �/��b��}ydC�"��1�"Ol��ǜ��cw�Тl��0OJ�q1�W3"���@4\rt��w�<�"�ʎa�gE���A{���<if���9��-�Sl $fcX��#�{�<�!���*�r%ې���l�P�5�[�<!T)�~��غ э��!kfbY�<�-�;��� T�Z5F�L�<��k_:fD6�Q���.���� +�b�<�F,۝��5`D�?J�.���N_�<�#�$�N	E��`���R(@P�<i4�I5Bb�eju#�#J�B�	Pb�<�F&/$d�5)��|�*�By�<���	�R�<a4m��t��lzŢ\�<��.ͽ&��%0%�(g D"�n�B�<�c�H#�X;��U<U������Fz�<����,;Xe2C��zi����Zx�<��#9��dT���0�E0�_�<���FF����
~(Tx3#��Y�<��#M�^��x��c��-�h���	Y�<4�4<�M�p����mٱ�IQ�<	�O�FhZ��%cX�F��A� [J�<yI���rק����8��FD�<i�-�$SU���U�ʔ���~�<YTBT�cO\`��b� \���\b�<毁?)���Ս�w-�2�iN_�<�1�X ���#��69\>��3��Y�<�t��XL�"���R0S�Oj�<�S©v���'�1e7Rh!Ш�J�<'�G�w�`�­�0U��E� c�[�<�$/Ĝj���B@�k����J
T�<y�@\ ɰya�S�
����F�h�<��O�z+�H8E"����8l��y2,^9  @E�g��0���-��y��P�,�@]I/I�;Qf}`�P��y�ݮX�ո�b�7��=qR�Ԍ�y��Ԇ9�Ѕ����/'��!##-L�yB�
Dwx*���$4\h*��տ�y�!�.��H�#�1Ѐ�Cq�[��y��S94|h4�ōV�'Oz]� ���y"f]�.�x<B�K���pcQ$�y�e1D�eK�̕�H���J��yB@^�g�ܬzP �65�L��$�y'O.h%bU�cCõ�ٓ�o�)�y�OҮFf�9�t���r: � "�Ǟ�y��ҭ<��x;��k�\aV*Ǹ�y�@�>u�*ۤ��iδu�׊�y�i�>p�PЁ&
�_r�r��I�y�$ĝQߊ���f��r�ᄰ�y
� :8i�H�Aezu�D��6j���CP"O
t�ѣ
@l�Ӕ�o����"O̝���A�w��	�pH�g�-�"Odɐ���$+�ܰ�[�Bj��"O<�A�˕(�p8�&ր7���YP"O\{#��i\x�Ju��k�B�#""O�A c�B7Y���	z�<4�3"O�h� ��vy���	�\���"O�U[V
U� w=؂�I�B�t�x�"O^�� �5�X٠B�-q�%a�"O�Y���F�p8�H�e F*MwX�"Oj@c�fh�*2mOE`��"O����Z�j�*U�n��H*p���"O���@�.-�xMȃ��DV�R�"O�� �.�'<�X���=Nr��e"O�� WF��I��HB�&f�$hQ�"O �R��/9Xe*v�	A�x��"O,��K�.\�(	�a_k�(p�e"Oȁ��U5\�L���`�
tM���A"O4���&��1Rx�J�IO@n��"OȨ� �f;���b��0U3��d�<C��2���!��&\�hw��b�<��cN%B�ʍy�K��1V����]�<a歍 w��0�ܩ.� ����`�<A�)XsЂf�I ����T`�<)�B�5Yc\�5H�%#��@���\�<�AL;��f�#ˢ���Wd�<qd��?S?h�CP��-~�1��σ_�<���,@q�u�8c�K��m�|B�Imj�;���DA�̓�ޭ*�C䉨;��+���M�&���/��$MC�I,��#w&�^(6�@��=��B�I	q$F�1/�9�d9����%�B��4ExơX1.��3�պh[�C䉀��k0mB�f@�k��Ѡ`I�C�I "�Z)�����&� �g�(c�JC䉇ZI�`k��@2Z�H '�H��B�	%u(k �B,.�V(SĎ�#��B䉣5��@P��^�j��G���9VB�ɇVw���V-1{���t 5��C�A  �*O>X��I$YrC�IvlH���x��B�Nؕ^�>C��8,�B\	$���N���ԊY�,C�,��ً�%O	gFI�c���
�B�	�v��}0�e�	*�b�i�CIPL�C�ɳJHP�Խ{|B͊�T�T�FB�� TV�D&/�_�¥����7Yf<B�	6x��ߗ%M�=��ߋF�2B䉨~�6�cAaO�w
<!EߖJLVB�I�w<��q�$W�JuZ���
L�lC䉞NM��#�&��i�Mު "@C�	�41�9je)]?�����E�.Ac$C�	p0t���˓V���8vB�V�
C�	DII�N�|����[(%�B�ɋE��0R�F�8�Z!1����^D�B�	!m
�aV?"��A�/�FH�B��~*I�b�4�Qxǭ��s�TB䉮`o��d�J!�ҡc��� |@B�I �*�r�A�&nol����to�C�������^�k@����X�C䉼.�����(@ĳ䭔�f��C�2J�0��'%�F	қY��B䉆_6*�x�A�<z�,9[��)8�B�	
��р�R��0���ܵz0XB�)� Ni� �U�!14�y�f쀥"OT���%@�Ml)���àq�,m��"OL��ɜ# �l��u�T
l@4�w"O�a��cL�N������)4t���"OhӄFy����M��1x:8�a"O^���FM|z�t&D98�p�@"OD0"�
����D&آcʰ��"Oڐ4
 �m:��Ӥ�N��x�3"Ovm�Gh˽	����C�$��p�@"O�����N���]!���E��z@"O(�xE��`c8H�K9��`"O��WO�E�4�Rl=\��	�"O*�gmS'���� Y�~B
Xy`"Oʭ��섥js�`F��6)�ƁC"O��w�� 农H��G�~�0c"O9�D��(E
4�ŧ<}>.���"OP%x���!��)���j�,��R"O���$�	i�,��@d[	NuJ E"O��!k����]�p��6e�S�"O�X�å
_��'�̫8X�(r�"O�t�3�ft�"�P!,H�)"OT�Z�G�hVځ��V%z�2��"O$((��8I�H�Ղ�Z�ݫ�"O�ܙ"`����M��a���r��'"O���V&�9x� Aa�|���e"O5[aĕC��}�w�ސH���"OVے#Q�kƤi�CQOƌ@��"OJ��D�J�t��M�ub�'b�ě"O<�ڕ�ўiy����̊C�ΝSv"O�:�i�?9�1�gN�.s��q��"O���$��Y)pqr�v�V�yB"O��b^R(|�x�J�hlJ��!"OJ�@�C7d���N�d�2p	"O���P$�M�dw/�D�*���"O��eD�8x�����@>`0F`��"O�c�O��.�8��(!v��!"O�0�o�TȔ��0�I�	��B�"O�]�D�٘P��	��	3,(�=�"O\T��cGO�\�H���6�%�"O@�0*��:y�ihB�Z�a2ܔ �"O�l�s㊠C	���n�l �|(�"O�1��bԴ�6N"|� ��"O�Y�b�i�������Ij̱�"O�q��l��[O�����H��"O�p	�oHh̸9d��!W)f�"O�1�A�
[-�(���)rbH�"O�	�0h{'��9W`[N憄�c"O��UĻJ�h�� �Q?_�p,��"OL���ō��-;�=w�Phچ"Oj)���,s,@��m�u��%�#"O%A��X�^x�Ѧ��3�pUrs"O���"�:�j ��,�%S��"O8ɒ�.�?Eyb!J�ZmXeT"O�x��	7k+L-�"�R��,�7"Od�!䄊�T��i0�ћ]�N��b"OP��M�+�u8�(�~���B"Oe�Sh�ZID�CVH�8}rఓs"O�,�Ej�7j�q��!ųoEΕ�"O��K0 �(tD�,�a�N�Ua�HB"O
PA���$��" 3�X��r"O���E�.f%�=1��ݡS��I��"O���2(�n(ѣr��Baa"O��b�	)@��C��ʼi�"��"O|5a4���j��ʳAC�d�$#`"O� T��+�%Jm~}��aV#.�L���"O��A&e���ӯ�
���*"O�YS��2/�TY;Q�� (���ZQ"O
�h���!@f.YQf�?b�^��"O�̘3χ�E`Q�	��}g
���"OڬAw�Ft�u��¢	L@��"O�Ҷ΃}2L���G�ZK*��5"Oּ�e�#	�� ��Q/�L�1�"OZ4�%�O�@��� ����鐥"O�d{�eP9����M�����a"O"�ؤ��
<���8B�+pG� ��'-1O	0�I�}z��Ԁ�3e<�v"OB�Ȗ)I*G�<�S���*:�pT"O��I(j���G/��?}���"O�#iM-H�ڜ��	tq
\�u"OHy�O\�e��ɹ�׶`�J"O�Ձ�a�O�(��&I?6�.8 �"O����
[<w΅�H�#�T-�"O�J�ߌf�T3c��@ጥ�B"O�21��6&:ƭ�gEǣȲ��4�|r�)�[�$�pOW�+/l��O��.XB�4u-��1�]ڀ0��J��
^nB�	&� �ٖ&	�i:"��@��.2B��4)!���`Qu/�%�B]�`�=�Ó.��:@!� P�����M4JW����Rnn�x�NH�]ʨ�I�A2uZ����U��q2ՆʚG@�	��%)��m�ȓz���9�g)>lqQ���.�ȓG����j�����*�W����ȓnf�y����?e�
�ҷ�D�]�����1Kp!��W)��U�樜�x֚��F� �L�;�x �dm�-<�D{B�O�8�@������bX�ށ0�'��T�Q��.Kk�)�+�NhNJ(O����<!�a�@=RoBL���-G�!򄁧)`j	83Mķ@<v��V��$#!��,��-���
j�.��F�!�O02<C�/\�t��UC�F��,!�D��c-��PH�6���e�? �O����i.lZq��"�䲠e��!�$�(zd��B�.'�T�Ĥ[�/!�4#����@&$C�����(!�䔜_2 �Z�ZH�8@�Ň!�!�d��T���rʊ!!�6U�D��ii!�
�`&�l��	T� גi
S� �e!�$��K䔠��%�C�,���oF�!L|2\�G{BN�lj����*���PUK�;R!� 4zA���1�7�Z[7ў����e

U	�ɍ�!:a��d�t��C�		Y��	ʧCś�6ّCmB;|�,C�I=J�h��$-G�F��(	]�!�B�	'P�0�R��0?!��E's����:?��H�78p�a��k�4�5���[]y"�'u�X�Ȓ-df�q��� 
��)�'g�9s��Њ	���{�G(%�}�J>1���IY\g�q���ֿ/��!3��:S�!򤂡+�2M0Ġ�))�LD:E-��!�䟚O�
U�0i��^Ľ�E�КU�!򤄌2����+F���piБd�!��:,"8��ٶ2+D��怲0�!��]̆|����d!�l2&&�z�!�D�46�G� �,v4$�u����'*�Ob"<���PJȀPd��H=X8�R/�H�<���E�~҆YS��[Wn��(�ϖO�<� �]���ԤvTt)��eLR�8��"O2�k�l�+����bץG��p""O��3�ˡ�L(�U ��Q�_��G{���T��|�┮��s���Y6��=;�!��I�|��J����S�P$#�!�ήuD��2�>Hxm��.۱�!�FC��bG'�f� �UG\�C�!�DU!�hĘDi�)M��[2Ԝi%!�D\�v(:ASV�N�?�����?I!�n�I�L�$��22hY��!�d�%h���1�A�.�D8�[[�!�Zr����f\S��C�f�.�}��Jf�	.?��ӷ#��<�|�a�.D������(��mRD/�9n.j�D+D���%�Ӿ�\�!�K&7�D�{Ҥ(D��Z7GZ'r�l�ɋ�,���'�O��61���"��c��xG�
,T��L��G�n@�E�%�.���C�hް��?����~�5ɝh\�s���pQ�A�Wp����I�q|�#m�9�M��K�5�p���t<٠�C4l��eEL4��|IbOi�<1w��T�.�"�l�ZG��k��Y`�<�G�B�V���C��7_�Nh��]�<���d��2A�3L�j��$F�dh<i��BR�RD��FV\�z�r2����$)�O��� oH ����2���d� �"O$,��#�ET�@�aA"O���"E�9|�8�S�S#�94"OF$�v ؃CqV�J���-	��5"O�Ő� ݼ5%ִ{C�3�ܴXu"O�jU�B9����d$��E��� ��'�!�d޺u�BI(d�R��,M�EE��)�'q���F(ܤhLX�K�3��5����x���~��8cE�'r�H�hQ��y�h�1s��1jD9�>tʑ,�y��&Z�h�8%�"{ݠ��h��yRL�&N�̘Ѵ�֣s )h�͆�y�P�l2�E`D	fʬ�P2%���?Y�'^�y2P$�*��+I�$�>ؑ�'��d��BʭUZ���@M3 a�'���'�O�6���k؄v� :�'&j��&dG�(ۼ)�a"�	gjj�'�FpA�+��*����E"� Mh��y�'�b���#v��� ��25O�0��'�a�@-�"X�i�t��2;|����'p q%��MN$£�JkaZ�s��y��@s["!c���T�5�L����0>���J�*L�|�0o]"���"�NX�<�Vd14�>��WFZ������Q�<	RE8I{��y���n��
A*O�<��bG�9�Q�Q!��@�K_v�<�wC9R�P�!�<^�.���D�=�'|�J���
T)e��0 �'u��)����<�e��5��6N�/M��;7B�n���'�1���!w��'y�@eJʿ2�%�"O��8�B	E�M�*M%"�2u��"O�Q�D�2TʤcRi\�}��,Ƞ"O�պF�8���v�a�0��"O���@�%/rص���
�Dy Er�"O%�'�B�d�#��Yl}xF"Op��"M�m3h��[ jTT4�Q"O@+��6V��z�ܝ�@R�"O��ӄߑ9'�X��J�r��T"Oj���3,T�����X0U�N$��"O� �11r됟m/n�" CXu��M��"O��;q�͆Q.\�%J1b\��!T�'��'�B�s��&"O���'h�>^0�a
�'�(]c�)@�t(����Ӓ.�A

�'�`�z��(F��VF� ��Ո�'_\r��y��sF'Ը-�T��'�Tq��߅����ɨ6��1��'8=å �#��h��,��c� H���5OTxkf&�3�TS�Q*��	�D"O�9���L2��������"O�]���>]	t���@@�fD���/LOlEiwM�/I%h�U�nl>���"O��F'bV�s1�OU�Eq�"O�Ȥ*Z�?�dl[�㛵WT�ȋ�"O �Ñ2mp�_']N�0r[�<D{��	2b��@��'؊U�SC�#4!��0 �	�bmM;0�
m負�"?�џ�D��"c��!ª#���W������hOq��y$���O��Y�Ea-5:$��"O�@d�2tt�Y���ݒb/���3"O2��V"��$�������!/4i�A"O�9x��I6,r5@L�G ��J&�'E��y0�{���s�^*x�^��2�:D��!�/C�9�dK�o].IH��� 7D� ���U�}�5ۗ`�	����� D�`Є��(<?��h�IB@�s�&?D�0:�HS�IN���̖&h� ��p�9D�$r�\g��yTdӨ~����� 3D�L��o�2α�C�n���S6!/D�<�vFүs `��2h�(�� e�<I��0>i�Bְ2���y���}�R]J`l@�<��JٴMNZ|K��I�o�,��Ba�zyRX�&��g�D2]�z��D։��Yic�ά���F��,�2��uu�� �N��S�dt�4n1D�h@�%�T�P$I�BR�_bb8 �04����/�vҜ�'�X�F�$��×^�<�� 6�p%���ɟR�t��ݟ\�	[����"��C������=���
.D�L��F��JJ&_�}���:td�It��(���!�ޔȖ]���Ɠ��4a"O�y��,6[ ���$}➡��"OfD�EłxARD"�F7��h�"O�=�I�� �BHk7ŕ�u�4��"O|�䕄UR��(d<Y�b�"Of	�k1(**%D��"O@p�A�.�����33�� "On����|Y��Ď�.�ޭ:3"O�<�k��]��]�c�7��M��"O��Y��4D�(1����<��#�"O YS@��W���1��x�Py�"O��'�X3D�H���DhX��\� ��I%*�\���J ?	��u+�$	�p+`C�	r�������h������F^C�	K��=Љ\�Dږ�����o�2C�	�:� i�ʀU�|�#�F�X�fC�	�=Q������<,[�J&�DC�I�-LЅi�Vjr�0уo�j�B�I;WQ�Ȁ��C���G]	4=����O`���
C�(�$�� ;B@ ���6lL!�dKx>E�j ).d���!��W*�>��l�b��Y[0�;X�!��6`ZP�w�1\�b�0�a�!���"t2�x3"O�`��ѥp�!��Vl� ڢ�Ș3�HA`Q8U�!�� `��G���,%`i�Â��w�	"�"O� )����~�d�SÂN�.�4�s�"OvD!R@�Z_��R,�*��8p"O
ȋ�X�|� ��QF���dp��"O�S�*R�];��@@��XM����"O������!`�� ;I> )e��X�<1�LId�i��Cˎ$���g(LR�'9a�t��Z�Ш��O�_*.P�d $�y"c�}�����ŝ�PJ��e�!�y�Ny���Zd/�A $ȋ�c���y�N]�yT��sC"��<�����I��y2�����ɨjC�_���@�9�y�I#8�H�B3#��L��V����<��$��M�:U�JJ8_�AP�,��"H�y��ɷI�j$AVa�O�J8[a��Vv�B�ɣu2|bf��t\��ڸ�*C�ɷU:���I+h��U�ܿ"��&��DxB��v��P�&c�Zѓ6�א�y�KeP��̠\%BmHvP��y��#h�.͠�C�>A����� �y�i tn��{d.E,!�Z���-���;�S�O�f ��L[�'wv�j��4]b��
�'}�ԙ����I`�
Zc9S	�'ˬ ���S{�k�H	�L2	�'@�r�W��Z�
��X�nUN5��'6�bC�֞E��I���`����'{0$񷌏*
� ��l�>H�(����z��83�A�GȤ��*�#�y�0 �(A��$-1�\��M��yb���
�qxW��#qЄp�+���<!���׎6�2[��޲H�ɳN�Q7!�D�hNdX�E,�c��yD,^,!�d�;�z|Q��� n�^�S�J֕6!�D̒Z�i�ЀU�
����!!�A=l u�F��#��I�!��4#�!�׮d���ըU5o�u+���>A!�$Z�k/~��%�����}���ѹ����L�UU20�A���y2s�/+����?�I�����c�
�Gp�5a���16^&C��Ջ3�U1Њ(P�(�C�	�T����pO�#Nv��sl�>9*�C�	*��Y�$[1a�* #c� G=HB�I�"g|�[���ZN@�k�a�$v��B�; �Ƞ�՗_��9���)ȾB��2ef,t�NU�/T�R��[.��O���=]AB���jY�1 29�D�o�!��g��!96����`�zs��9�!�P�U���d�)�������.hw!�Rt� �"�?-�qPw�_�
�'�a|�k�'��t2l��^�-���&�y�啣,�D2C	��U+DA̙�y��Vt��	ÁS�D�k5HL��y"�4V���"[� �rpX�(�&�y�g���pZd�τ�x�(0j��y���,����C瞽-�i�b喬�y"B��S!�QH�;zوAE���y��Ķx^�u����4��T�'!��<'k�\�e����&�  !�G\Ґ]2QJĺ>���!�!<�'�ў�>����3\���b(ХC��K��2D��bw�P�He�q悆lD�7$2D��0��m��5�d ;hy0�% &D��@e�ͻ��z&k8s�.0{�%��0<���ݎ��0�,U2b].��"Wx�<� @ԁ��GA��Yz2�͙w�����'���H��-I�����m���O:D�@���RW�&� �!�.r
ƹI`�$D�H�f� �2eq����c���'�0D�`� ��=�N�)&e��ZH��E� D� �(�0O������	W�À�!D�����Ǫ`;H�y���9}�h�qB>D�H2(A�}���Sv�E�0��p;|Ob��01��wDT�� ��_z�Qr�n7�O��\���R��m�����pw��ȓi�(Ѩ�0B8F��v�ߓ\&��}�Kb�\0q�@��@Q:d���,��p��C1K��"#"	�X�l'����Ʉ/z����.T�����N�C�ɥa{(��F� ΒЉ�/��C��,�(��`��2a�ʽ{C�ŞqưC�I�r"r����g��m����K��B�	�m=���	��2i����)׵%�XB�	�D�Ǟ,Q�d��T �Fi��?���i�.��5(��� 2�)sl��fN"�)�������G�i�HTҗe�LW�T�
�'����Q��"��q��L�@iX���'�~H&i�uP�8��54�d���x��UjD-��,N�9�%	�G�2�yRș�e3\�[c,,����'�%�y�"T?_!�2���1/b��׫�y��H6H��1fg��"HR��Y�hO���$X�C���c��X�eyb���#b!���kR\bc��uP��:�d��:E!�ę��P���a<���%�[� Aџ�F��( �q(�q�F��N����ybI��R�~������f)�$F��yr�[�a�N�:5�N����#���y�B?�$�Z ��L����B)�y钄q��C�@��,��#��y®��YD�T�u�����j�%�y2��2Tf���5��8�T�;��1�yRb�,+�5�ԕg��l1ǫP��yD�^	4���HEZ��|
'�I�y���7z]�镡�$X��Kfk�&�y�!AR�<�T雮���x�H[��?)���{q�L�ĕ���(��X�2ޔ�ȓ3�H�as��:40U:�dG-\b>��/����w���<e -� &B ;|���ȓ2��a	��*3���a� G�l���'HX��jޡ��k��i�"�8�'���Aa��y�ؘ+�!ͬf�tj�'X��3���	����=�R��'������
}��x���L�$:1��'sv���+kA�yC�N�����'[,|�3�P*q�ZA�� J^l(s
�'���K���?�� 1!+M�%<��	�'?��� m�g��,Q�BË	�|
�'� ����S;9�`�zV�J�:��
�'�.�1!+l�J!FS�%ˀi�)O:��0=�a�2^�=�5넬���I��<Q��ۗ���i�.�%.��ųӀz�<qc�>^���s�@ �H(���qyr�'>F��`e�\���	;3XЧ"O�C4��0#�	 B!)�|�A�"O�� �,Hb5���"K���i"O���v�"?'\ѐf��Vz� 	��'K��1c`<("�A�&`�YW��N�RC䉫5T% �k�*a�F�SL+<�JC�)� �Q!���T� �(��A�a�|��"O��p'*Hd)@DM�"vr�"OԹ��I��3-�	jk�i���t�<�,�Gȥa���]3P�Z�Yq�<�4�$Fa��zs���N
�p����j�<)�Y�sxDHɇ�ԕ�m�5��f�<�Q�H=c@NȜSk��9�Z�<	��X�M��u�`gZY��q#FU�<a��6�0���oz��x��T�<�c��$>D4���
��E��ˀj�<���D1�|�2�ˮB[fqW�#T�Ly�'Ȏ
;XͣF�6�`hBf.�"�Oh8�D�7# `ecfϛ�(��	�"O��&�I�R�0��H*t�:��"Op�5�A�WI��",��Yzj�"O�Zr.^*<�̐��I#7d4=��"OB� Bd[y�< g��W�n`� "O�(��i\�9``��e���fi
�IC�O�$���C	
�@'
'S��):��4�S���z�x�7C�M�\1)���q2!�Ĕ�U�]�%LG�J�j8�F��B(!�$Y��1�`E�DE��?!�$�$Hc��K"��wB��1�L6Y!�+�I9��S�L�uK1<
!��$rH��D���̓ 
�>:�!���Fo���BJ.Ԯ����)hx!򤁮F#�H�A%uþ�q T`!�Z�����Tl��T����eN�-n�!�DN�%(,�`ʘ	]�@�8l	���	�'nl�:�*W.qk�\���
%�$	�'&�1:!�4:��Q2%E�V��!i�'x��OE�\~4UI�E�F�8��'&M)���s�z��r%܈8����'�T����:l�ڴ:b��z��9��'���%AC��ږa�3s=�X��'<8����6�m[&L	�m�����'X������"���q�<�(�'��2���>K���4CE:S�NY��'�$mB�b )7(4`��Z�X�>�'�Ndh��%!D"A�fӸJ,�5z�'��\cjSϲd���Lάh�'�ɲ6,��/ʌё��Q)Z�1�''�U&� O^b]P&@�-����'�K��ݷ��M�E�X��'� �!�LW� ^���Ѣ8�z<��'h�Pà-�B] �hTJ�. 	�'J���̊	�ܴI$�^.��i
�'����mގz��:����uC
�'q�x�IQ(*�YQ����dA�0�	�'�4�g�0Z��pRR%͕Z�D`C��)��O5 8y@��0����4�B�yRgʃF�(Ţ3�C"˘�$�K��y�c�r<��uڶf�xф� �y�`ϳ�b�k5'ӬPN�Ey�Z��y���+����C�B?Z��F���yr�: <�H����"E��УSBյ�yr�+{˲���mB$C���83	�yr%W�[�|��B�<Q�8�u3�y�d\ KR�ڔ�6���C��4�yB��0s|
` ���20��D#W�W��y����Q���)!r�Q5C ��y���m~L��$� �b��q�oX��y���׌Px�<�/��"^���ȓo���
 ��#9�]�@Μ��ĥ��S�? �4 �޽w�uz�cW9=����"O<ź��S� ��`[a��\�j�8�"ORy��b��k�%�!���Z���2"O�lX�"��oOX�"_�/���zb"O�!s/Ԡ]P��jE�٫Q�F���"O&-����Xj&�Y��8;�N�p"O���u��e<X1�
�  ��� u�Ir�O�|ዃ����l��JI���	�'���A	?����f�M'F�FK
�'��)� �	�>��� %�tZ䉳�'ذq�O�3~^��Ҧ��Z��'�D�r�抯u�lJca�!L��UY�'���iA9f� �Z��I���`�''Ɖ R*��4��l���	J�(�'qV�;HW/nfL�x2�R�z�"���'�b��!�ƕD�J$ÑkV4w��ip�'�:�R�)R<}����h���)�'�&`P�	�u��E���`

m�
�'���A!����+���_�j�	�'�z������e`C[X����'��A�g���d�WA#	i@�y��$*�'nv��{0���[��8`�����ȓiZz ;`�ɭO����/�/�`a��Na��	D�T/x!@k� ܅CnQ��(�����ZS�6�R����c>���<7�e�`L,8�pJ'J]<!�����	�<I����I}`��!�,�D��Ї$T�ض&��WS�M���^?<� Q$� ړ�0|:F�ծ{^t�#�U���B�AXc�<���<�\��@Ե@�n�Vb^�<)Յ������L2{��TcR[�<�r�A�c�i��+!em[���M�<���D�]z2��+J^���@ʟ�'�������M=hU�Ȁ:�X�y����B䉏�P� �"� �j�ӆ��a�&B�>;��7���̳�@�)�!�99Lt�j�@ǫ5�2x�㠘8)�!�O��d|*�16z�Q�Í�h�!�dCas�L3p�C�$��8���$��Iq��(��D�`#\CӖ������T��%"O(Ƞ�
_�pQ��D�]�,"O���5�� �`T	A�̵,�dX "O�j�I[�"q���ǀLDJt2f"OԵa�MY�hl)W�v�����"O��,o�n��C�ދq"ځ�"OΥ
��A�k��
Ɖٱ|����'5�	� �zM���#Eez -�:NtB�I(B�詪扥;� `Pgᚻ�6C�	EezU)���o�h
�o�%"~�B�ɜz��0ڒ戛M��5�C�C��B�	�b2.{ti�4[fx�Z�G<�C�I.aD��`ض�X 0�ޟY�B�ɖ(�Ѝ⡇>zF<躕�.:�z��� �ɛI������((�(�7n2]�B�	�sn�����Z̐҂_:�B�	 ���C�%\5`S*�cG��st�Oآ=�}CB̭ha���l��0B��\v�<�-�jb�*Ԡ�Bv�T�q�<i�J�;I!�q�"�6K�L��R�<�d���X X��5t�0d���M�<��¡P�.�d�N�CN�5`W�ZG�<ĪϞQ���D��T����FyB�'`CT�O�2RC/Ɇe�~a��'����&i4ќ��H�4_ٔqC��� ЀcFLì#v��\6C�$Qk�"O\����ǿ��L���0��p���'1O}#�*�-: ��"�K�*�\��b�A>U�����d���$ �b �Ł6D�4��D'B�4]i�ӯ�6�`�!�䗺x��Q���ʢy��M0�!_K�!�%C�^�����ܜs�/��)v!�d�>`8�B�"�	�:����#jf!��T� ęY#����KZ\j���'����#$_dKh(�)B�U�VHc�'�0yST��!Ƹ��Bؠ �<�L>����H�#z탐�۩l����7���;f!��_#Kՠ����*<xvpb��yO!�ā�@�Ƚ�`�:4l�Y%K�0!�DR�����-I5
N�j �ӎ<�!�ę�!v�@S��8O�QZ���|�!��Ӏ.I��SZ�b=�L��"x!�dL�}w�(ǖ�8:�=�M�y)�P��(��i:͘�~�����Od��E�'�ў"~����-L��x��J�&�tp�B���y��\�<	����O���.=��y�)C�1��)@�("͞�yB,� �~]��&��6��-{����<و��S�Pl�����*[i���>|�!�B0�z�;=H~�Wm�!k!��5�&��%� �A]�%�r�!��7Q`v�:�C�?Z>}��d�Q�!�$ۊ5���#)��Doty$ʄC�!�<9L����W�]>��R���)�!�������Ѝޝ}1���$�i!��HHb�Z���� �ᩜ� �!�$��F+������\�rt��臒C!����HR%G~܄����ɝV!�DΓT�f-���N;�|C�'��!�$F?�Jm�ĭ��G >��%�`�!�$�"f��t��j�q��I�R!�������b���͙ H!�d�.��	�f�!����K2 !�Dо,����,�d5���5f�*!�D�0n���c�'W�?1
5�ǥ���V��(�
e:�D�!ajvQ�C+hv�[p"O(�e��S�� @\�G���"O�}фnP�e"�)�4)ܜNv���R"OL3'�74�TaW(� ik<�AE"O�h�
�ݚ�"��U'��-P�!��&���`⚏��9��P�9�!��L��YKEf<�����n�M�!��-}��r��N?f��I����<�!�DR�'S�8���T��Lrq�Έ�!�D\��T��VC�s��ACV��!�$_�f���/St�u:@,�%:��{���ڌj�i��Ғ# �u:��'a�!����\�K��N� ��X���A�qx!�װ���"�O#���r��L�!򤐨f�>+'�(�d�Iь-!�dQ�s�h
g��T~rTh2B�v!�d_:|"���'S^��a�IW!�M�V���a׏�*^4�bO"[6!�� ��p�c�5+>5��NT�J!��{�
�g��Br-�
D>!�W GX���x<�컔#�!vل�qL����[<qe��+�D�*(�P�� 8\���Z�Bd��OY!7��4�ȓ_������#I�����cTp8Ĕ��S�? $!�e��!����� 6tV��	!"O��r��<ڜ�#!��D]�"O�!��	�o�.�R� ZB͒���"O�,��Bأ!�*��q!�.�&�q�"O�թw�܌g�� A�/z,p "Oz�����0m,�	�J�%Θ�1"Obi���"A��d�:#�g"O�Ab@V�X��y�l��'
�}��"O~��E���N0Ӓ%J�*S����"O�Q��C����,��٦"OD�# ��X�3���8�B'"O���6h�{�~\2�(�!L}h�"O����� �A��lKè_�}����$"Oz��єOS���p��;N@`��G"O��+a�ٲo��)���-<�Q�"O��3#^�9{NU�e��]��	w"O�� �
Z
u���T�^#vl�c�"O������}gZh�'*-	�)�"O�:!��YER�4�Ě*�u+#"O&�jvm7�n��!g6n��E"O��aa�F�O=D�
�h�\^�4Ks"O� �r`T�~JL�EAT*x�"�"O�؄!���.T��/_�DA��`�"O*l���
?��貨��O�|�Y"O���LȐ/�x�b�ԜT�ڐ��"Oj�:�kL
oD��ǇF>��ܚ�"O������Gg�;S�@�k0"Of�#lX�](("�W���@�"O�8� f��_��ɊԠ��e��X��"O��g�/��Dh�/��Ђ�8T"O��H��/�&3ϖ�l�P�"O�y���67lL���B��р"O�cr�<&�$�##ϐ	^�%�"OhPQ��ǋ8٤��w�N�ygt z�"OQ`��O�pcf��.0��ظ�"O&�3��;����!Fۈ4�:Y��"O��{�AY3j���sEI�k�t�"Oظ�ʘ
c�p��e$ρ`|)p"O��8��^X�j���×9x��"OZ�*B�d,��2��3C��z"OF)�cA�d�8`��٫_8�12r"OH8b"�B���1'�,�i�"O���g�3#�;�eԌRtH��"OP�D�,0�N�a$�<�|�� "OX�H�� )/ŸAiD��li���2"O��`%��� ]:D�e
)[VvU�"O�M��KShA:���.xG���"O:M	� C6�94��A;��#"O!�5�ȹMU���G�����1"O&H��<Ab�4� Q�\kf"OT���kǗ4������*EF4�""O�U��'	�1�X<�扗=�f�Q"O�mв� 6a;h�O�
�x�6"O�pP�#ؿjt��i���"O�CC��&�23EF dS@"O\�#�J,d��XhDν`��A+"O�(��̈/hƵ#!��6z~��0�"Of0Ӂ�Y�0�$�����pkfeK�"O����8L�pa���&;R��"O�y�'�%@Th� �(9
}�"Ob���~�@��e��!]"�4�"O���F&ٲ0P��'IÐX����"O2z��?H�=ZG��1[�!4"O���0�֧t	nm����;tt%��"O� �zvʛu�*p�n��sJl�F"O����\�LRv,��vbfZ"O�x��i�Zmp�]!��i���y��e�T@�¤���@�-]#�y2��b>V�P�� ��"P���y�.Y��`݈�+�}��Wc��y���h&2:�J�/xc�	�֬���y�Y@�8P��,i���� @��y2j@�:���1�ʚ�I�PL��@�)�y⡗�W�<����MQ���y��_��ti��94}�I9�D��y�
	:]z���"��_��9�kK%�y���,7u���7)�)�(��)ة�yR*�?,��g�9"�X=�4#� �y¦͘�J��I 2 ��YD��y�Μ"��"�JD$��j���ybl��`�8��h�'��iP��yb�Z�L�.�DM@ `��������y��I�gI���p�)]v��9q���yr�\�q�2Y�SďQ�f��0ٗ�y�B�t �A�ˠ�0I
g���y�2-�r=b����HT�����y¦E�t���`��6U��m:���!�y2OE�5���C���D�Ht�D���y��Nb�pP��k�'q)�a3A��y�&V�P�|�(� o�(d��E��y���L�����_8�Ѐ���y��\"c;t��&�
4W���x�Ȍ��y�ɺ;P�	�](L��$�� ��y� [._p�izP�P=T�I�u�	��y�
V"�`��Q'E��U��]��y��B#wB��
�fUt��T��`��y�/�@��%�sdpm��٭�y�)Z�����]�ε��)�yh�29ޮ���HJ7-��)$#H��y�	?f\�N�)T�a��ݮ�y"J�~6U02���'𒈒����y�����j���65�<
����yrl�~����eO�[�fj#��4�y�F&.]�TYW�ST81a�C��y�^�TY�T"dM3a�0�Dl\6�y�'1DU6��&��Y�T�Q�Ƀ�y�k�F����QB�P�B��Y��yB�G�<=j�5��,]�&�S�ؠ�yB��i���!!�2T�.�yF����y��[�������O)S��5O��y�@BV������i����y��M�}�h�Q'���
,�X�́
�y��ݱ������	8T(7 ���yҏ]�ku8�@%z��-�7��B�<�EeB� �Hq����k���]{�<qwᘲŢ���aI26��a��G�y�<1�)S�<��L��˃"@x)cf��^�<�$.�ԋ���2T�#3�Ft�<9D'�{f t!��8yN"���ɝn�<���A*��!����X���&TQ�<����'������-+��1)�o]H�<��1/Q����<�Db��_D�<�P�G�W�69�D㍵Ch%JF(�h�<�QiO�d4^)R��Ӊ\�ĸ!��o�<�/�2��R7+Bi�	��k�<	�%Q�,۰��J�F9;�f�c�<�7�B*J��H5�@*{�n��b�I�<1��3v�>�33"�5�&$
PI�G�<� ��h��;S =ۆiH�&���F"O���&U)�������@�"O�ZB�G�E�e�Ln����b"O�ժ�(ޔlHy�e	�:��w"O�U ��Ů"�,ɘ#D]D�� "�"OvțqF�n*\�R�gi����"O��E���j��KON�F		"Ou[�O�H�jru*�438ƙ�"O�4q"D=B~������%"8e"O��Q��)I�5t���_���k�"Od�9���Pϒ�(Ԉ� <83"O�Z�B��<@�#��
�p�@"ȎA�k� ����&.�1��8�t"O*���&ɾ	|��D��:Z�*��"O<}���
&�VY�E�9RV���"O�E#�Ј1d���'$����"O����l�a58uGF�Q~fIs6"Oք�`O�Dm�tz�@�PzN��e"O�̉G��0���Ȍsy���D"O��å�!�J���6%]�ౡ"OR���j�),���)���/DX|cq"O����@�j�*��Q�Θ}�&��"O���%J�-��,uv��"O>!�bdA�]S�I: ���q
��e"O:��c��a�U���E6ܴ��"Oz�����V> �օѭ����W"OL�a��+>�F�ŃW�w���"O�}0�J��?����P@
=\��)�t"O���A���\(fE�`��i_��8�"O��y1%��*��3�X�PKj;�"Op!�b�]�N���3��t�Usu"O�p��b�b,	��^�"0*'"O�\�A�H%Ab�q�$+��xˀ9�v"Oj��-�k�<`Z\?q"���~�<��*ߖT?� �aJ��t�*�!�f�<����!|8)Y�Ջ1Z�˷��K�<� �,p������M�Z&��B�K�O�<�0
�M�b�y�[����J��ZL�<i��:G4�MSDI,'�b���]H�<��G!.L2�
��_46�cE�<i��";����!D�r�7P��y�*�O�����U�z�֣��yR� 3U	>���D�$��!��J���y9)��]�& �H���$�Z5�y���2��#4�'h�0��"���y�,� zBZ��m�>u�0 Z����y��ҥn��Q��@\%����*�+�y��'j|�`h�ck�Jw'���y�a�� d���.a���M�<�y�莓L^09ѵ�K�[H��y�/;�y�!n���T��]��x�� ;�y"���r8Ĉ���X�]J�Q�VGN��y��YF���z�Pi�=���Y��y�GO-%vH�y ��O��{�$��y�h
b��)�S�OG����M�&�y�+U�@yBH���W.C��l:���6�y�k�QH�o�:�`|��D��y�!]:�I�iڵ6^���u�ݫ�yR�G�
���H��L�H��4��y�-]�d9����K�2U��׆��'Pў�2|�����.Y�'Y6"�e��"OTi�O��I;P GئI���i$4�DhVG��4J́{$+ʈ:� �:D6LO.#<�FX������Hw6D�� 􁉗��r���B��,D�P�AQ��9�S�ӹ`
b<2��I�7���sS�-�C�ɯm���[FA�
=}@łqJ��͖C�I�@���D`V���2��B\��B؟P��P�^�Ԥ��*�r4�l&L)�O&OZ- D�˗v�ڔ3gH�jMn���"O�\����(E���åc��>B�30"O�	)w��5a���P��ͫ�d�9P"OHh�R�_3`����'a�0�p� �'ў"~�3��[�����
\��z�@K$���,�S�Ć-��$ ;W�HE@���|�j�	A!�Y�:�yբ]
�H1Aj�'S?�'|�I��HO�)^�eN�z���>OzU���&P"!��?~T����<Jih�i�`Q%��T��$�"~���ہ�v�2�.ҵ3��%`�L���y"�M�<Z0���i�8$��0��y� �7�8�j���`��"�����'\ў���X�%(^ĸ�BP�� �"O��H��՟)�*��vf]�"F~��0P�l�<��ԟ��8��#W��z %ę6=�M���'�˼�;�B�>�-�Dюc����Ix��������v���ڣj��eL\�#D� ����3X|4�Ge�#�<����/D�d�Հ�jD����r��%�>!J~����z0D�1I2o��d�F��w�\C�	.S���J�H���(�G�"c&C�I9@v ,&([��nA�E���,�C�p��TE��$!<	�@��RhNC�I$
�|q�?9Xx�X�a]1|s�B�I�,��(PB�ɺR#,��
%>ɸB䉈]|8�*�
x�M#������6�S�O>T���O��ݺP�F/�"�S�"O��8&@��E4m���C�A�,E�!S����ɪ`�4��b4>ѺM�������D<�$@6z�N���K�4�>pZ�(��-(!�$�.$xD��34cf*R�J]�џ�E��Q�
 a�#c\�"9�AƁ�0�yb�1a"������������yB ��g$N��g�`��iq�Ɋ�y��=d0������Z2��q�[>�~R�)�'$t�����H�LCK��Y���Ey��|BV
���G��8�֝���^y��RX�D�cHӧ	*M�D��L����O���'���	�����,yz��� \�j�:�;�o�	}�&�)��5��/ޟ8'����	&q�a��������yR�?U+Hʻc=(�Xb(�6b�@\�W�8D��ŧ��M+&��]@��@w�&�o�`�S�Z��#hxdX94k 8>!K��,�rC�I�g3�i��.�?\��& "Vu~�[����Dx`O:�����@�],�MC ����0?Q-O���M��hg���f�ƻL��r�|��'���c�O�f���9�ѫs����B(F���S�.A����J�g�� �!�~?XC�	&��u;����(����t��b;�QI��D2�g?�G��2" l0 �j�EiBL�a�<)4��1,d(��r��I���������#i:����)|�-�7��D��ēxj��CO��u��r��w-��"O���WB��<H�4r)��0�I��O�����L�8�/�`1����Yۡ�d�=/�sC�$�.1xcgQ���*�S�Oi�:�b�+(�U��5����	�'�n�0` ��.���k��?4�	*O����ÉX���˗*Y�P`��"˺{?�}Ҝ�� �9{�AB"c�|C�oD�_�xb�"O,S�K^'� E�c�Yop|=��"O���da�.z��3��A.BL�"Ot����D�!�Ȱ#!�T7����U�$*\O �*���1�
�$���@�"Oj�	%��$���Pg�	-MH�"O�d#�AY�T��H��[
4�ҜI��'�O�Li�C1�^�X+����{6"O����R�2g�f�BI{����"O���A�w� L[ԈK
��"O��	�ki�"@Rp��*�|0�"O��.�(�H����+@׀xb'"O8�s��/ZA�=õ���O����G"O���d��q���ó��
P�0dca�'��I�
���	&�[|��!����UЊC�	�g�� v D�@7$�"`k�4C�I�n]���ǝ�/,�#ဇ`��B�I�8*� �V�^�<�#on�|B�I��tLy��85mT����&skB�	�"�.u0�J�
C���Yk��O��=�~��i� ��93`T�1�L�2��[`��<�'Q���d�D�0(L��#K1O�}��}��'�V0H�
Kk?u�$�}�B�/ ����E,T����X�Oϡ6<�C�	$i�fpʗc[�`fɴ���g��C��=1��PZpH�$t���`E	�1��C�ɡ3RzH��9��	�C�87W�C�	�?�X�Ba���gN��uɅ�}xC��c�@E��JɆ����$-хQ@c����	0G|􅠲��@zm r���C�C�	���g-N�Th��_�Z ���9D��Z���2i}�x��B��-ʈ�u,6D��AA�ڏM�``V�Z�l�n<��/D�4�5%L�'�ґ(�KS$�PE�,D�8*v胢c8R��E�
�pv <� �-�n�
��<����a��@�1�����IS�IG���P���Z���.�+x��V�7?����hO��O\����/X��i#��J:b�F��O��D[�!Y�U���+~3�IcS,S���=��<E��Y�m�"Y+��Z��$���n���yB�]�(ò`���P�V� ʔ뜡,�Ni����O2l�b/�)� �6�J��i�"OX��AGƗ\R���63���`b"Ob�rv#�U��`Q2o%=�T�H0"O@}��$�Sn(��h�(]���i'"Ox�aG	�s�x�t苻{���aѓ>Ɏ��	P�P��[��27H~����R5��`F{��ԴK�HB�i� ����3�L4 ���5lO t�wS�"N`0�\�@���i�"O� �PY�`4� YG+��p2�h�"OF���	N�a���钵(2x3�"O4hcv(
*�|��v���]���"O`)���!F�e颡�;W`���"OViQ�R;6GL����Q$=��"O�]��i
�%�^����ܪU��]�B"O��� MM�	b��(bN<�,e�7"Ol=q�l��JzNx��0x�F��@"O&��,ӧa<|XUn�0��ͺ�"O�p�	Y#pNUkA��1j�bG"O�`�d̡|��u���C� ]�5X�"O4��⅝4c3�tQ� \�3�"�b "O"��Ɔ�2�b!#�A�]��BF"O���3A� \����3
�p��"O�X�b�=qGl�h��ٯ<I�s�"O� ���w'Q6� G�n_,��Q"O�����>nX�ˢLJ�$O��:c"O�*�
;���K�
D99��"O���T�WQH�Q���o;l9[@"O&��CՈ+]����'	V�h$"O��wkI�\q�ȡd�<c <E"OΕ[�� �G'��Ҧ�T)K\!��"O�}���K;bF�ʇh.?�-+�"O�Q���	:G
�����N��"� "O<@��^hr�X���φ!ʚ�9&"O XI +�� ��E�>��|C�"O,�rt	�A����E[�"�hx1"O�`mr
�)��N<S��j�"O�is�!/]������9>di[�"O0C�J��8u�Y�#�L�ʴz�"OzŠ��
S����T��(���b�"O�%��ˀ+b*m��,�Kh@�� "O��@�_����Ql�Q}��IT"O��2`���
a͡'a*�b�"O�� GB8���qK�<IX���"O�	�ƿ3�@a2Ɗ֔}8�Ԣ�"Onl�'�R"! ������1SJɣT"OK;)t�|��O�(���.�y�MN�<$V��jF�YI؈P��Y��y�BU!�jp3��|�|� ��<�yBg�?F�);�G��m!�̰���y"���rM~yx��e�j��"�&�y" �;o�px� >�P���W��y
6*�\�j�ӭ���b��y�*�w���2A�U	�ve���5��'�hY�g��|��X�;@	�yBQ2]��ͺ��Q���%"2*�yeQ0bYF�BèC5P���ч˳�yb�Y)gF���횢W*�1�FM��y�@�#��p�d��J�2�{a��y���|�N4�sH�$~�r�S��yrc�=;�vl�­\�l��07N�yRf�$�Z��tH��+�ꝃqK��y��+�aH�U�����ҽ�y�+ڢ`�´��hPAep	q)"�y�'S�O"��Bf�3(xn�zjX��yn��E;�MQ3/L�p��ybc^��(�] H�2d@MI��yb/N��qp��-{A�e�0	��y�IA�s@I�È�C~xY��,_�y�iK[/@����Q3<������yB�ú h�@ ��"Y������y��m����cO�jX�r����y�gB7pl�����X�&�y��E���y�AL y��y{Æ�#~��=�5d+�y"(�>W!X�˒gE�l��$�f��yBh�lT�-c��a���84�+�yb�0^��H���-��ZՁ^0�y���20P���)	4�GL���y�E��T�D�ƠA!S��7ᖋ�yb�2�t Z�߂@���DX��y2oM�k�t�A�c����1����y+�:�����F�䬩x�M.�y"�G~�P�Y�*�*U~����X!�yR�S �8��e$`�a�	�y"-ݫm8*8���^�db����y�@Q�.~Б���VA�H�a����y�	P�8���v+M�Dܾہ�� �y�O�,7P�x`G�-a�^8z�/T$�y��$��FEb����/�y
� �ps��A0on���I	7����"O��"�(��A"81��A�K�i�!"OZY� M��_�Ĺ���մ2-F�t"O�T�7ñjx��Y�h2Vd`@"O�9�֦Q�_"�#�쐏i�y�u"O`�XqڍNbF܃f�Z�&eBA�"O� Bu��p��Mw��=13%�"OHx ���E��|���:2 h�"OR�ŧ��t�U0N5.��"Oe�B
�V%đ�6�4&7�8�"O��"�W����E�K�|,�:�"O< ��n^*(��q�u�m�p��"Or@�P�	C�X�)Z�Ҵ�hE"OZŐ5�Q}8�b'莵W��t
"OB���ٶ(<l
'��!�n�;�"O���g�� �!�vȉ�sLP�"O�|� ��C�����m�K��3"O$�+�S�d� B&��4�U8"OZ �Њ�$%Ux��1��?b���r"OD��0N	�(�k`D��P��(�"OXm:P̒�1Y4��g�O4���""O��c���s6�ib"�L��:I�"O�Y$��,P�聴��9a� �"O�Ur���h~t��N7J�p% �"O2� ��]7tX
G�1c��0�w"O����˔�`���v�
ň�"O ����LΆh�ID����٣"OĀ�m�!{���G�� m;��"O�y��L�`|��!g�����"O80����  ��f	dx�d{R"O2��5/Y�5�H�QEXa���"O��p����D�
`��U"O�U!�M۰: ��1�$�88/��<�`[�SI��Of�h#�K9!$��5MC��=bd"O��c��4_PVx�!L Ԫ7�����GD�B�
�E�>E�tF�'��r
�!�h ����yR����ڷ(J�\�}X� F2�
Y���O`��;5��$>c��ఫ����R�RQ���Q2k%�O��B��/3�}�%�;k�����[k}�9bd��6iU����A��\����#�qO�
6h�0�c�O� �y��3���E}r�	Q>z$��ꀝ(�!�aX?9��L�ph8��cf�<;�5�Ǣ��.��D��|��-�g}�D�/�P�����>kD$��!���y�JŮz(<E�3FE Y.�Y�Z/�R"}°��8�^-��:<B�΂!j̜SA8��\��	$v98�X�B6n��gÇ!#�`Z�#�7� |�Ylt��q��y���n���G�!	-���	~�h-��Ê�/���wc�B���D�)C����ȗ-3����d�B�{wҬ��b>>9��j�I�
H�&|���(*ȃS��-5���7-b��ȟ:����A�H~ T�f$��Y�i���Oa`1(�iSY�5� #׃z��ԩ4&<��X��M��;�� 7�@�|'�a��鉦�N�'���'��>Y�b_u��r`k��H1��CWڟ��)��٨�.�3l�	q�Zr���2���&^����rOY�g$���醴3="D�uh�-*�����[U��W�ߜ7��! AK"�@��e~y��1��\$��P"�Z�'�"u�\��C1Uj�D
J�=���|��y�"ܕ}G�}B�@��� ޽���w�s��S�!Q!{2��G�I�wk<lYGa��"!�WC?x��+�lXDX?�`��P0V�f�
C����Y��ўh� M�d���@�G�0>
 2dF$
��� ��Ehs�T�H4��k�@�^"��`O=?��&��>�d�|�O,1�P��9?L¼I&��7�hZ�'\�ۣ��`H�P���"VW -� @E�<KΨY6�P����e6�<eI�o#G/�����Rs4��Ɍ(�CNW;Z�	SN^�w����� ��3�x�����%���+7J.rW��!m�yb,-��(8�/ѻ<2x������0?���W�a>H��
�	z4w��tUtP�˛H����� G�p�*%���6*����=�b��^���	?h\U�&���,�4hkbk�Q��>�V@U��#�i�!�u�(H��qK 
U�A�vݠa/��^�,[��٥cD�2�O� ��"F$|��Y����R)jF�O �C���#M�$p�ʑ�3yl{���s��8��[�5P�u�B�=m�l�@
�y
� �d{�O҇:XD���)P�����O��V�&u�S�Ķ�n�:%��O6�(5
<?14ܤ*�nL�c瑢@u��1�q<9M$R�����)�ЅA�̸(���:���=o�n7͘:2n��!w���0<) �B�x.���b/��
�Z�[��h��ca�ܕy��P�k���@��#�l�2�ӣbM���� l�&�3
�'J��i^6z���KbGI�a��,O����I�&ˌ9s�'�<��fv�c��|�U��+�N��h����ȓ���2b��[�� m_
v(��љ>�c�ڼ�D�J~�=��M�b��A�!KC�DH���L��ĸ��}������G� ��Eo�9k�8tz'��a�cɸ8 ��V%�N�"�0W�T��O~���N��
�4=�L|�Q+��G�E�(�9qG�A@�<�PM�` �"'��Y�,����FYyR(��i�~��`B�j���{P9���
�m���7�ĒՄB�	��!ۧ`�����b�*MnH�0I�0�Q�D.P�̈&?㞔+��1}��:4M^U�Bɒ�$3�O0��k?c��1;�D�dʥ��@��6:>��i�3L��Ja�<�O�|
ѥVH�.]X�N�)(�:��'��P�%Iuc]iaH�E`U4}z\�q����$��yB��hpJl@�M�mȲ��Q)���ٔm�]�Qkƽ�EMI�Oڨ���iS�W�<�s!�P�R����
�'��A�#ƇY�|���טWN�e�WIA2v\��7}B�h�V��
5�L�!�o�/�\E�ŀ*D��Qi�o���)fv; %9u��Od����tk(�p�R�荺v&�0�� 
w��9Ō�� r������ِP��v/��QWM�/8�>Y(&�Q��yC�LM6��B�&1&�h0ŭ@3��'��	8惇��dD�$�O�{�D9���3�L���B��y2�ki����,!$����_�� �6F�/?��'-�>�I+: �PdaI=+�:)k�'<.B䉚:��)��@��0mh���:��(j��S�=��X!o��򭔝Xv�բ ~���sV�3����	E�p�����Iz��#e�ո �C�D�y�)*�h����+PV@�<	EEE�#~���?C6Li։N�4���D�f�<��{��I��)���#�J�<yR"B5Y���ƿxq��;vB%D�k��^�ê�솗p�����%D�d9$��@�0�C��S�J�X ��5D���B�2_��Q��>�豪0D���)�`�1&���QG���j,A�'����3��2	�Fp�F�>`�J(i�'�(�Á�E�X���i]%_�t�I�'Hf��bbI�"r6�����!C-���'Y�E���	F��)��=��X��'����`*�ES~�qK��`�2�'_,m�D� w*�&oۃ#�T��'�R�V��?F�0(��%��|c�'���TC��(H�@Ť�7ڀ���'�H��A�B�^XV��;�`��'���#�I�q[���X���C�'��(�Ȗh-y��� Q�8��'�b�p�
C�F*�G@,[����'�\%
A%�\�ђ� �2y�
�'�0y�W��I�N,�� Q}�b,�	�'l>�[a�N����v`��'��}��L,cT��*t-a�j���'C� (�(V�<Eb��[�TZ�"�' ���$��y��R��O�;_�<��'��U�ؓmަ� �H��$��
�'�̬�D��><Q(���&���	�'b9�l���e����+J�R	�'Nt`�GL��t�B�Pd\�����'�F�(U�7��)`��aJ	��� �嫲�@��^�[٤����"O�8`�ϗ�;��|C��LZ0Q �"O���:H��<zAϟzD�"O�A�V��
_X� GM9�����"O&�����#p��pc�Б�X�"O`����g\�a����6w����"O�����'s�$��bY�H��a"OJSd%�N|x�.��0�U"O �Ն��1��h�c�C=Gp:Ŋ&"O��0UΏ�z��K�)torq"OdT���3(��	�w�
�:E
�8%"Od�zD�����"#<4d�z"OF�k�A���@��2i#���"O�h!��;0Q��T�ƒ*L!�$"O���bO^'��T��7��8""O6�z�J�@)�%�1 �3#��٢"O6%��`^ oVDu���4Y����"O��`������*�$�.vf��ZV"O��p#�-}!���C@9RZ��"O [!�N#c�1��m��n��"O�"6� `��H2 �4+V��W"O ��#"E;B`���!A(*x�&"OL�s��;J�,�C�@T-�d�S"OxZ\��$P����,�H�'�.�y¯�,����*ۤT���W+ �y�&�>wZ�M�¯4Q�%S��@��y��!�����
�/оhu�W�yBi�5+� �AS�LMx8q��Ȧ�y�_QR]B��99UPi���yB��	5�6=���œ>s*D�(�y�i�='�0{��?O!��R#/��y#��PzX���HBȤ�/��yBm�2V>f�q�v�COR��y @�lO��x7f�u�@�C�A��y���Iu0p���A �f-�!��y��=-�>��GgːX�өǝ�yr�9^3�h�@X(Z38�Z``E��yb�D�.�P�ɠ+9\������yBEW1vi����f�d26���y��B�rt����n���\�H��y���a�Da@��� #F����?�yR)B�s3���4T|d@����ym[| ���)	�R�$"��G��yB��K���a��*1���� U��y"E�84��Qlְ3�`���!��y��L�2�S�
G�}eb�@ec���yr/��p�h����m�[f�/�y���@����� �u��L�(�yC�g���:R���J�,��c��y2�w�4��$�h#�� �ybAh;$��!b�"k��CǊȐ�yb'��1CHT)C�M�k��Q���� �y�����p�jL8~�6`Y�� �y���*1[W��3j���2��P��yb$�+fHP��*
�Y���2Q���y2b����zr��ds������y���"�l�@�Ê�fJ�� C!O%�y�߃~�����!��S�C�,�y�D�#R: ��3k��$ N�+�I���y"��]�~�jqh���#d�yr�^?E1�D�6�q�A��y���6i`丢��L�(FJ���y�'SN<Uҁ��Gn��1�e�$�y��T�Fq:=j`��49���h�2�y
� "��S�9Z[�����:b��T{"O�&��t�����$/z��E"OŘv�Q9v��}ې.ӸJŘJ�"O�Q�`'�v���-B�ڑa"OH�p0H��5�|P9"l&j��q��"O ,1�DQ�c�ڐXcA�*Yh�Q&"OF���� - a�Ё��<W&��"O�;b�G��dY*�`�!MA�@"O�m�e�K\-V��e�5)P)+4"O �G#֜�V����"撙�7"O���U+ �Е�"��.6���o"OL��D�4!%�D=M�-;�"O�pS�)�	�Аu��=�
�Z�"Od����I�$5ϔ���U�`"O�x�+�>y\��Ba�̓B���A"OzT�a.ū��]�f�Ebvd1�"O(�4�[#L�(��
$t�P�D"O�t��	��Y^p*��>r�Q��"O��Su��;FU0�I�$ı_��=R"O���/7p(!�0����!($"O��*4QuL1a�cãE�0Y��"O���	B3I�@��0��:�Z�I�"O�p����V�%�g _�N���C"Od�	ǦR'���2��:1�hM!t"O��lNA^�<2���4}�,82�"O���&ʫD�A����P�"Od%"EF��I�F�Z��ӂS��X�"OPP���1�,��Y�-��aIt"Oh�x�
K�Y5�M����<P	��"O�=���3R�T�� AD�d��"O#U,ņrD؆�P�4�X�w"O�!iPJ�X"@yY��Z�]���"�"O������%�ϝWG�EygƑ�y�12UĮ�0�XE�V���yR�¨(RE�Qh��+R�mx�M���y�
+0��h¡�$����% N�y�
Y `B���U��a��J>�y�A��d���F����/�)�y �=)�@��a�6<nH�B�ʌ�y�JJ�J,��a�brܜYSN ��y���j�9��Q$c8����H�y2胨�n=14ɚQ�$I��V��yr�_�|�$)�Q��J0�-������'��#����O�~��#�ߎ+H���d�^����
�''<D��&�+˂=Qd�XȰ
2b%zoּ&����Y����ף0*���A[�Z�Jm(p$�	�ʈ��ɯF`�>	1��A�+Ӷ1�N,fw6�[�ΐ�S�|�B�K�q���dգ'r*� ��$h�޸)qֆx^)Rr'��`؈A�.Ox��O� Q�u�̋>�:���'ĸ#�ʪ�J�P��،*��:�'�LA��E@6dx\�t�$8\j��4xY
x{�'��Js�!p"¦P�@]�/O(�Q� )Dl7K nT��-N#&����2%XH��h���ȣn"�dY�b��7޸�ǀR�*���SA�Ix��r7�
�w <i��X�`F�\F�g��kդ`��ˆHq ��׊�	l?qO��S�l�e�hˆ��$��O�~����0�t�1AV?��m��C�9b13@��va|��Xag�YA���(�L�a&Q�攩q�\Ry��'���O�:$�C�9�4�2O�Q�����p�)c,��y�"O��a�D�F`�F�W�08��`IȰC" +�,�k*`�rccN���+�Q�������?=��I���IR��t�۠�Ӷ�0���E:^�"@�4�E#I�*Q�v�?b�|��B�\2R�@ M G9|�v��N~"���D�f���L�Pp���%?ZP���U/@V栂��"�I *v\��AB2"���B���O��� 7m
ڸC�K�X{����}>l����{X��@��v��`Ũ� ?��j6�^�V��HGnS���:��m�D��O\!���h�~˓X��a9 � 9|��2��<}T�`�ȓ
�B�/������:e�:��	(�(��b�ݮ4���M�K������e�� $A���J�\��'�2���ʂ�'�������%�P� V�[�|ع�K��J��,�U<�@��n�ԁLXTyh���z�'ְ���@-�l�|����,?rB0h��T n<�=�"d�Y�<a�OV�BaAÅ)HHE됣V?P�+N�hqj:}��� ���	����[G��0L�!�����R����E�*<���!�� &����۸�~rE
� ���\�� ɒ	�MI��Q��A��JC�� �Gs4���+��4	�7-���g��~��3�V4��q�
�'n=ҐI.#b��;6�D�-��h /O��y�������'6��E�r�'a!`\hE@
+ounP^IN;�"O�i
Sn\		�2���`	+�2)�F�f���U,�M0M,�����4�Y��\�4PpcCL�I_��e̚��@"��{��c��2�PE��$�0���Ɉ`���E�Bb,��td^��?�⃗/v��@h3�i�0hɀ�����I-ΕJhJ
^5!򄄖TT6	qnN0Ex���Qn��I9;� u��`��E�S�O�B�f_T��s'R.Q�F1�'�饤U�&�:L �dK0H�4��TO8}"fI�d��Aha���{�.8 ���jTC�� (�4�co�:��?�Ď��Rt��s�Rl.���A��#>�4aW��<�.�Ƣ�=�0>	��K�#h�p��N�g�xA��q�Qd�vs�8��gKZ舁�ɋT՘�aa�U4s�\��Gȃ�C�ɡ�F�B�G6�T��I��8�'=0 ��o�[~m�b��Sɑ>��g��-��d+Q�L����/+D���AI���Py�Pm
�a�!KB��p`��ʕ&��	D��~r���I�"D�c`��J��S.���y��P	W!�q�Dᇍ�6f����?aEb��Nf��)#lO����$FH�qfL�p-��A��'c̘Z��Qo��lZ'^n������4�Д�0N�T(B�	Y��pH0Ɣz����)ά���̱�C�<���ɰ�+^�F$R�$K��s���4B�x�ޘh��3R�ց�+ֆOa����3�(3M��G��'^̔�A+�5("}�&T�mڈ 1�'W�a�`�/l�Pxd���iҝ������F�E������
��D0�#_/^|�$��U<ja|�eх��A���'�����V����QC�9�V���'�>(b��P|(1��J���e���۶y�: j��I��s���u,��[�^��%SV!��[2<�����>��b�H̼eK!�D�-��.���h� �r���"O�h�䀋?T*�)�!ˠk�%*F"OX� �z}��څ?Uz�6�O�ybJ��&�-����9J>�V䒏�y"��9J�8�\�<@&u�t��yR��b���t�*�<x����yR��>sOe�C�*%sP��,�:�yRlC-5`�i���[\}r�U�y�bܺ�s����Y򠚭�yb�E�z$�Ȣ��{�.i�O��yb��~��� Yh�ĀAƉ���y�����q��+a��-�^���z�
�H�Z9,L�Aj�O6b�TQ����E��\�U��΂� �f��ȓ��e���>��0"�4AW�L��"����F�)ry�'@ԲaoȰ�ȓ��= s ���jX�"�-,1��ȓn���#LM�4�L$�W�/r��х�yU�|��� ���H&5F���7�U�s�ܭ)�҄��L�DE�ȓ$!�}aU6g@���S�u�(�ȓK�H�B�,'�9rU�#.�y���-C�m�����#����#1���j�l�af֑ma2y�׈;w��`��S�? @�Z�얞�����FתLŚ$z�"O�Tb�X�hP�<�vJ�X���"O�Q����dc|�X����f���"O�����:NP ���-K��%��"Ox�`��7 꼢w��vѨp�w�<���=`�|iEa����@b�T�<�v�׳�.�k6oQ#X�X���<ɱ��9�]r�3!���%&�{�<�%M:�Z$��K5q��b\�<�Dϖ����	�ǒlƐ��V��_�<��
+۠��	
�=+�@�U�<Y��	e���b5���X����CR�<֬�r�$����%�t ���q�<i!�����(��LR�fL�R� Xo�<�w�ʯIZp(+w�/j�V��R�<����?��DY�/V+?�I��G�<�bM�{w�IpiU�sT: ��&H�<Q�᝖A���$$*T���a�D�D�<��hP�~l�J��h�B��R��|�<)cN�4 vmQ�	5gUz�SE��}�<���K(y������8h�Z�QU	�w�<yV��0e��K���#! �����n�<�r&ԃTșZ���S�$au��c�<A����@��E�D�)Ȉ%+�BM\�<I���;&���g��,"�(��2��t�<��D_)8���m�$ ��A0`,�d�<y��Adȵd�G46 ��E�`�<��C}�L���!�
M.�i�+c�<q,M�YN��p�o�.���A�Bt�<��k����!��jJ(iD�(8��_�<�3jն4���㓩���xb$WT�<q&�����0J��Wy��5��R�<�g��rD��$ !����B�@�<A�g�PY��jtM��Z����<���3�hai��č; U8��{�<!�I��*���al2��5��)Zr�<�TJ�>h#��(��%+ d�ㅦ�e�<ɂ�� ���ҫQ�V�	i�J�b�Q�54�@!+�P�H��K�,�)�<�-��S8 {7������r�\�<$F60��
��T7��uf�U�<�r;E�D\�l�	;��]�<�N�8+&-��@�u���RE��W�<�G��9J��"	��X�z�W�<��ꚯg�p�K�=H:�Ѐ��PU�<��oZ<tD�=���(�S�<����;\a�H�ǐ�?P�, $"L�'&��Dx�O~�q��@ 49��td��ZB�N����"-��$�����S�'d�>%�%���fRp�!@�`^��I�XV�{ �6\
4�����0�P�v���A�]Hj���	2m� 5(���I|��h�t��.�����	��7t"�JMy|���_�	�8i�'E<��	ç!�F��QB�!�@��0&�
�8���9��dJ6 ���i"�i�:} �(UO[T'^���B�TkN��'X�XB�C�Z���S���䫤���uD�YhT��'�\y+�@��!F �b�O�>ź�d@�TO� �7l6D�.��&�[�)OTi�$
3x�~ҧ����x�P�q,�@!�"��4f\��p�'��Z�$��
�$?�3���%o+�]�@C�;~��u�\:!��L��"�t~k�x�O��S�r�v�� $(B�Ѐ�!�*��e
��j}�=��D)��OD:�js���;8U��ʆl�jl�.O�T���+>���:�g?�flB�z�̪��?)���0��<�g�˭8��鳒�x��ɓ��^����q��ě���^�<9��'T�J�/[���dZ��XJ�
��'P���� ֱvN�����-:a�d�	�'�z�`OW� ��a�Q=-1��'���  ���   �	         �&  �/  �:  �E  �P  �[  �f  �q   }  ��  Z�  ��  V�  ��  �  t�  y�  8�  {�  ��  �  K�  ��  ��  �  b�  � M �  u �$ v+ �1 F8 �> �D K PQ �W B^ �d Ck �s �| A� Ċ �� � B� �� ɭ �  x�y�C˸��%�RhO5d��pJ�'l����By��@0��S�F��L��|�t���<d��46����U��(&��M´$�
f	"��ǇO�W��I0�d�>M����Kՙ�uG��^����+��4��m^�:�Ń6U�E�6nج�X�B4h�T0�#?�0�*�	\�E��]�9j� ���M�4ȝ?'��05���uCT�[6h��K�q*bl�-1�R�
 |�u@�N�]9�6͎>����O\�d�Ob��Q8y��x���o&U���%W�z�$�O���O�����O���f�tj!ݽo�PY+�o�>�L����O$�7���O��H
}���<�d��Sx�����n��@X�<�!/E!�IQ�dH,<J܄��K�ӟx��EN�J�x99T+��3@�<�O���	2�\�
��V�o�PaĂ�>j�@Ä3s�Y�,�O��d�Ol�D�O���O���4�,z������y�Le�X6�:��X���m���?Q�O��o�H�4H��	�y�9sF,		
O��%I%�(�G{�N$�']LH�`�-J9A��{���&?D�ԅ��{�'���&aǠH�j0BF(Y�.�)���hO?-3��E�B9KUeSf����v�ZPyr�'����>4���q��̏a�$���$�<���K��B�^�����Q������ �?���S�!���a���v�,�2�@-�� D{��dI�7���Z+{��5���S���ydlUd�|r�'��*���ȴo�?C.paZ���PGΘ��a�4��?��82�i[(�v��]o�9�6��#͢����0�tM�ȓq
X�!���U%��L�R���	4�?��L�x��T*�텽/ J}0��H�'ߜ����Z�p��+�, k���Q��z(��OB���Q�E
��P��uչ�OP!���u�hd�". 2��ix����!��X�^*��f�؛0s����^�
�!�d�3g`B��vh@�$���B4���џ|��I����$x�O̪l�Z� 3,��5�B�=�O�i�O`�d:?��gN��D���BU�Q&Y��-�m�<٦ �+&,��BM+"�.�i5Kf�<Q�
/2�%ST闦Q�<��R{�<1g��T��[ ��~�l5bKt�<���(?Â`b����4q7ktyrf&�S�On�+�择�D26�ł	 .�I)O������O��$'���&�Q��D�w^�e��`�/B!�S3}@�gC��s ޏh,!�DA��(1�b�5��-��.A�!򄗜X� �1E䝋"q�u��J�!�ׯ$]���D�K�I��9q�S�,F�'Rpb��3�w�(�'Er��V��-�� � U/_��������?��O���A��ɔUo�e�OD�d�n<�8( c�V�6�Z��'�8�r����"�|%�OX�Cf�K�"Ȩȅ$K�~�8\(��'^p\��?���?���[
m8"�E*���* ����O�⟢|�'��7��+`�d�V	ؔ�D@�����(�x�bO�p���BAwל���Pybg��6_�9O�瓶id��ꠃ��t����B�
�%Y����O(Q�����qO>u�7 ә� �Ҍ�[9���<?!���-;Ӗ�"|
B�,�Nxccσ�?C�� k�v~҆���?A�����O]�����nz%�`[����qN>����0=�!�M2
�i��U>���hA\T�'6£}"E�!J��C�����n��v�ϟ�YӇ|������?��OL�����	h!���b�
��S4"O �U��R<ՠ�$�K����"O�ѡ��Ky�9ۀ�\8��c�"O��&�U�\������e��Ii�"O�E�7� ?-����+7h��Ac�V�,����S��:x3傌.��8H��X�V�Z�c�mi�8��ßT��y�)����^�Ή8ŉ�|�@=H�� SԆ��'�])����2�@q傶Ҽ���	�x⌚�?K��8���.��$h�ۜr��)���?I��?/O�3����1��
�>��-G1<��ȓ�ڜȄ�P�l]PL��èR�'���4�?	.OX�*05OP��4���K[�����O�P-���IN�IڟP̧Y�l%Ex
� @d��;)�(���\���'�����
�Mr����F��ZM�$Î�ax�Kž�?�y"�X��SD�1�hܡpk��y�IF3=[��Ʌ�;~ d���Ƣ��?��'w�H���S�1q��R�i[�� �L>����F�'�R��4�'���cA�0ZMI�f�
MJPs!�'v�%��_$FpHf��,$��)��ӫf}���%�O�;,2z�1wOfU�tq��>o��3�t�H�j�4!P�CB��	�3*�Ļ#���`���A�P �eM;k=��'�N�(��GԛF�'-���$�'0����@S����B�0g�:ъ��'���'���'�j@�ؙa���*�b���"}���D�~�OD �%OĀ�Jt�֍B�6n݉�iFt��4���O�_�,x�O�,N�`��!Ř?`#���Ht:2͙+EZ�9@�3�r0��D�]#���;uh��@*��X��z���TaX)ed�]]�w7��ȓ&A�%�"!
�'�$�j&��
z(V(�'S`#=E��O�qR&�����*;���� �����<T����O4�Oq�b)��ׅGܡED_�8��P��"OH�SB"W*����m�|����"O��ӡ�@�T��[�U��l�"O ��G㈈A4�C�߆�@,�"O��PQ!�0����'Q���җ|��#� ���P�~��Q� _\��1ain���O��d��O4M���E8_�c'�*,���;�"Ot�Äc�:78!$�L�G� �"OZ��d�X�	��L��3^�`ͩ�"O��F*�@������!�LX2��' ���dDy�����9i����P12ў4;щ<�2�a��Kȥ|��,4�~��r���?I�x�&�9�+<��|`�)Q��ȓk;~3O��&Yx%g	7�j��ȓf,\Y���V��f�W/"��ȓiHP�d)�>C���s� W5\'\�D��-ڧi�|��8(5�DK��&/>��	�0�4"<�'�?�����D_51����N�4f�.YAg)��y�!��]eJ���2��e�%�Q�%!��H�p�4q)ӭE�a3�d���;u!�2��i���	6@#a�P)%^��d�!AQ�$�NQ���pQ6��6��DE��(������K�J`�$h�o�v���3]�|�dO���(��p�)�-Bru;�h_6M�J2+���C�I�{�XřA�H��I��MB�UvC�<62v���'ƠWn�u��f�i�6C�21���߆@�RY��5	C�I!EMV�k'�� ]0�I1Uꘞ�ȒOd�F~�����~2�^�)�pUq�oU�c�j�����?J>������p�  �Pb�5����4��(��B�:9D��`��>[�DUB�O�6^@\B�I�-�V	Җ��;:ֵ����.B�	�P��T�N<.��%�3��Pg4����ן��5�؉K���.Y�0k�!��G!ړz�0G�T�ZG�>�R5�Y��[2"B�'�a~��79� f�6qБ�����ybL
2��p�P�\�Xx����y�8\�9���RPE��q5*ϩ�y�IłZ�|���]�~��su���O��D��bye�'m�pR����ך�?�a��Y���4�'�2��`�Z�|a����G�=�
=���4D�\qB�ƣh��m�C�
�r�$��!�0D��:�n��V>��`ᡞ�r�L� �+D�h�	Y�Y��DҲaް:�~��)D�,�UCV��<X�afܿT�8)���<	��)�'���I&"�I��A"_7
f)�'��ٚQ�'Y��|���JU�gE���-e!��!T�y
� ��*����w�^L���fG���t"O�Q��N0����Wg�S"O<���n{���k��[^GD� w"O�r""S�C�h�!�Dd�� �|�,�]ͺ��(!�JF��G�u{'"(1�H�	k�I՟���O��:Agl�����5i�� '"Ob�#�N�Р��!�	:Td0��"O�x!a)�^�PAс�=�a�F"O��ë� R����/�IF�'K���	���d)4��/q�Qh$ڝr�ў����;�M�v$۷�
�O/l�*R�^�1J(�)���?y�~��2
��
��)n�v�����c� ��U�3��0�$�^R����X!�#�B!0�XG�9Yz���"@P��RG����kwő��pG2�4ڧioh �P�+aL& �G�32::m�ɏu��"<ͧ�?A����λd/p<��A�&j&�yJ�(�!�H= tH�b��9wm�]����L!�D�8"��X�K̍wcLP{%�
 1!�$H�rh���ڪTcҰ��L!�Y�MD2�!��<QI�Ó��C�I��HOQ>I9c��0ΐX�@�,��9ztO�<���ܞ�?1���S�'Z�n��(ֱ$�<xP�eM"��ńȓl!
tѐCһ�RT�ub�a�D�ȓ^����'^�jM4PR!�wB��ȓ������Z�B����y�@Q�ȓ^f�s�N>zb.��f��nD�&�L��$�H]��C�`�z�Hq��F���qB��]B�|R�'=����ŐaT�N=���e��S���ȓ9�Ш{�
1��ӥ�%tKt��ȓ0�t�+2 S�e} �B��$|�ȓoK@�ꆃ�yQ�=�)��i#f����?�S�V*�� �+>6�9��l�'O�S��	�I�����5B����� "QU���O���$�V�����t2�`R�f?[�!�$�'J��!c��+�6�0,͞p�!��A�=SS���F�&�+ClB!�$NO�Ը��Μ(�������#(Fџ�
��	ןxK��j&j@�]�����ׂ�B���O�i�O��$1?ar�����YƦ9L
uӐN�[�<�_bD�`�$��.��%��FX�<a,L�\^2�� jX�k���*���O�<���3iQ�HCș*o��y���M�<	�K�A	F1�dO�;(�P�GKy2�-�S�O������&`��zg��}.�H�+Of}b ��O6��,���C*�v ƓUN8�q���;x!�R�{2)�E�p5
�+"ڜAv!��>���*$L�\*�"MT\�!�$��EYoB�qPܸ�̃�!�D�o��:�LK�����@�@o�'|"?Y��_?�Ǭ��A��PiE ;�uC$n���&�p��q�g�$�q���FO)䂘	UT 
!򄝉V%�Qh�($=Ϊ<S��K5X�!�d"@5hŨ��i��-��BJ�2��B�IqV���EW>J�^K�G\`����$��܈��'q= �Q7�CqP\!:6�+ړP�@F��/�>��%0UFN�M;�L"���)X���'ua~ra�8i�RUZ3'�sv]��:�y�n@9L)�)D�
y 	��	�y"X�$a�=@Fm>t�6,���y�Ϻ&5¡��o�17�IqP���Od)G�MM�_���!l��8�B�-���?���D�����'O�������4]kT���F�X���e�:D�D���C�P`�p-Ͻms�-4D�� ��u	
;n= �'��Q�"�;�"O$��S��)dt�-XC�Ȋ>�py�f"O��#J�g����r������B]����F��$���5?�D "3�ύv؎�(���?�N>�}*��:|n��C�u<
 �P�Dc�<�a�ʌo���uh��f��"�`�<	ˋ9BN>,���EkH�D�T�<�^`،Q�
]-�X��"��M�<Qw ��9��DcU&A�p�����G���O�p"3�OX�1R#�?9_� #'��@��DQ�'%�'�R��>AS�O�0x�����ے4Z�-�n�<�Պ*(�8&nʑ.�z�Zc�<9���4��좳�O,Dm����z�<�􀅂I��DШ�E� �B$Ly��lp�~�&lQ�lW KE�x�mU$���D{�l ����((sҞ^�T�����>b\�L����O��D7�O��r@A��
�^�2%�ƙ(��"O6@��`��;E���ũI d�Z�a"O(,�6ec8�y���
)��Yc�"O�����}a7���\mZh�`��g�џ؛��銙oc���]1+�Bk�27x�	�A�"<�'�?����$��^� ���ۃ/jT`���	�!�N�D�b�߉g�TR@Kfv!�$�=�<�r�D		�0�S��h!�dߎe2�5�&V�{�j�j�τ�I!�� �|�B"ʝ�a�>;Fn��VA�I��HOQ>����:����� .���Qǥ<q`팛�?����S�'�DSq̅{���2�	$�I���nሇ���(��@�a\_�����5T�%M��-�@��4hS�dk�	�ȓtA4	��m	 [�	��$G
kb�݄�V����R� [�eh�aI^�=&�������>�$�3>���w!��^�2ǇS2�b�|��'���%В$2�BH�'^�K���'����ȓy� ��j�X���dÐ(��ȅ�	R��DB�|��X"rT:3N-D����ډS�"����@�j%h��Q�8�Ot8��8Ku$M{�-����	`cA�|�=	�!�b�O��U구� ?����*Y�$D0��'���'㮈	�C ��|1K[�$+
���'���T�ǲq~�� �$HO�)�'�"�:�ꇁ�&<�PJV;��Db
�'����]��PU��IQ������_E�O������]�w������ɣ_2p���"�Dx�O��'��7�I$gC'27�b�D��kB�ɑSDx+C (w��H�%L4f��C�I8i�$(�G�
�p�3G˦`�C�	�"t�V̆�<����N�h�tC�ɖ������/p:L�A�Ȋu��H����|:V��+�߁3�r	IBm~y£��"�'�ɧ�O��=��D ��4kG���a
�'D�49�@�-}��%�F���)[h�h�'k��R3�X�Su|���ԍ4�rL��'���*pil��p N2%n�q��'U�Y��(k�\�zw+�� �֕ K>����/-����`�<�@��;��I `�&TX^�d#�D�O��?�'xջ#@Z�h��AU"i�t�P	�'�v��P!Z�Y&�t����<1����'{LE��N6̬ �ިxlX�'��rNP<�tY�Nޝ�؈k�IYr��2Vz�CCNJT�(�G��hO�a���S�;����`�� #�W�fȢ��I� ��	66�
�b �\�_wT	p� Z5?4B�I8>�m�5&LIGEY�aD�B�)� �u�R�׺_������$,���@Q"O���ʳo�Ș���>�&��f��?�h��-% �CC�R�k©Z�f-���'��ˋ�4�����O0�\��JQ�$$�� ԎҦ A����$(��_.U��=c�&����ȓ[�T���
)�n�qI�B�ԅ�{�B�� �sQ���C'X�P5��\�j����G����$k���'I�"=E���K�p��3���EH:A@�`�.��$��E���OԒOq�����1���k��ГY�{c"Of�5��9"�	[$��?WC�� �"OѹB�H('
�T
 �YO`dp�"Ol�	@�V�^�b0 �y�4A�"OPţ��A�ma8�c��g)�8��|�,>�k�b��s�
�Xa����6{U��4�i��I��ß���O�����Jٲ�"e
Vr!�d̂me�IӢ͆\�u��K
G!�$ �m�У��ڹ�4��-B�S�!�d���5A' �f�lٖM�L�����OEÀ/��S�f�{�ˍ�� (@��ɜ>.�#~��%�>:��DkL���ᕀ���?����0?��n>=j60H&(X¶�2@a�<鱧�FѤ��4��=m0�l:��Z�<ieΜ�}�X��m�;7�4Z&�Y�<1��ܑ Cl�Í��d|R�1��T�'�|�}Z `	9-�nI7��4(*2ȹ��Οl(e )��|���?�O����X�:JE����7���t"OxQ��T�V��NI<'XT��"O,D��b��T+��@�G�1EiP�r2"O����i�%#�Ԁ�3�ҴjN�X�#"O*%)g <v@��h��͠IÒ^��Z���S�5��8� ğh�M�E3l�Hq�I���$Q���1Wi��b�Z,wL�u�w*�;A^�`#Ũy%�O\�$�Ō�C��M�����`�pYN�i>�����T���`�t�v<� �7����c@�Vc��X�A�_��F�O5@0�3d�[E,��סT K������O���.�S o�ʁ�Va:N�d���@B�(��0?!���vyP��;9zt"�JEx���-O���ש�d�JXR`͋!P�z<FW���d�g�@�	[��<i��~��a���5)����H�C����W1��!�9�Ը'-*o���i��N�����ٌ+�q� �?#���6[Bu���m�Hzь8��Q��A9���6���G+�[�,� �h���̟�������\�q�A�G2!眴�w\5]y!�ďA��PK�%w~��j�FZў�
��I��4��Ṓ�sQV��!"^0���O��$�%`�,n�П��	����'SbnY�T~�p�I��eylA�&N�iqT� a�O$�!��.��D�?#<1���8�Rh��������2�5��w��XC��=���O�|i5�^�5�����v	������OR�=ړ�yRa����ӄ'5k5`\���+�y�-T$SSf�6e��a�i �D��?���i>q��a��ݒi�2I!�E�4�|m�	�Fn84��̟&��|��â6:��PD�gJ�Q#[�<��B�]��l�F��֝1 �L�<!�cRw��% ��2-��H�<�^�e�d�S�EƖ6zT0�7��{�<)����%�v�b��E�`9!1,�ty��7�St\<�OxE���8�Y $��7ON=�e�|�'/b�':l}��Y:1p���a'ʙ8��5X�'f�!@g�C�-�1)�8�0�'l8��B�/� �PX�O�z
�'��5��B���0B�R8���-��t�:���֣3n�+�ެ`�,`�c?��|b��~��;�mQ*��Q��v:����x"JS�-�8@��ۀ	9�-8W����y��_ (B��mк\ia���y
� ��ѲG	8q�u�LV$�&�
�"O6�2s.�& N΀�c�37��<J1�	+��
��a⍙z�X�1d��9qH�X�M��OF���O��d*���m����-��fGb��D��Z�"B�ɝ/7�[V�I�"�ME�B��lلP��e��?ϴ̰�!�pY�B�I�yž���	ӱ'�����
8# DC�I� ��	�K�7�jT3�[	����F_�����}"�,3�L�'�/-Z)�7��O�<�o�O���7��A|T�2�ާX�@���E �I��B��U��j@��8iC��*��B�I�P���;V�%�aI���b�jB�	�Py�P��3o/�����p&VB�	=e��HP���"9l�k1n���˓P���$� �#}�n܈n�:� �ê;�D�'P%���?���0<1udH�hJz��a��Pk�@�a�Z{�<����!e�!�e�<|��౓Ë\�<�Q$LB�V
��h���WʄT�<�u(,&�R}�`�ϊ6�̈I�ĎUx�t�)Ot<ad�G'#�M�눛bx-�'R�$�I%��|�`�]o��V�4:^(y�"i���I~�Xf4����AS����)F4��?i۴���\b>��d"�	R>���ЫC�TD	q4?���O 	��>��yB�U�l��i7�f�؋�����Q��p1K��PTF"}b�=�iN�?x}��G�
<Æ�LR8�L�4��'6�>�ɝE���[w-�rޔ�u⇒�,�p$i"}R�'}��5��I��雞���G�Giس���!B�
��C,���i���	���7����/L!�?�o�b�Dc�� ������O3eQ�L#�or	� 3H�ŗ'��MbO��(���§�
�qddS/� �#��Q�B�C\?Y�Wu�T>��9F���D*^����W�H��q�-�"$� ��e�9�򄍴d����X��>��Ȇ�^
��$��i
�9��M�Oh0��'kdMC�O�s�������$_!<
�I�lN�r)x��Ag�O�)z��G��I�!0jFpy�Ն����ȓ�f��um��rVe����q5�plZl��>�>��s���� U3��RRe��1��)�'��'�ў�V$M!m�O���J�d��z
F �ȓiN�=qD-U,�Ǣ�E�1�ȓ[J&�8�ΐR��	�oPG@y�ȓ4���T$�?-�\��f��:C�\t��!�b�TM+�)�q��9N�P��Z0Ν�b��k�*0��g��D���x�l �0,�L�X�R˜<������x*�
��5Jj:|-<5��1�|�@t�|w� j#��sb�ȓr�~��t� Un��i�(Z���ȓz������'E4�@�w ���UF~��'.b�'$��'�`\�SL��?+�+B g���bӜ���ON��O��d�Ob�D�O�D�O��z���p��+d)ה9T\�F���}��ݟ���˟����� ��şP�	ߟ�s�f��32y�񉟥N� ��$DH�M���?���?����?!��?Y���?��@�o� tPZ`^ҽ:���.1N�V�'r�'B��'��'���'�ޫFZ�`4-�xϔ�+cm\�zJ�7��O���O��$�O��$�O���O���J�$TD[ՋȜsADE��CC�?`�HoZʟ�I�|��۟P��ߟ`�	ɟ��Ʉ`����橆�9�,��ǀ�p%��2�4�?���?Y��?y��?���?Y�t��p8�$Pz:����	��4|�U�i�r�'���'B�'�r�'�r�'6��2���$X��/�bt(��"KpӦ�D�O��$�OR���O2��O����O�;�*�)������I�S�|aJA 䦩�	ڟ$��������\�	ݟ ��ߟ@�"�_	@��a��%��.&� T��Ms���?I��?)���?��?���?�(�~��zDXKr� �fÞ$ߛf�'
r�'�"�'�R�'���'7�h��E�^��C��3_�f�{D��r0�7-&?������%�-��9�,џI��v#ނIȼAJ�O�ʓ�?����ArӪ�ɊoF(|��i̺��<�Ef߮U�H���O��Ic}B����Q3��&�O�9�Ğ�[\� Ғ���H���'A�M���x��i>��C
X��N֮u -�u��K�u��Ey��|"�4�SßP� ��9�,��:���.�+4yjI ��dm}��'z�?Ol˧��ы��=�0؛Fǅ�b���'?'�����s�O�)��?��hd��SJ�&EP��]{v�ɪ�����$�<���h��$I?v%��sb2{?�`�&J��$2��>�)OL mX��-��r�ǁA1-)������?��?y��)����4��dh>�*�'�u��Ƒ!�$H�`b� j{(̒T(�hO�D�<����N��ޚ�ʶ��?[� ��pȏ���SJ}�Q�d��v��sTIKr�X�+n|�4%�1:��� W�\�I�����H�Hb�ɽ���oMG*@��S�Пx��ݣ�����I!?�R#�b�ay�P�F��]J���M<�p$'��(��{���>ў'_��d	N��0Y�H
5���k�4��'���?�4c]�a���~�+G�,�@�$L���4�y��'�ڵR'H�?�:vW�P�S�+GMZ�y�h���nFpN���7����������!蟂�$��U,�"� X�	��I��D�|� �i'1O`X�f\��$z� %Pt���|��'���'�9h&�i��iݥYF�־o�|2WA\�4�<Y��2zGl������#bφ�v��|a�g	�(Ū��?9!V��Iȟ��	Y�䁏�K�dq�\>SG��4���_}��'BB�|J?���_� �t��UI�&b�N��Vj��4���f� ɔ'��d�DO?�I>�����(F��b L!�jp ӝ��?���'w^AHŁݼU��<�g�J3~��e�����d����?�gX��۴A X����[�`�B��?u4��i��7M%d��6-`�H���|�.��t�O[Е'�DH*��F	�P����J_20�C�'x�I̟���ޟp�	��T�I\�dJ�s���)"eA��,��n��IП��Iҟp&?��M˜'�&�8��D��AIs�p����O�� ���O����O&-��f�J��s��� K�RW<L
b��m����ɋ >�L"U�Ol�O,˓�?��ک��N�,��%����uP�h��?���?.O~e�'rR�'D��ѐv�8�h#�	'Вq)��Q�[]�OP=�'["�'��'�4)z4�҂<�����֞5����]���F��&��o�=��'PL���<q���j���� 0��x�"��p�	ɟ8�	�lF�T=O���ʝ3&C�� �ăo�<�`�'������¦��?��'t"IR�K�X��D#N�b$X�Q�5�&Dq�:�l��2�|m�e~��ƺL�N��%I`�q�fBɥh70�V��,[(���|Y�l��ϟ8�I⟔����|�gH�_T�h���*LL�
�H�yy2�>I��?1�����?��k�0ee8���ޮS��!���g��Iퟜ�	d�)��xf
�(ȕl���ʀ�¢c~�������*O�h��Ž�~b�|�R�\i��L%ZD! ��}D ����t�Iџ8�Işt�IBy�,�>���D�$o�\i���d>T��B�6�Ē|}2�'e�=O���E��+D����kC*6X:��C��֘�l؀���#�Q>�λ�>]�a�U�HRڌ�k�����<�	�X�I�@��F�O�4�����X<8(`�� )F����?��F���~�4�g�c�P�����  �q��?�:��J?���O��D�OXw �T�y��i�՘58Ӧ�'4vr��g�L)nN���Y�vy�OL�'��@�N��q)oH�y��AO�18pB�'��I,����O��d�O��J���c(@^�@%k��ܺ?GBt�'?z��?�ܴeuɧ��|�qYu�b���J�C��:���oE��O��	���?Q,7���"Bd|AVaUZ���։��sX.���O����O:�$;���<��'� ��'��;����θ	� �C���?��@>���D�O}��''��3���p��yR�P�,����'�RR��ƕ���p������i� D�bi����k�P iT])��^����������l�	����O����6
�}X@(K�e7u$Z9R$[�������p�s��+ٴ�ykԛ'z�h(�(�;&DP�]���i��O�O�]`�i���H�GB���i��Y	Z��+��0HbĘ�+�P��	���'��I�h��>�R�	�5]���Kҭ�>��X�I�������'����?Y��?i�.E;y8�2BϑO�Z	/w����?1T��>Zf�7��w≉GnT��!&ԵAP�$�An�W׺P�'�)��j�20:\I���4�\�R1OLK�,��B�9�j�(R8f�c��'���'���'��>i�n�D�Q�"��L�p�D[am����$�<)ֽi0�O��	Ƃ0 ���/J��(��T ��g��PΦEC�44��ڛ���H�Q���v�D揢1,�X"	�	�\���^N|%�ĕ'^2�'H2�'��'-���#P.IB&P�%X�(��}�U��Of���Ov��(���OD�j�銾N?�|1�-ΌHrt Tj}R�'1�|��Dh�
`@ �4�`B����ң.�] �i���3K�J��G�O��OBʓi�  ��	+Q�dsBX�n���?����?i��|.O�H�'�b� �hB D�.+$�YR#μ����'[�6�%�I����O��$v���E��0#ę��N�?aF���.^6WZ6�$?���J8Q*f�|z�w�beؔ!ݜ/P��G�@�L��J��?Y���?y��?q���.@rd�8x�	���7&�E�F�'C��'����?�Л��	��-9��N���谆D�nr�'���'zC?қƐ����G"dC\����/?ݢ(Ub@�~��I�O|�O���|r��?��V����s����}��-��z� �R���?Q(O`�'T��'�?9��EĖ=�d��G�W^��9`�<�[�X�	П�$��O��zD�?��Q�I�&f�1��o w⤙3�4��D꟔���'�'�$|��h��qּ}�͒HƑ"��'�R�'�b�'��O���&�?���@�'��<2�j�-��ɋ�L�V��<iU�iX�O~��'�����������s�R,A�I���'�]#��i��d�OH=��E!��s��2F��n�H0�1��/1��h+��Fܟ�'���'^��'���'��S�=�D���M�* �EU��'o�������i��vz0�)�	,�A��v��'��'��O��	�&�i���YnDM�BKV��%SEO1��FT�)�fm������4���� M�p���xD\�(��Z�\���O����O�ʓ �����<������_�Bd ��`� �gk��
��Iߟ ��x�I�S�ް�T��V(*��+Z��]�'UX��숚t����3�I��~b9Op9��Y��V�Q��>�~�F�',R�'���'@�>�͓k"H\CЊQЩc��L!O4���I%��$�O�����I�?��'I�hq񦏔j��= Fe8���{�wn�&"r�YmZ,���n��<���dVЁHC�����t��9��G�T���vD��R>��O���?Y���?	��?���7�TՊ@�\�P��1Mɮ!W|#/Oȵ�'@b�'2��t�'��v���I��!2KϊI&���E��>��i�6ͅz�)��Uqra(��]�xkAU���g���rB��"��4�u/�O��cK>�-Oڤ��O6c����rˆ<��P�(�O��D�O^���O���<Q\�,�	������U�����, Ud��	��Mӎ��>9�i�6�Ɵ��[�{W��Y��;V+D1��"�}�7M*?9ń��fAH��?�����#}X,��5�I�d���2���4�I�<���	��F�4��8� ��-�� �0{R,N�?���?)�[���	ݟ���4��' �<�@�ʂT(^�qQ�WFX4��x��'L��O��q��if�	" 2 ��О"���0��������J� B�I`y�O�2�'�"�ד,��Dif��>S��!ׁ�;L_�'��	��d�O����O,�eiF��)M�>�r��
n���'o,��?Q޴v ɧ�I�k�L9p���h6���S�2Nd5�&�PH*Zt��O����!�?�P�&��<^[�53.P�w"����O��1><�D�O��d�OP��:�	�<�$�'cfM��G�jmx�9���[.�j��?��/�����K}�Fl�|���?P<n���)ް� �h��!�ߴ�:�+޴����<\��'��'�ԕh%A�-!:�#�"Ηm64���Hy2�'2�'`��'�r�?a��LQ�PP� �D��815,�Z}��'%��'7��y�i�h��W޽��M\klPd`i��QĶ���OғO6������mӂ�I �PQ`��ثH
nݒ�h)l�d%9̹��'b�'��i>��I�g�@P	��:J�	KEA��>i�I��p�����'D���?���?A0�Y(d0��%�E�J�����I���'�"�D1�6nn�.�&� 㨓�c�������+�j-)�VbyBJÅS�$!!�ȾX��O�"=���X����o&T\y򧊅oL!��EV�sd��'a�'A"��<�Tk��h�xJ��_稡�@#�ٟ��OD�>��v���Ε�v��F�L}���¾;>H(k�J�O���O>�E�~��6M6?�/��˖�N��d�&� \ʉ�Q el�`%���'Y��'�B�'	��'�T
��	͒�q�����`eR� ګO�d�Of��9�9OPК2��*o3`�Q�I.>��`FBm}�'��|��d�� �(���헆w�XƤ0Vd���i����P��O��O@�l��� l@�rM�䉓�N1t��p����?���?����?�)O.��'�b��i��b���'$p�Q%��"'z�|⟀��O�D�O�I'-7$=WGF�c�غ�O��"���Bw���`���É+ʧ�y�O�bP�t�Q#ȵ��u ��?!��?��?)��?1��iC2�h��5��h�Рb��>�"�'����>	,O�lZK�U+�I�Y�P��a�0b�4�%���	П����_��lZk~�FU�:e(9{  T%��J�A�! �~����r?1M>�/O�)�O��d�OT$�wE�	f����POB�(��Y�U��OH�$�<9D^���I۟d��q�dI{��T bdW
o��A��A��D�Q}��'�қ|J?��Ņړp�8���* $��c+^�K\����d����J�ʲ�P'�,�戃�Qm��� ��<nP��#K�t����`�	ןT'?��'���� (�6K�K1����HE"\��'���'��6-(��(��$�O�mg(�G�� �O�OD��UK�O��V�2�6-(?� �'>b?���Ԇ-���z�
�[=��.�OD˓�?I���?���?i����I݀_,@�� !AI~U��Z�k+�듆?y���?yK~�-֛�6O�F�C�ho� ��c��H_ِ�'�B�|����O�*Ms���O,��+����M�7L�9�w�'߮y��i�`?iJ>�,O�I�O�	���Id�Y;�b�Gc���'"�'G�I+��d�O��D�O�1(5��z�U0
\(
w�(�	�����O���4��G\.>hc��;��$J-_><���, ���$�M�O��;�~b<OJ᳑M5<�gH�.BΚ�P��'��'���'��>������6�^%08jLKbeǄ	Rm�	���D�<V�i��O��	^,!�t��H1�v5��KߪQ�����O���O.�`��|�H�Y���ʦ��~���`�J qC�҂V��h��,�C��Cy��'��'^�'^r��'9^�!���:(�V%
Ƥ�7�����O���O����d����+0Ɉ�'��{�a\.���'�"�'�ɧ�O����̑!I����筗.4r��yT႟�1��O���񈀅�?1t	6�$�<��F���	X�I�9DEA�?2��O4�$�O6���O�
��̟,X
̭f�
�K�;7l�x�_ɟ�b޴��'����?��y�*� Up�)�.E�}��Y!V@�A?���ܴ���Xr�Z�O(�O	�.��z`ah�g !!�4� ��ϱ^��'Sb�'���'P��/�h���	."�N�����n)��$�O��d]U}RW�p��4�'H���Մ�zQ��SmK�q�jL>����?q�+�`� �4����.ĘU��?!�>!j
ۅ�DavC�>B��	i��`yR�'.r�'�bA�'T����&d�=h���w�	(M���'�$����O,�$�O��$~&�1��8��qCW xm�'M꓄?����S��I�! ��ɶ�Ut���Q���?w���rΔ�o��֞���ӰS��?��؇][f�8�ˏ%h߀�$L�9�6��O��$�Od�$'�ɼ<���'�t��0���b�#%ە� dj���D�Ԧ	�?�#U������[�"G1������?����	�@V��֦��'˖=��!�M���U�0�L�%x�Yi%��CǞ,��Tyr�'x��'q��'t��?�c� *< ����I�SU�(	��u}��'O"�'j��y�ei��扤e�CG�
�qK����D�(���D�O��O����iK��k�J�	 �<� #�S�.��I�t�Ɇ[s���S	�x���'O�'��i>-�I"k�}��(ܣ��b����@����l�I���'���?)���?�fD�$5o�Q�fT�,$�2ę��'D��Um���m�D�&��ٲ��	1&	P�iER|2����wyr@Q���Ѝ�6��4�6�!��h`��I�o�����@%@%x�
�d�OH�d�O"�D;ڧ�y��9Fn`
�)�56�,SdL$�?A�U����؟��ٴ��'�����Xo�A��+�JC�(��O�@���'[�`Ӑ��y�h�$ ����G�����q�̝�#S�}/<�Pw�,t���O0ʓ�?Q��?����?���y)lӵCd_<�P��<�R��.O��'z��'������'�P��c���F�B� �J��x��,�>�'�i/�7�\�)�S W�����	�nc����,��T]BB�)�2N���������O !�N>�,O�m��ب>aj�a��ۣ\;b��&�O2���O"�D�O���<��[���"^����p&ɷܶl����4���I8�M�2/�>���?���'�ԡ��^,"�%��M�]�\P����M��Opђr!U9�ҏ��;��z2��,�V���\������'�"�'��'�B�'�>h�hжA�B�����K�V���L�O�D�O���'�R�'3d6M*�� vz����Cf L��I&�@��4~���OXP��c�i�i�����|\�{��Ċ
}v��v& NB%���2L�OF��|��?���F�ڌA�ᆈIR,�����l��}r���?�-O8��'�"�'1�?y�p&'�&4	��j�Q3��<	�T���I۟�&��O�zy�C�B$KN̹�`���k�]��=�s�릭�'�$`M?�H>b�!*iڥa2,����!Ô�?����?��?�J~(O6L�	��2)�	2�������*x��D�Od��̦-�?Q2S�(���0�;������A����?��)i���4����2���+��Dc��֭�%���@�C����?�(O0�d�O��$�O8�d�O��'��}Kā�*R�X! ���Eu} �OP�$�ON�D*��/�MӚ'BF틆�T�gl�q��!Pݨt���?9N>J~�Y<�M��'�z��נ��"�p)p%�E�${�z6�Z�k��,&�(���t�'�Tܑ�
��C��Ӡ�q���F�'��'5X�T�Ol���O������8A�O�Y	&��W�1-�㟈K�O~�l�/�M��x�/К91����+�C��;�n���ɮ��;hs����d�������;O�4�EG����Y�GR�C�N���'�';B�'��>��S�? i�d)E+T�.A�������C��'�6ꓷ��M�?���iP��͗Z�|8c�/�y-X1P��oQ�V�|Ӝ�o��pPn�M~���"$�\��S���U�E�#ADT���̭=I2��|�]����͟����8�������H�u��}���F�\T��h©Hy���>�)O���2��>	�(<2�.V�LB8��)��&w�$��O�`n��Mc��x���K�&�xh`H^�l��鸁�� IM��R%�Ǉ$��	;&$A9W�'�&�L�'��H�%m������-/":툡�'�b�'���'�b^��Z�Ov�$܂�Np�Ɛ1�p!���:�b�$G��9�?Y�]�`K�47u�6+�O�� W�_@�%jaD��8��Mqa/�=Vu���H��ř+:�Ā�R�߼���Jb����	QP��2& �����	ܟ��I��D�I��E�����mkQ��< ,��$"��?���?!�T���	Ɵ� ۴��'�><��%٧Z*=�d��AU2�PL>����?I��AvR8��4�����<��̘ L����dM��q'F��`��JɈ��d�	dy"�'���'�2�:_���viǒ�� ��K�.�R�'��I���$�O��$�Oh� �L-�Qb�=б*�Cbݦ��'l���?����S�����k6�<T��ɳ� v�e��W5u����<�������_�	�Mߌ�
�H�4�(����z�J����T�	�h��Q�Sby" �O�u	�$��1w�`*��b�H��'H�Ƀ�M+���>�Ҽi���/��=%�	r��9{��P8�o���m�2k*Pm�|~�o�=;���8{����
@�l� ��y�a �mU�V)��$�<����?����?q��?ϟ��3�ܴ%�8\B7�\@���>���?������<qհi��D�;�fi��Zf�̀���'�6�즉kN<9�'�R�'@^����4�y��������Y�0J��!eB��B��s����R-�'r�	˟P�	�=��]��KY'7*��!T�8�Iԟ$��ϟ@�'@��?����?��F4��4Z� Q�x��P�K��'�R��?qشz�'�i�^nB�5��/ƙDe`	�-O�	� ��j���u���Ӊ(���<1V�Хy�C���ɒ�0���$�����Iǟ�F�d:O���CeUC���q��X9y��'2���d�ӦE�?���#^��K�7�X����
����?���?��oZ�M#�'�2ş�.	�O�`���Q/t�T�:5��6Up	ZL>1-O�$�O����O��d�O���-� K���ag]7zT��0.�<1Q���'�"��4�'ۘ��f�=b�Z,���\�>L�6��>!²ij�7��`�)���L�g��䂈 g�ۢ3�Tm�6cU�y�F�Gg<�2��O,��H>*O&�:�a8BN�C7��,|Ƞ�q��O�D�O��$�OJ�ĵ<��[����*1��	���=~��!&�@�`��ɶ�M;���>Ie�i�7�؟ "9J�&�rK� j�hvn�#Ow07�4?����9i����3���J��drތ���|X`uG��l�	͟��I��@�	ßD�� 	"S�0'�D�<g��`释�?!���?�QU���I�Л�4��'�$�d���Ax�E91�&K��J`�|�i=�6M韲�cVMyӨ� ���&V�rP�4��0-V~�	��=n9�{U�'�X'�������'��'L�*��>�^`�%��K���r�'�[��J�Oʓ�?1ϟ�	( H#K�Pe�q�U/uܲ�`aV�hK�O����O(�O�'&��P�)ɍ9��F�3z`�a��@Ԡ��1c<?y�' %��$�8��"�\e �I�|Gb���B�>=������?Y��?����'��$�������܈2`�zV���_ĝJ�l�O����O��<���O�ʓ�?(�
��a`s훿Xv�ɹ�,�9�?9��H��#ٴ�y֟ac�����.O.p�E햤NjA)�AM+E��ن��Od���O����O��d�O"�D�O��'v�&��v���V�9��M�
r�@�O���O:��*�9O��j���V�]��,��K-}�I�5��O����<��?���?Q�=�M3�'2���B�+Y���GQ�Iovx���'/� �5��{b�|b��t�')"@�4&5 U�Q8F0l�W拭S^r�'<"�'K���d�O����O�|����p6�I�l�|�0��)��Ny��'��T�DΧN� �aT��MX5�IEj'n���ɟ\ۄ��py�0l������ʄ��':��3uº��BԬr"�|å�1+��'t��'b��<��>�z�+�b���XP�K��$q�OT���O(alZS��jb�܅�x8Stƃ��m����?��?q�/��a�4����@�ᯤ?-�6�j����w���.-a��Te��EyB�'��'C2�'�K�P��QT!܄B$�%�TcB�	{�	���$�O��$�O8����D�8ʴ�Q�B��)�D8��&F�(u�8�'�"�'2ɧ�O��	VA�9�����I��w�� a�=��v�<�g�݀j���i�Gyr
Ɏ������H�x�Gպ|��'\��'��'��	����O�e1��-w����.ľR�ʀd��O��ny��o��I؟��	�<i�J	e�48a��R�~�� ��9.�m�G~�'(��'��'�y�I�
n��aOG�s�z@c��K��?���?����?���?���� V�b��44�HeQ芆�=�'��'�����d]��<�`/<�����>���8to�x�	֟��	��ܢ4�˦�̓�?Y�̎O��dC��};R��A�҇K���5L���'�䖧���'���'�`��!i1P�@ ũ_7}j8��'�BP��p�O�˓�?˟NY� �D�6�q5ɒuaJ`�"]�ӬO�D�O��O�'2���Z ��){=��� ���b-�m#�[� �oZW~��O�<(����O�R< ��iI��ܒ#��q��ɟ��	��x��̟�%?1�'#x���<I ������� R*mMP���۴��'����?	5`�,�0��D˯saTC���?��Y!�%��4���+?;~������#���pB�A.鲼��$�?*OR�D�O����O4���O��Q��a�".&��0ӂI�=0劬Or��?я�4Ao���ɢZ�4u��C�" �&�AÐ�L���D�O��Oⓟ�I@z� ��;@��beơ&����6���d�.V&Z�'q�'�i>��	�~��!gH�'^�p8��ׇ'����ş8����d�'R�꓀?����?���ߔ@��x{��@��TyQ"���'=H� ��� w�&�3G��*vx�Y5	��H0�S�AyrgU|&��#be�O ��Ie���P��B�Q줱�&�۲j��'���'���<)����{�<����7Aa<EZ����+�O��uěv����mAĕ�DO�#��#+���C��O��lڳ�M��ib�9��i��I4G�vez�O����a�r�蹓C��#���B6�D^��iy��'���'�B�'X�j��z��Q�$\�?�LX���(/l剃���O����O����$Y�e^���bJ	5��1I�M�(Qp� �'�6�KӦaM<�'����~|)1e!���a�7� l�Pm�a�
Y��)O�ɒ��D��?�# &�D�<�j�"*˲�a�۲Ku�S2挝�?����?����?�����Q}��'}PH�3�l�R��u�W�j��H�'�6-3�������O���o�$#�k�,C�mԫ��Y"���%x�66m7?igImӐ����䧲yGO�?	�pzV�8K�:�س.U�?����?9���?���?���וZd �ȁ��	'V|�c��v;�I���ɨO~���O4En�X̓OGb!X`�7&m>�@q�Q'5�$�,�I����� w�2n�f~Zw)b(�/H�v�֥$��P�H*$� r��,���<	��?���?�����!��u����8��9�b��?����D�G}��'{��'���1w��9+'�-?��+A.S*y4�ʓ��I����It�)�4��C��(s�_�v~rQhd��b3$���X:�M�W^��ӅO���=�D�\��(�JT��{cgY,����O8�$�O��*�	�<���'pF�0Ca")�Ф˗c�C��ٳ��?��q8�6�^N}b�'"Pq�)�|�~�1m�<h~|��"�'��
��V���]|�|��'��IFh��l�%�~�j���,��F���<���?���?����?�˟>�p�iܧ,�᳡�U(kf�D@歵>y���?Q����?�3�i��$��X�~�"dva�h]��� � �'&�,6�2�Iܟ�7��<ж�Յ �JEBUbP1 F)�т�OZ]�P�֤�?�@4�$�<ͧ�?�5���76 �P
�Ѝ����?���?���BL}�'���'V���ք�6�hA��22&����D}��'	r�$�� >���0��2y;2�QiA���7�P�@E�<+<����iJ��D �<O�����6nI��Ԛw/xX��')��';��'��>�Γ&��hR-���tF�1���I����O8�dʦ��?I�'3�����O�[������ɭ?̝���?��\+�ƨǿΛƒ��Zq�V���T��F��E���sRH����G�X�:%�|�_���	��|�����şd�F���^�Ly��Y>kؠ��-jyb��>Q��?������<!��
�qq�uq%�)�r�����,O�I(�M�v�isPO1��$s����/�ع��aP)A����gψ2&�Вϼ<ir���/q���K������N8Lp�'D�PP�C@Ո\��$�O����O����Opʓ8��	ן舣/WR�p�Q��
K|�DÓ���X(�4��'H��?����yre��j����<��	�;-4�lX�4��X&w�Y��	}�e�%��Xn@���m�lq�$�O����O��$�OZ���O�#|��C)G�t� ��;y�q��g��	��+�O�˓G���.6���Ξ2r|�zs� 2sa�'�r�'j�N��8����!�K�c&f��d�I�8�˞�\Z�D1�O(�O���|���?A��[M�q�5OV�v��0"a�Β�� ���?�-O���'���'-�?-��@�YM!p��6K��ؠ'�<��P�P�I֟�%��O�x����b��MЗ�U#?�~QS�N��8VT�0�4��I�?��O��O��rU��J6����6S���@���O��d�OX���Oj����x���x
9�0�?�8��S��?�/O�dl�s��;������T|�,8&AƁH# �b�����ɖ���mZe~Zw�, џp�'A������#��*k��	@yr�'�"�'Z��'���?� *PI�._�&����]�X�6I�s�>����?������?I��i��d�:;�
���_�&���@R*��R�'��'p"�'��.�,(��2O�Őd��>edj);b֎N�� J���O
�#E&ײ�~�|�[���ן(��Ć>4��7��#x�Tl��ğ(�	��x�	uy��>�,O<�$�78/�y���*1pg.�6"Y�㟬ۮỎm���MS�xb]0"p"��e,R�43���ȈH�剰Hw�@��:#S*�'?)�v�'V*��JR攚b�';!x���Q�C�,�	�����p��b�O��2KQ�m8@��
j�J�JQ��;fb��>�.O��nE��� �W
r,�En�2$=a,�.�?y��?a��MY��Bٴ���a�h#�'�u'�ߧ�P)��x��=p �I������O����Op���O�����YZAȥj��9��u�D,��fo�������������%?����!it0&^VuC�M<U��}�O����O�O1��̓�G � �h��<�J�W6�T��i���5 \�b�O�Or� 0ms�D`��,+rF݉@XM���?����?����?!(O�T�'� ]%_¥8��$F�j	I�N�=�b|Ӟ�P	�O"���O��	"QR>D�g�h�fa�`�/9@�n���Y��0�(4ʧ�y7&�R,��8�o�LV�1�+E!�?!���?���?)��?A��)��sq(� EM /h��a��yR�'�bư>1-O��o�Z��֑!R'� %,��e@H���`&�0�I�p�ɌZ��o�D~�įupN��wO�3��c�#�/~J�X������03�|�]��ܟ,����JaFP}0��z4`�����	Ry�ĳ>!��?������ͅlO��HC��[ڳ/��eS剽��d�O&�d)��~�d/�@n��%�
����Æ�L�M�­�'E�^X��.<��DJ���?ܽ��
N���	���`����?Y���?����'��$UßqƁ���~5p��B�?Q�4I�c�O�ʓ���dC|}2�'�݉���0�왙�@�:wRj%2V�'�2&O\e����(�A)��{c���D+D$#u�+`��MU@2��>�?*O6�$�OH���OF���O �5P� �`ŹG�@���-�� ɪO����OL��!�9OpimZ�<y��W�2<��,� �|��6m��4��r�	T�o��l�q?1��p���"��E~|�:「ϟ�i���{.B�Gm�Iy�O��ǼZ�m�q��F�hXS�˦V���'��'=��3��d�O~��O1�&پ))̑x��@$m� ��M"����$���+�4��'� �icE�([t#�ᇉSfZ��gU�|Ё��5F-hU�W�S;4���<�흴"0䙫��݀c��+@���,���h����F�D:O��Ϛ?�v����@�c�\���'�����Pզ��?��'^�E	��RV���}�@�&�?	��i��7M��a��x��U~�g��>�Ν�Ӣ(k�5�@��$2M[� ��,�N�і|�P���	ݟ4��ҟL�	˟���kP�q`Ҵ F)��uA�]y��>����?�����<��H�F�z��Q&U]�X���1*��+�MSƵi��O1��	�ɏz�K�ɟ1(tJMxs��9����� �<	5�޵nD��������d(#�h�2�ĀXQ�ha���Xy.���Ov���Ol���O��t��ӟ�颩A�wn�`CC�ߑ}�ظ.P����)�M��B�>9��?�'��9�U"T�Y�Xhq���x]F%3 ��*�M#�O�u)�L�3�(����Y�tkA�F4)T> �g@�s�X���O��D�Oj�$�O�$/§��5�
^
���4/��l��(�����ɟ���<YQ�ix1OZ����!"tf=�6O�2s���*P�%�d�ަa�޴���f���M��O���1�^�/9�,�8�XP*R2�~����h �Oz��?A���?��5�Z��b�7�%Ҳ��8A�0Y*��?1(O��'�B�'Q2�?M����+�R�z�KԤ;D���'�<��[�X�IʟP'��O��Tۦ*�"-�|<%�S4����r	L5)r�}B�4���럾�y�'��']�\(4I�<{�9 �I�SN����'�R�'���'��O�剹�?a�B�8�}��#��"�K��e,��O<��ѦI�?�ST�X�	�3	�Ѩ�8��p3� ;O�0��`#g�Ӧ�'z�j��N�PJ�#c�)s��9oB�%��yyr�'�"�'���'�?��޲�eDV�@���B>`Z���?���?�H~���1O�A{��B)~^j5e��9{z�p��'9��|���4b�5'���O�Ղ�X�Z�jA���Ƃ/��	�f�'�����Vş��|�^���㟤�S�@[~�e�
e��d�R���0�	����iy�l�>����?a�E��pi�L�r�L( 1���U"��#�>i��?I>if�1LslSW#�= oZܠè�&��]�l� �V' �W��i>eH �'�<e��A_�0)E�hp��/_1P8^�$�O���O���!ڧ�ybH٢Ԗ(��h�ȼ����?Ic^� �'37-�I�?�I��D�x�XM5�B3p>Y%�[������$�I7I�n�H~��O�D��к,�D����'/�ܢp�_O��ny��'K��'��'�� � s�ƊB= ��L�/�\��R���Oj�D�O�� �9O*|H!O�j�X��fDE����wC�G}��'��|��T�	�`hipt�D�xW�܂ԇ۩IL@�Kƺi���n�&�	�O,�O�ʓ��P0�$^6@>]h�b,I��E����?9���?���?+Oi�'�b���^�����"M��:&��#__�n}����S�O��D�O���u��jA�=%+(-�5CA���K�e�*�t@���'�'�ywE��`	�Z.F���O�E���	$�I֟��	؟\�	\�O��%1�o�/w���q�, ������?9��;U�INy��y��b�y�D�U�����F�#� �1�0���O��d�O���&s���DER,	��30^5�RB�$&9� ��Z���IT��Fy�Opb�''��^��#���}L��4#�98���'�剝��d�O����O`�'=���`�G��J���h�"��Z̗'�(��?�����S��F��i�%�1L)bk$b��\�n�ڡ+Ԇ`���)�<i�'Y�2�	J�I-Z|����4HPh��Ŧ0��ʟP��ҟ���B��@y��OXA�	�c��Q�2f�HC��'��	9�Ms�b��>��i�03`˫l��``I�90��qB���?����M�O���J_&��O
�D����H!���9-��D����O$�d�O��d�O��d"*0e� OuB(��B� G��x�$����d�O
���Ox���ćæ��N���!���7��1�x����<&��$?��˜٦���=�NA�'ʺ)
*(A�	�
}��T�(���O2�O���|��,tp��I�T�|�P��5Yv!���?���?i-Oڰ�']��'�"�G�J���[s���X �:q��Odq�'���'��'����E�c��QV�����%��\�h��F-�=nZO~�O�z���yd� hLȴ� LיA0�	;�H��?1���?���?����x��Q�,S�4���]�V�@^���>����?Qu�i��Op��Q�f���bP����+@��
7T���O����O6�`�z�2�Ӻ[CM���D�̺s�Z�a�6s�\�+$��Q=�'��	ϟ��I�x�	��I?DqD�*C�S2h�-)NL�'�*��?����?���4(�y�JT*ׄ{�����J0��?��S���O ��BD.��X���FS�IT�;ϐD��� �+��gpBe�myR)�yd(t0�"2E�Nћ7���*��'n��'��'}�ɢ��d�O�|*�f�X^�Z1��>;fH]ZĎ�O
To�Y�����㟐�	�<��Z�j=��ɾH�t=�쓞L2��n�b~Ҩ�O���Fܧ�y���gUD`D���sy6i'	�?q��?9��?Q��?a��iH�T�^fg<|�Ě��׭rb�'z�c�>�(O�(lZN�l�����.|�Pk�N4<
&$�P�	ԟ�IBUoQ~ �m���Џ��wdv�["��~#J�A�ޟ xW�|�Q��ܟ��˟t����	f���N���BMG����Vy���>9��?�����AY`N��p�Ǘ4�(��A�b��I�����æ1h�44%���Ӣ)��Nֵi������"E)���M�K���?���'>��'��e��C� 鐉�[~�ht������۟���t'?A�'� ��!J�v��A�t+
��-ș���'�"�`Ӱ㟀((OJ�D�,xi:�C�L��nb�e�"E�Ţ7-��%��V��m�'d>�A'-H�?M'>��%��P����͗	~�$��wL�O`˓�?i��?y��?����9�@�S�E�K��u���$���?1��?�J~:����5O\��0F˄o�P@���Y�x� ��eӆam��ē��CzH1�ش�~b�� �|�	�.`�B���S�?!���7���d(�䓜�4���d@uB\�� �����>�j���O~�D�O�h��IRy��'�d��Q�M)a���q$Z�9���"����p}R�m��mړ�ēB�*�#"$](*O6U���O�f�Ze�,O�<P�Y�EH��:ő��51�Ҋ�<Q#��$[���B\�2��L"զß��Iԟ$����E�t3O6��@ty��C�螟�5#�'�h��?���-��F�$��iH Ӄ#�fa�QC�F�~9�&�e�0��֦A��4̜H�4����7�L5����u�]�Yn4����� � ,e�5�䓁��O���Op�$�OL�D��b�����'��	�?�4ʓ^����x�I㟤%?q�	�`
���M�*� �pIط{b��O��l��M�V�x��$@S�eA�#C�&��P-�62�h��Д��Z� "T4���,M`�OVʓX��z�䂐\���7oC�(��U���?���?����?y.O��'��,�6Bό�y���u��=�����R�b�x�P�3�ObHo��M6�'#P�����O��Є*�<2�{�.�M[�O�p����z���:��=P%�N�����)O��QQ�'#R�'y��'&"�'G>ia�ɡZ���3��#P��!�$��O���OR��'��'��7%�+�Ƞ��N5���oM�9e�O>�d�O��	:��7M<?�'�5��K��5�0�5
���᯼��$�����D�'u��':� �QQ���^�,l�Ų[=��s�'�\�ࡩO6��?�ɟ$�3�!�*w��XcF�S: -H�I4\�d۫OZ�d�O&�O�'X㚑Kc�+`E��)�I�P��i�լ�~���l�V~�O��������%Cݚ4������b`i��?���?����'��$Fȟ�Pt���"`BZ=v��bE�:�5�4�?!��6��&��}��'� �I��"lw�kՉ=5�4i��'N�#̠I�旟֝9lx�������TL~E�H��I@$��T�\��ߟ���ܟ��I�t�OVD��g%LLI`��N!�|h�AV�8�I�,��^�s�@�ߴ�yRk��"@��J&-��Q[�C ��?)��䓳�AT��cߴ�~"��d�r-v��=I45�"(��?Y���d�H�	T�Isy�'&"���`d1���/:�h6H�YGR�'��'��	�����O����ON���e�>az0$�T<�i�,'�ɱ��d�O��D9�dɷ/k$=B�I_�O`�tJ1K�<�hʓ|�⁹bȺ�M�Ǔ��+DP?��'��x�R@@�(����$@�\.b��?Y��?��h�b� h�D�K�O�܌0S�¹X��
z}�V�ܚ۴��'��T�H)e� 	�%^jڑs��	�R�'���'f�#�i�i�)rΝIj��M'Z�2��`��[�����CC$�Od˓�?y���?I���?A��w���zK�TH�h �K�i�A�*O���'��џ�&?Q�I�����ըDZh���&~Pi��OF�D�OX�O1���HB�)l���3�Bf���IC�M��7-�Qyr���M`e��䓊��	���Q��%�=�lY[d�$L���O��D�O����O�˓g���֟,�iW�Q�F��@`I��$dv��ϟ�ݴ��'dF��?���y��V?�p,������}�b��$w��R�4���5P�p,��O��O7��χ `T��C.�
g_�l�׌�xx���;�Z7��;f���1��
t|���-�{g�̃V���!��c�h�9���7k¨�$�"6Œ���Ԛ)�xXr���{}�؂���w��3��+S�X&�7�*�9�������V�z@|hб*R����:����w�UFG�	�J5��+����	�'S�nh,Ȑ0(Y�=�Z��#���uS`���H�h����E<x����Jz�(e	  4�@�G���A�%U�\�80��F�):IT��w/>�d��`jcP�yf���T ��1�̟v�p��&�'@�J\���O��ǣ�԰Z���o�X��5��
|&4�bV�F,�,����d�O����O����<	��cJ$�gM�2]��+TA�M�T�u�M�'�)i�j��<+
U�wfz����ɒ�H�>l�$2j�&%�2�V)��}C��;d���P'$oRu12�Ӣ]O���E��U{��]���K�H\Iv���P�I�fҬ-���Ex��<8�����(
��O PO��#�H�&�kd�
8$A���v ��s�Pb���ҥ�~*���fR
S�����")�}@d��Jx�@�ę�df(x��:4޴X�m��3�>j���H� ��#�H�{�n��Nλ:� ���"�~�a$K	7�?Q��i�T��DZ�Q�9��5
���g�'���ڟ�$�@��ڟ��%춟�Y$�"�yRrŗ�e}Dd���<���?9���'+������P�^�!	��J�����៌��Z�ៈ���O���<��#ȷ!�9�'�h�ԔG��ݟ,�I���'Gr�~���?9���0��
�D<�@����@�JH>���?��߃�?iL>Q�O��kV�̄^^��&�F�W��B����O�Qm��� �	�Ɋ����L�����B��1FڗZ����O���Ħ|.���:�<�VN�	�"}k,I�p�����O@ n̟0���\�	���$�<����w�,M:E-��r�@V��-�?�fkí��'�����;y	���G
$�9����K9t�oZ�����������d�<a���y�o�5f� 9J ��~������?iN>��փ���?���y��G���w��	�д)��?q���?�GP� �'��|�HF)9��������r��ĸ,�	*D�*`&���	����^��%�<�K�*8*��1эG�@H���9��$�<������?��*���o�9W0���&��.$��f,�A̓�?q���?yM~�Q�O�:�꓆X�&�� ��240�1����O��Of�$�O�8�Ct�[�BTC.0�DeE"�:Y���<9���?�����aB�S�DH�ɨe5��3�ǎAbbq�Kʟ���s�	ʟ��	�~;���I`~⃘.`���%">���i�I��<9��?i)O&��E���'2�'��QA�,�y9����K�v_�M)W�|�'^���v��O�!rL@���N�LY��pA���+5���<���P��V�'#B�'{�f�>1a'w�¼�D�4w(�����?y���?鐎����'�1��ᒥ��:/8��$��a�
̺��'��s�~�$�O6�d�Op&��S;�"�c i�j8��X,=���D�ON���O��O�s����l�޽Ju��&=�i��'�/#� U�޴�?���?���>؉���o�$A�]�/���! ��V8��H`�O��d/�ĭ|Γ�?9��?i7`W�.>8�b��*u�����?����?��xʟ�O0�[��R�w��}�t�Ų�T �f<��O��O&��<�'L>�0� W7g*���iس-~�Uq����D�O���5�IП�Γu�
��5.٪
`���YX����#lb�(��[ybV���g�? 8�(�_J0���t�ۿP Pʦ�'ar�'��Ol��<)0��0��1@ng��ڱm�.	��`YO>�����<�)���䁓G�����v�r�SeO�/����1�Iޟ4�'�TIH�D�Rp������AR���)�O4���<�.O��'�?����~G�ߌ)f�X9�dW�E�H)ӓJ�[�	�,�'�Xe���dF5!���e'�Bh�9?��Q���O�ʓ�?q&�iT���������D4T�^�k'*3��j��:��Z���I�4'?�&?�:%�C:c&2B劫���:ã�ky�'���'���'��)B��W�&�d�"cS��, "�Ċ0��DU32f�"|z`%Y	X0�ځ.��PKȁd����ȟ������`yʟ�T���@�&k�B�)�aļ�$m�b.���'�?A��?��1W���02Ŋ�v-�[G�P��?a��?)��xʟ�O^�� �E�8%t�b�,.��7�!���OX��?	��?iɟ��ٗ.� F���A�A�����'�O��O�Oʓ ��"'� 5�!�w�aZ�2��?YI>�����<9�O��e��lƇk��#��)Wv����?	����'�B\�p� �2PL�Ty�Hq����T&�*F�Z��'Tb�'������3�Ju3�r,ӣ}�(��0��,#��d�O4�O���|�����)��^�l�r�Q�4wĢ��̱L��'�bW�8����ħ�?q�w���jrBB%��hѕ��/\��0J>�-O��d�OF���!�q�3M�-5p=:�,/(�6��<��5��6T>������-Or�+ǪOk�0��w�#RL0��'��	����	_�u��"��	[�%G	���0"�T��e�	��`
ٴ�?Q��?��0"�IHy���g�I��MI+4VU0ao��>Y�!˻���<Q���'�@	k��I�p�:B"G;H���ZjtӨ��OJ�$�O���'��	�,�Ff@�𱊈f�p5��?SEV�	˟0�'��5!��t�'���'(��Q�,�Dl� ��s�����')��'������O�˓�y��	�/�4�{ #��@q����+A"��D�+ca�	ȟ���ϟh��ey��ad�}˶,C�3~R ��eB8Qi�)�>�+O��<���?I�|ULdJ��Hg8����!'b�����<y���?����?�,���'%������ s'R�N-2U�2f��?�(O��$�<����?���0o���>���B�?� �'a� `����?1���?�����4�&D�O]�6j�xօ�]�LDr�a�f��'N��ǟ��I���q6��`BfH`�A�@VL�K��Їt� �Iן��Izy��'���?����?���O<�CG�N�m���g
���$�O~���O��W5O֓Ol擅f�%���>W@4[�&T���d�<��-ƛ&�'���'�2��>Y�g�(U<�`��`����rvkؓ�?Y��?�RF�i~�Z���|�3�D�	�:���+����..A���O�o�������P�������<�5�@X�f:A�<k��%�E����?!����<����d6��؟�����y<}#�"��*BB2Q!D��M����?���?IbQ�|�'��5O���@
H�=0A�>!�'�'���3����'�"�'��*J��p�09{R�O�S~�����'�"�'�����d�O\˓�ywHB�"��P;�O��K�4P�i�;��ރd �D�O����O����O&˓"WX�_3-+v���bY�>? %��m���|y��'������IΟdof��E/6N��A՞&�"!�,3�ПH�I��&?�:��A[l@����|	��1�� �	vy2�'c�I�������@�ki�@��뎬I��̃��խ°�Q�"�Qy�'�"�'F�	��|AI|��MӽI`lItjC�R\ M�𣑢�?�����?���C�*��=��` ?6*!�G��u�j�������ßL�'���/���OT�Ҩq8�ˇ.���DْL��K���O��d�OX�ᥧ�O�O���(�J� �ڷ��ո�cL�r
���<I�^6�VS>U�I��)O���Z�{�PBmS�� ْ�'�"�'!LY`��:�S$	S���D� 4��e�Ǆ�*��$�OnMoZ����ß�����'�~��E#im�$#��4IJ�eJ�'S6�Z��'��'Q����Պ�e.]s5��B����EN�p�i�r�'��'��O�D�O��r<��1!c�nR�ٛ��&,����*�DU��쒟����O����5�u��mL�+�J�IS�E?����O���[��?aN>i�' �<����� �e�h�h������X~$�<���?��4% c,��`.V�3d���3���?��x��'��|��'�B�V�EU �����B`d�)���'l��*D�'��Iן���ڟ�'?����pŸrLGu��� tiȖ%�8�'l��'J�	̟��	ӟ@�SHb�Ԙ��ՂW�t$���P~洀+�doy��'u��'��O���l�f��s6ĕc��Ź�����O�d>���O��q�Z�8?!W.N���R
܇�d9e�]��l�	��x�'��(&�	�Ov��.� ���H)_[b�%9Fi�R�|r�'82��>�y��|B<�R$2�(�*O�.!c X�a���'��	��|ش���O���D@y�%'��E�D:z ���� ���?y���?����<YH>���T(�� �#��ۙh�V���=�?��KX�6�'C��'y�f+��O0�¢�H6!�����&�V�N|��O��HP8O<�O��?A�I6��!agN&$+f� 㙈y,��{۴�?���?�l�OF�$a�4��j�l+,@����C��x���O��O�1"�3�i�O2���O�A��߄_���J���!O$m�T��O����O�&���Y�'j�9���X^��{C4R���L>�����D�O@�D�O8�'v	�Z �C'=~��d���R3���	�ē�?Y��D}�h��5
N�Kr��Sr.�P��OP��<����?i���?�.���$�F�t ��A!��� ��y8p���O��O2�O�$�<92Bι#&(	ڕ��xdhu	I��,O����O��d3�i	M���'����)�phq��*%�"�'aR�'��O��3�	�V� ���ú-w
U�#!O_��D�O����O����Oʧ�?����?� �I@
3��V:W����F��䓺?�/O��ҧቤ'���q��`	䵹���wCZQ��韜�	ٟ��I㟌�����zyr
<p+Rl��mB/7jp��:���'��I��#<��J%�U�;ad�Qq��K�'�B+v�|�d�O����O���'��0c�qi�&�<�D[T-¯g�r�DR%ZS�㟐�~�	�h��� �@`��݈uؖ�K��\�l�Iǟ������֟d�O�29O�8��R�V�(H��B=<�f��$^5�Ofc?�%��[X �g̷{"�8p7
��w��م�.e�,���H f�TE��lS�Q1z��'��?���?���y�i->�v0�W�+u�X葤#Ӎ�?q���?Y�4�?��P>��	��`�'��X�!ϗ?��2��^$O���7���0Y���,}R�5Rdώ$i?�	p���+4�<rf�[.Sڴ�2���	˔	z��t�ȡJ��*l<J���˗�M6���J�"�b�"��)�$i����`՘
� p:H:rȐ����sG��;L�KV�@O�ਡm�%Bn��e\�n�P0�	� ���%��1d�u�׋Gw�@� o�/V�ށ�S-�_���0��D;rt��8�j5����
yNC�Ά9��!��/�Kٖ�&�C5nL�xCh!W��b�[��4eͅ7:�rM�p售'�����*N���	��X��zy��'�b�i�4˄JE�.LĜI5��ݛ�4J���6�M� ��T�`F\'�p<�"�T��<P��V�+0E�#�	����QDT�4�nIK�AL�>���	�Q��I�'.Rh�b�L�}bt7��4J���'eў�%��QG��>U�T�Íz<�P,�\C��+ � l)��!�d���&H8R�r�<�V�t�'v2�����0k�K��e��:���5<pHsqj3�?�������O��$s>�@�B�+���ԴA)���@�>�UpsN��%ۓ"&mص�Ĩ7!��@���<��ٹ�ץm��f��-�a{"��?���M�CU�gEp�tKW.6bx���b�E�'+ay`�y���ӊ�1,�\�S��3�yB���Y�.w��ԉ�-Р�t��'X�*H�^��O���$�
�4zt�ˇ�$���A�Q?g���������I�6�Q
�ΦZ�M�D���?�O��[��`�q��!j��h�L��O@��""~��p�����d�f�>ib�ϙ2(P�j%�5Y?<	�i8�	�E���O�"}F��Q���'�!*-:��/aW!��� w��lfHt�!�	�#��z��$�	1�t$X��l��\`Q�0(Y��e�ɛW���'������Or��OL6�H�N�ic�ӐIC6�4I�EL���\��lv��I�Z6�eJ ���,�0��:V����fп��-P�ɯ>��>	��; ���rl�_���cF�@�R�'�Tʓ�uE�����`W���4�q�Ƅ�
Q�ȩ��`��?)	� J�M����$;�(�
r#ڌ�t<pA-[�i�f�'�>�lZ5Q�����ؿ���JBǔP�|T��Gˌ�ӰiN��'��Y�����._�_��0��+֡$afI@�_}X6���K�<늙{q`B�74v�@�#�y���yRU$vz ���wM�p�����LlE��t�pǂ��y���]	b�9�Cm�*C4O�E�E�b"�5�f�5*�dt�L^6_�pd�I(�MK��iX��'1r�']��'ћv��mCd��GCN),X����y2��s�X9" +�&�M�7E��W3��l�k�Iq��	%�I{?aT.<�� �ǧ�;�P�/r�4C䉅9��rn�1&�h	�i�.&���M$n���`�����^�;���
K����'�͛_h<��'���s� 	~������-J�\�;�'X��X��>4҂Q���8�p��
�'t�(�E�OR\و�锈?a&�x
�'�����oox<��oۼ)�,Y��� �z��-QTF��ֿ]E�]��"O��S0�26�$l�q��iZ6��w"O��S��O�*X�Q��0ZD�s�"ODX $JU?5ͼmXqJ��G��p)�"O����)u8�9�*B�Ǌ`�d"Of�1�%��-dT�Q�	�&��Q "O>D�G���$F��c�_�k�L( �"O�%k$���x�p��h�
� "O��'^'����	�?���K�"O4��DM�9,}��@A\�\@e��"OFy��k�zt�(z�k	�&\��"OV�Aƅ�W���I�L�M���"O.�CqA��Q��@�π%�4Jc"Oh�c��/P����Oع'�V��#"OD�;f��h���#4_	�6��S"O�ܫV��`��Å�͞Ѩ1 v"O�yUȟ_ ~q0U+�� �Tl��"O6�Q%֬٢�QQ�F/�l �"O6�A�)��3�G@�W��i�"O�xy��)ϐY)���4O��	��"O�v�ގ&X$h��E�J �"O�`J�KHz?��q �v=L��2"O���F	�b-j����.Ζ�hg"O�� ���|L1���D hAld�"Ot��qo_�JUR���պSUP��"O.}!�� d�<�"ނVi�
"OR٪sd�=Y�����!�>8�P��"O� �T��~�J���%���33"O�h3%�7� ��/�q�
��"OR�	A���J�U�Ȣ$��AQ"O� 1��,O�MQ��T�{-��"O��h�0��I����nQ谹b"O�!�g��>
jd#�I�t��l��"O�1��J̦Gp��P�f $?�
y��"OԤq�Զ/���/&X����"O>�ї�ԓWm
A�gXT����B"OjT��P�V��,wx�s���!�����4Sv�Үyl�{J��i�!���.A&�y�)��[i�h��
Ci!��IV,B��"�8c��:�!�m*rI���K�(������C:v�!��M���b�Ś��Y� Ȁ�i�!��T4&��CD�B+b�b�(��$�!�d�7cm�ՊrݎZv�3aE=w!����n�g��o"0�O �<k!�DU7B�"e���,T2��.��w�!�Ē�h0A��C5�P5�%�W,>T!��?Y�A#b����!��Y5$�!���7i��b(���xtK�1�!򄝼eZ:�"��O�,F������+�!���O 0�E�� !jA��+
�!�Xt�IÑnTTȀű�̊(�!�ʝi��'h����+��6�!�Q�e�����ذWn��Xu�΍n�!�d��h�̉b�F�3 ^`��V�L�0�!�$]�m�R�"`�n<�a$�R,a�!��K�e�ѢW�^�HH���4�!�!K�Ʃ2�o��(H
Q�l�j�!�D��*�8	r-G=Xl��'K@$��x�(���<I�f� 8�v���D�-�0����C�	 �PAr�՚k��)�!�|�>�5&�'A(�~B�N�B�O*�� �G7)z
���Lq
r��P5@�B�ƌ(#$�� ��ə����L<�`���� 梚�[�&h:Ĉ�e�<� �Uʥ!ҙT�6Ukǎ0����""Ou��|�<ݛ1�F<^���6�'���&��-���B5���`Ka���n9D��1�E-5��榈:$VF="��:ʓ����,7���:%TB52�ޟh����7+�(�DH&0��:�"Ot�͐EﺠQ�	W�kC��Gk� ��y�.˚$�r��&�H�y�~	 ���vށ`���b�ƐQ�Ν��|B�2�O�1����?!���
+�pR�W2E.��`m� �����_ %r9k�BԂ9�;)�d�7`	�]��K����6|��s7H��i�4Q/ʓ����R	B�y"(��}l�,9!�O��M��͒�06�Ԋ3�]�,^�Q�ȕ�&�9��ϯ=�֕�R@�юX��	R(!0e�#>YH4�)LD��05A҃@W�-�i�b,�I��<pȊ�Ez�� ��U����!*�$}���ƈ�me� U T:7� Q�ׁ_���?y�A�+zȐ�%o_�g� ����E:��A��Z���:�ƈ0>�t�t��*v�f޽X�0��M6f�]=_�Yq� m
^���VT,����4���q@ހ.��Lz����m<֤���)��E���& 3����+���P��6��Db�c �i5�BK�+��˓T����Fd�����MGƽFx�I�R:����Q���!�B=���e �P���{�hI+&0������%�Z����< ���2�c�\**mZ�ꔠH�џ@�˞�H!�e@��v��'���|��y�q��3Z�r� !�q�gk���X=ۥ���s��gH�5{��5@�#6v���sF�?����C A9xi��ɐ!4P�����P�D(��!5�Q��Ԫ=���4��qc�#F�.THt^�� �B�q��I�`��T;p���F�3V� �$����R�'"�3`�Pw�X���kJlb��	a�N�H�W�I��,"�dơeۊ�X��U�!�`��d,�aKjJ�툎d�T� ��֋M��[�4��!_�0�vPB��O6�Zc�Xb���3�J��Ů�#H��Cȇ$0��H C)T	^���쎮F�VYW,B7Z�=@@bR ���J�L�O |��͑&$���B�<�ʄ�gID> �T��ƒ&p�6���O�z�F�o���H��nP3r��A�/	~%���i�O�Yx��^��T2b��"��=� .� -0mP�
O�my�!wZ4۶�� {F<A�	�1�5A�a0o�p��^�%��yAc��qT ˮ��	.��	�#��%]��T��ܭL�R����/h~�Di�'�~R��(R^H���!L�6= �ضe�y���
��E�9�D)S�	o_@)��;��EQcJ>
�(�e�H�L7J`�<�%!H�I=^@�c��<����%�*���eU�1 !V_aD��kɬ^���c'���Px��U�d,2�����,�D��LV�z�b�Qy���7$0�Y
C6�Vߟj���9��T9�c�.�iq'K]2 Y!%D�k�mZ�nDţĄ	�tE��1���1bҺi��A�=KO�TA�'~Tc��$lL̟ͫ�I}4������8h@�1B��&M���$�5Dl�,Or�S�D��[���S�aϦs�M(%�i�|\�{�2��T�5LO(x��C�2>�P�XY�d�����`��p���>-�	��i,���t䝥,r�@�6h�=��'�LyC2A�67����D�h�*�Ў��%�����I�186:x�ϒ{��c$�A�2�!�&-x0m���'yV�X'��=�!���ʰ$(���>@�!I��!���b��A�f��-q�i��n�a�!�'l�!��.L�b%�RjNBay2�C\���Z0�xro�MU8��#�P,�2ur�*�~�<������6�ͮ=e\� U�u�D�_~��@Q*���0|
���?��w��)(�~i��j�<	pn�P$A�E��z��E ��-OHL�u@��1�1O�
+�]u��uiU��2��fO�:������1�ǩ,�ʈ	�ǋ& � ��@Z|���f������ȫ%�|���]ax�D�@IF�&�D�6���Xrhb�@�l�t�����:u�RC䉨j�X�1��ʋU� XJ#��'B(��pi�d��E�D��I�U�<у�r�j]i�Dɦb�!�Dɪ	��*Ej�
 �r��a�1={����,�<�A����|�<!7&�V~���2!@�]��[\<1w��#|]�ǪC+w�*���9/q�E��V~�6�b�#cP��Ȝ�4=�m�am6,�\���IF�ȸ���hִe�'��E���_�t�ڝj�v̄�"!��.l�Lx#��2���X�K%�e0"�����5H>"~�K��6�,(���i]B�JvN'���{�"�H�a��+���&+ԏq��P�����'��X�������Y1j�@�O��T�S�c׼ �#e�-v��4�1D��Qbœ!�Ľ�t� �:U��(Gm�>iN�%8v́�e&}��� ��
�5rV�;U���'�V"O�x TgI�K��S�l�&j!�s�%,}�DYI�V���+���[�7ǂMx�f	(
�:U3��kAaR�H�Cc�����S!�P�q�Ӑ/�6�q��?�4݄�	�P�� {��Ot�^5*��ݛ+ "?Q��X�s*�+��1�	L�N�<��
�#$�8��9&!��:H�U`�B�yu�9貨�a��&����G_�S�O��i��HV*�਒�ջ*F,��
�'�Ph ��&P�-A��S90�TQ��>I�!xtD����}b� ?$A HB#Ť3�^X{����?��bƀ}O��Q��/�(CG���C�t�F+�W����D�9O�ح�2�[ZURY��N[�\�џr���mlQ�|*R����Ur��.PjLp[q�j�<Y�N�v���`�.wʠcpL�~~`@�\�E�=E�ċ��+�8��ׇ/;Ѷy{�	�4°<!!�5_t�e�N�8Z�nөe�\���Ɓ�;D(��-D�dX����A#�Iɘ7I�he���'}H��m���fo�O>s��XK�Zd �g۪"�j=��h(D��h��-_ �I�k��,5�¬�+�Ֆ'kd��l�2��Ϙ'�`zLE7k*���N�B=]Z�'�h:bI 2��M�tD҈R'�}2'oD?x��)p��YJE�}��8i2zѺ�B�/}��}b���?�0<��kV��f�k�S���d	�:�]0B-r��9�)Gu!�&Ss�<���N0���UAX�%����L�t��qK��Lj=E��9��|Sᑒ,gԌZ�I�!��]�4x`k�#/�H!�E�mv����<�seDg"���|�<�Qc�aPy�N-L),��C�_<�������`�H�-?�
���M+P��i0������V�%	EN�� �\���Ȓ�7�h���	(s�0 ��DD����'��ШS ���d��A��s�'�l(�EX���$Ӻ��M�����^'w8�a��O�Q����(�j�4L��\�8a�
�'��E`s�Q�3��QQ4d	�S4f��A�D�I�R6b����L<q�E /���s�� ��A2q+Km�<aÀ�h��iQ��a�@bAO�d�<�Q�CR�)�cł��-³��k�<aDV"��-���0O�j����i�<�1v^,
�t�>�Q#X�<q#����h%�V�+2*���Y�<yŬ�W*�E��BT� x���JO~�<iPA߄/yT\�PUX�s%9�C�ɟ7��1k�D.JPK��tC�#3<س5ژr~  ���^C�J�r|	� չLNx�r�,Дy$C��2vK��£�ה?dx��P$#�C�	�*A��)	9tt�Y�KO�(�4C�	5L�L����q2�ĨF ]�C�I3m�,(�Bl?~g֥��}ҤC䉜6z�S��Ƹ/6𔠲-�j�DB��+E#R5�k�_ݦ���.�$B�IXP�+	y��H:�k��	�NB�I�W�b�)�OM�Y�����A�4�FC��=[����U�ӥY�9��!��aXC�I#X��Y��+�6~]؀�! EHB�	�-�`�s*HKcʸf�̑t�~C��f��C`�%4Ɓ@�kٸ=�hC�I�4��R��u�� �fdjC�	y�#��l�~���e�T�^C�	�W� �G��|��$�P,N1RC�)3��z�	��|N�!s@δ$B�Ɇ%��ᑦ�{ H�0���B��"\��x�6L����7{�6B�	�)���Am�4xI�I�P��L�����h�pLH1��0;��-B�l\�3:�;��+Y.�X��� ���lъ�]�FN(�8��"O8Q� HE)1�h`᢯� W���r"O��p&
�
X�����#N>��H:�"O�-��	�������g|88�"O��I*z}����1�^p�u"OZ����M���8=o�8�"O�4ɕ@қM/hdsd!͘5~�	R�"OE�C�ěx&����Ir12C"O��ٖ�rH���պm��b"O��!diK""���t��#�y�w"O��K���ye"4�@�"�����"O��A7*� 4�z��ukS�Zi�%:3"Oؠ�',¶D
Yd��p[X""O\YӀ�4�J1c��M^���"O��%R����M�<��Q&"O���P� �(LB�'K�r2�c�"O@�ڥ$�~'؉y�*C�b� ���"O�!�e�-���a���=��]��"O�T�o+pr�4
6*��2��m�"OP��C��?Q"�bt(��B2"O"e��C��đ%��3\J�p+�"O�	��� h[t]	�5:u
�"O4i�G��b�\�q']I!��"Ov�a��\�]6j�A�c�A�0��"O�[���X�@4w֏+�����"O�ty�d���(�h��]:'���3�"Oޭ��K� ���z�.B��3�"O�y�����O�$z���P"O��"���*døa���#do6�Х"Oh��0M��X�@Ge;��$"O��I�^� �g���'$@L�A"OX�4��5@�J܊Q�C.,"VUk�"O"����������0F�"Ov��@/g���*"c�
9 �И�"O���5e}!
��dեm�C"O���G�@�����`��3h �"OL�K�Hd�J�9cmK;^U�t;�"O2�����]���(f�Y�<���`"O4�դ��ȪQ��+���a�"O��[#��R�v<z0JPl	@P�S"O���2�����1�]'�d0�"O	���b�)S祟1;�V<0&"O��F�S�R>,�E�Ծj���"O����l��,�Y�%U8ag�z "OJQ�ąT �z�pv�Y/��"Oɓ�O�`M�h�r`�+P!��"O&x��A(~�L,.xn�i���y(��tn��)o�P8�bR�zC�ɯ"W�)�a�Y�CPl屴ٻE��B�	�h6�q���<)���%K�LB�	 ��(²#�)*���8_�C�	�M��q���Ӈ�x���C�ɂ|�C7IAs�|@kÑ:U��C�	�/ޥ�����K�F�8#���,4�|�.���1tMEn�-�Xxxvǘ�L.d��1MD�̐b;���S=B�IDx�h�"j��D���e�-!3�M����O�y2��<Ce�В�mZ F�p���L8�(�s��
o�S��yrc1�^�8�=���#��=�yB�ۊ�*�0���&OleRrjݸ�yR�S	��!��R�@Z$��(ςt���Qc2��Ǚ:T�����tc�*�������Ȇȓ_�QW@B5a��!�gB
5���ȓQ���R
?2�*������S�? |������
�2Q)ӱ0��80�"Ot=�P	�3F�q!�N�,O���"O����ąH .�	�.C<�p���"OJ��b�C.Y>b��W��;&��9"OJ�@B y�C�Q�0�:�3b"O�l	aȖ�X��a�pG�X͌���"O�l0e�
�<X��Pqd� S�:<�"O�4sUK�}��'dɎodvh3�"O��#RO��J@����3�(y��"Opq�Q��& �Zz�!�%�:�+�5O�m�m����|}J?�O��oS!�ŋ3���e)YX3
Of`�3H�
؉"��	aa4k 
�	�8L�	E�'6��B�j�p]���Q�}�")���$�����@�b�4ժ��A�{�(�c�T4 ����	�S�TX�朒Ƃ|��;iM����	�>y����ԇW��tI �<b��O\�>�L|:1�]�@���!�A	�^�D���̷+�uK�t��^����
����	�7�B�ɍS��D���Ծ�� ��$Ԅ.���:&U4h���r�i~���P�����{:�!�߱��尚'�:���ʉ(*F�@CJ�
�|$��2DQ��+�-��y r�ũZ�r�	��Z;����<�&Ǩp.�ਲ਼�ʁ.���v��I�'"D���� n�nHv9{�����dC� �D�H�=@\��"��26��
BK��1@!R�ǉ�L�kve�&���uE�	��'Ϊ���o�>��yR��e�v��Z?*~6 �W�~]���LI���8�ԋ��-Hz���O�9��y�P��0�%<&�����"O�#K��YY�)�1�01@W��p2�����8�r>����k�2��5�Fh�dY8�2�r%C��9 ���!Y��|2�ç$1baZR	^������֢)fa2f�͸����Y�,��n�!`!��c�D��4d\R�p�&���~d�<��O�!#8D��0lL=2t�� ���}��3�G�1��'���C	�͓Ј_(dB�>NV��c��6�]�i�Dw���Z]�,<��.��+3����(\,U�W�*�s���p��K�Y+_��X�.8D��X���z�vay2���bt�̾%����b���q�D�]&gN˧؞�A�yR��p�vf��wu�8(歉��>)⥙9
� ��]ވȳ����"�\�yRA��>i���ぐ{;j�*�Ý��0=9%N�F�܍�*�1���VZ�'�������}RD�EZ	&z|�Iu,R�`	��S�o���Icߤ2���P
�'�%�Nȴ<7ک��EԄ)0u��'¦��F�n"&M����7I��P!hB~�O�,�0�'X
�q�S��
��'Ǻ	�q2`��QІN-K��\�r���|`�#�B%��հУ��ħ|�1O�qTĔM8܁d�V���A���'N�pP�	6(xX��̓�Z��sÏ�K��aᅊ�%{�(#���[�az��ԵLE�!�ƌ�(!J���盛�O�\3�f�O�AA�	'Q[#��W�v���	�3b�b�ح`;Ąqf\�!�!�d�F��< PM�a2�� eɀ(�f�+$���e@W'h�EKYw"|λc���
_�x��	�bܛb��Z�,Q)�L������H�)C������4�
�'�Lf`e>7M�O�'t�Ya ��`�$Q�嫈�+&R��[M�}q)O�Lہ˔�&��4�ٹjL���'�۔]8L�b��'�a|��E��`lK0&�^�pi��T:�OĠ
"}2�G��'[0-X�cɳe����P<~�ȓ����T�[YL@t�$��:"ͅȓ~�V)8��r8ʠ���\��1\
`�A��1��:W�� ] �]�ȓE��$�$��$��H���'Z�VU��a���;iä2�����;n���ȓYP����@9X���q(W#]
���aƈLK�� �(U��	�A9���ȓd���dLM>2 � �����+D��<�&���#T݅�ӆ� �y'��#�p;Ug@!y�B�I�v���!ϗv�x$bw�*���)w.�	(��"|�'��EIG��Kz\�q�R)e�f0��'�P!I��*h��g�P�V�2�c�
�`�����k��q���!x#��+�aͱ?
���	���5�0�9?��hL($L�{�¼
n�q��l�B�<q���s���5lG9 0����bd�$8���ubf>� x�Џjc������<p�(�g"O6�3 U9N�QR�-� e�	4e҃81O��I��3?�@@у%�l��۶c��{Be�m�<9̞.$s�H:u�7H��ek�ʕm�<�`��y�f=%�\�eL T÷(�g�<qE��XiaB
�'�h1�'�_�<a3�\1u���k_�F�t�K���^�<�3N�+ �%9���2�.���h�V�<1qD�����ga�'m�`d{��	h�<�� �&'��� l9=9�"`��{�<)�-���f莩\��}j�AH~�<9�˘�t�s��:v�x��HC�<�f.KT��x3kK3,ц�h��U�<1��A>A��^�26���q��ͦ����#�ا���F*A8x�ʩ�#�շsExH��	W2�y¬ޟ&�ekBG�s&�H���$Z>����	�k���P��$ H6NV
T&��d���l�ێ1+%��4m!(@"%H^t5�ȓK��X��)L�o\���BS�[?NDz�j�'^u<"~Bc�H� N�0�0+Omu6���|�<1E�f,�EP$ޏ0K;)��D1��"~�b^/b֦�ó� 0� �[�h��y"�ʐu��u��M	�5*y�gIց�y	��#}�����\�r�� b��y"B�#6R򘨃�Ͱj�z�iTm��y�I��#����`�_��%ãD���yrk�	��5�<Z,Z$@"+K
�y�]�@���

�O1������0�r�k��=!�a��AM�O8.��pK
�6�v�c�jP��yB�,i?� oȜV!рvC�"d����v�>��A����'0X�0�oJ���E�k!�ٛgOR83�*�fh�� ���]p�Z�"�!6�W=��>�iؘ>�ڰ!1@J7YjrQ�".�}X��!�b��j����U�lڠ��0^TIHV⍧"г!�!D���(��X�@��F�#|�ٸpd-�D�'t����dLy�O=`1��ҳcw ��0��wf�+
��� �gp�HsҫOsd��!��T�<��h�"5��̐����!��w�<!ªܹ6i0��֏N�+ DA�	�X�<��j�;7 P �� ,#��p�m]k�<iU��_�za"A�@�f�1��l�<	7�Νr�^Ab���%Nv�Hu�Oj�<A��c������ ��h�ÒO�<I�H��dzr�A��^z\<ȅ%�K�<!��$���F�B�I��cD+�J�<�uݎr���1 ϓ(\��k��D�<91�Ӣdt�0I�l��Y4����C�<Y��:�����d�f�;�({�<q�
�D)
�s 'ӥe�� ��o�<Q"ბ%��XBG��)g\�6�@i�<a���*r�iZQIW3:�(E�FP�<�G��|�ĄL��	���&��N�<Y4�GZ�!#��$	 6|��J�<�ÂS�{���,Sr��d��H�<��kŨ���ɫr%��x��\�<�7O��l���]C,���YZ�<�vfƇk+&��P[�MLzU�EK�<�G�1]����b!;x<(hP�K�<q %P��Z��&��[��Pn�<���?I�"�[rC�+섋��Ai�<�a�<UB������8���M�<y���j�"0lP m���B��K�<�t'�
.1��)�3t�P,��N�H�<yӆ�>1���v�[�wL�ڐOTZ�<� `a� �
�g�B��뙉-�~9"OP�B�!C��2J\�
q�Qu"OZC Aҵ&����E��U�b"O�]�E�_'(�Ҕ1�(J�5��\�S"O$)�Q-Ң%���͵W�ĩ8�"OF���U�-1:��OŶ��t1�"OT6�W!6����qN�,W�`B�H?D��)�ʆ���8���"\0�5�>D�,K���'�v
��]Cې� �:D��h�ʃ(j]�`���5sT��Po:D����X(U�֡;�M?bN��"�6D�8s�,�.�~  �n	5�.�F�.D�X+Soʐi!٪��k�T(K%-D��j��W�Y�r��D��EjV����*D�,{��N.c$
��	 x�`���)D����OƸW �1g	)}�H����$D�����Z�l� '�7A�֌�R�>D����.�8��G�v^�8�F`<D��A!���4���VFBqZ�-D�<�S� �K��΋�;;H�:b�>D�H��a�.f� ��bI�R`���G;D�$�Ȓ.M�B*B	5q������:D��ad'C ��X�Ȇ�r�j�ñ�9D��{����H�hx�RhÅI�L`��E$D��``ĉYdv��n�H�xQfC"D���1IW�i	���q��\���&�!D���p	ҲQ���<&=\���G=D�P���8��"��k�(��A�:D�H����!֜���3D��Q�ی1���2�ғg%��"1--D�4:���F���!�%rsl,��&*D�p��@?)�(��%��r,�+�+D��j�F���`E��M W ��UA+D��ka���]/� �V��?#���B�+D��#�L=�����/uX|�5)D������l�ZH�C.�F�*�A�#D�P�C���0�T豬£O������&D�h"6h�ڰ�rgLd�=�Q�#D����Aڻ]R�É)N����<D�`:Č�IȀ��l��]:��a7#<D��9��̯0�(U땬�TyD�!��-D���0Ʉq��\j�
 L2��*D��z\EC��7@[�2�&tz��ݤ�y����a�h� Z8�� �O �yB�q̑�%�źN7>���"�y��C�X�ap��y����&�
��y��T�R ېe�s��C&l˨�y���"(�B3b��8&H�Y�Fȷ�yr(7Y��e��Į6�R$�4#W�y���7� ����7:��C+�y�K[��Nq����[t��B���yR�-@/�0����ڬ�q��$�yRbX#v�.lx1�E� �݃�ƌ�y�X�,{X��ā�jG<���� �y�.�(g�ĺ@$?�n��l���yҭ��#:m����',8�9����y���u9 AW�H}p�A���y���,C)��@�jß=M�� g�ybȅb���& ����t����yr쓱\?­H Q�	��ْVC��y�F�W^Mc��
5L ����
�yr��D]@�3��|tm���U�y�Ϝ{�d����
F+.ɂ�N=�y���g���ق���8*`̢d��y
� ��p��0b2�!�ㅞ�^��i[�"OD�
�JA�6��P!���c�qs�"O8��RJ=r�"2�#�YI��@6"O|��w�A*0����C%Dќı7"OL\"��i]xt�QAL���@X"OX,"D+Řd��2%*�=8��$�"O�}7�E4p�����N�!<�\�IW"O҈�q �m�uZD�G�d`y!�"O�<��,X�n��Q��
 u@D��"O�|�e�ʪZͲ�* ���.Kd��"O��g8e4"X�D9J~�@�"O�P���D�R���V�5D�t"OP����f���
ӆE����t"Ohe��(Y�*��J@��+�<�"O��Ϛ�/���X6�!"�|c"O�	���R�[u��v$
!xq49�q"O���Q�&o��؇M�A_ <i�"O�Y�ѯ\A��3KF�sX�H)a"O
�� l�Mk�%D�"O5�PɁ�r�4i1�fZ�<
�Hv"O�!��(M6�ؼcW+�`Bp"O$!�&�>G�.|*6#�0p�HYQ"O.Ts�@2<�������f���P"O�l���8(
���A
;�@���"O6I0�$�~�"���6<��u�r"O�Z$��zh�D!�����Jܨ"Oș ��B)�������}�����"O�X�D�xv08�G�z���sU��G{�􉕿{��i�0k�`��gTH!򤄅8�05��>\`U��B!򤕙�l����=BS���u�ԢvV!�Y�k����_Z*�R!�D��P¦��C��+Q�(GB*"!�Y3�2lZ�n��+����"��!������	
g-�IR�a-!��*�L�B���'���a�\!�D�<�ˢ�ٹM������t�!�Q/��X�Q�b� 	��j,�!��[#oU�q����>�~d�����g�!�dE V2�u�#꘳RY:��哹,�!��eA���D�>P!ʨC6'̩�!�ׇH&�W��[(�0��^�!�䑗W����v+S7((�@@�e[�'w!�DF�LY:%AU;Q�ȕ��]�t!�$��gWp3d��)����+gn!�D�,(����@Stɾ<[��G�~k!�$_�d�z�A�Jԇd�p��#M�:R!�D�b����%����)Uaʰ�!�D�/%HQ��.8�V\
Łܻ !�D��B�)Y�M
-^{­q�ŝo!��X�3�D��2g~f|��a��	03!򤘒Oul�s⪇�n��<�hY?o�!�dY�Gk�Hْ�	��~ ��X��!�8(�Tl	��ɀl-�a*F�_4'c!�Z�Gè���D�+~\QG�0i�!�	[%���B��'k	X�4��E�!��!-n���-��(
ȫj��U�!�;:�M�0.͏|#~H�e.�5m�!��تd+
��#�	;>I�-�k�!�$EF����#��>b�b��\*j!�ć�rS��$�M�-�<�c"��<{W!�D�<(���+H�����O5\:!�$��H��q�s+ݴ|�V�@��ŕ'!�
U,h A�
� ɶ�I�$�'!�� ��Q@ȯWD�S�Ȝ:�p�D"O��s���AU��i6�BYF9b7"O�y�B�+6���j�V0 ��"O�,3aZ�9�
T�#������ۋ�ybڿ! R8��S�H��̱�L��yRBڊA�б9H�@:�U����y�G�-Hh���ƅ�K�����1�y��ܞ1R�Q�7FP�.�hX9���yB�q��+7���|2d{�Ǜ<�y��M?/g����HÖI&PІJ ��y"�5*mf��edw�d @�T�y2�R�O� !3��R e����C� �y��,w�F��Ǌ�V�ց	U�>�y�)�9%� h�Q�K��B���y���l➝jS��;3��p&&�y��U ��D/�c*d2�/D��ybM/q�$�4���� ß��yBA��.(~TA6k	� ]�����y��؊r���b��
�TA��C���yrF�*�� iĠ�wh���E$�y��ߒD� bl��� \3�y��?����wT�1�L�s��<�y���'Z� ��i�����Y�� ��y��8+iLK���
l�  K¯�yrlՄ"j�4C�y�컶���yb�D6b�J�1q't5ʽ��G&�y"	�-�j%�����s�RE���y�"��������9<)��#K� �y�)�	��US�e�8k(�����y�C�5��M�֧.a"����)U�yA^�-�B��n\�I�Ȝ@P��yr@�7C�9�L��I&$���Z��yBě�D�F���K�?�P�أ�]��y��*c�8GaҶ2�$e�����y����p��̺QB������yb�[+8��;5υ 
�(�P�c��yBh���x�q���3-L�I�F]�y͉�gJfش'B0-X�@X���5�y�D&+r���'"�Uڦ�p}B�	�X1<1J�(��N�~̰�Z�ws B�c���9�����$+$n�41�B�I� ���� 6Ӫ���.��RyfB�I�q�9r��Z{z�7���NB�	�3����ʂ2^������u{ B�	�E6��1.��{$�+� [�6]�C�|�Jd�bÅ}�6%hUc�#t��C�I�A���K���92�*g$Մq��C�I�Y0��FI�&ّ3���y��C�	�/��P�Y�sN4���	�2qzB�	!Jc�E	�����2�n� ��C�I�W��i""�C=J���/yE��s�"O�����\�����
?��r�"Oj�b!�A1X�����N�=�qt"O:!�޲6����띙p_ڸx�"O
�"� oI� *� B�R�`���"OV� �H�� `D�nB%�U"O^����vCj�JF��XQZP��"O�hg�/}�vh�ču��Ԋ"O��aEmF�vV�� iR�l{Z�y�"O��G�]�8�BՑ�Ra@�:�"O`����IgL��!��#RE��"O��ۓ�X>`�x�EY�lBԍS7"O\��ǩ�,e�`�j�F��I&�H�"O�(�H�*6�:��cƏ( 
=X&"O� (m��j?>�LE�U����!"O&�뱯�8���8A�Z�>�Z0x�"O�-�D�ͥG6��W��rՒ}��"O�}�Rd�H��P馨=��Q��"O�=��T�MG>�Ja�1y�.U�"O�\�aߣhpD�f�˼:�h��"O���@H\�]r4���	&ϢE�B"O�HHB)0K��X�R(U�|��19�"Ol�SU	eaE%zwD Z2e���!�$،O��:C�A.<p�Q�dc� I!�$�S�\���]�Nh��J����}1!��'8��Aj��uS �0�Q7>!�Dߑ��U2�jN9F]���@�\��!�DJ�e���"�C�F����N�[�!�Dع/G����#3���HʋP�!�dZ�kzᚰE�).H��HF+o�!�D�r5����̶f���;�-�.�!��M�PI�x+���0�p���p�!�DΛi�����T�'c`p2&��u!�䚾u� �"J�7b�x	#�߹gp!�d^&>���P'l�!>N�ĲdĲ"4!��s��;���%_�fLKң,S!�DB>��H��R;H#<��"�H�!�dN�G�A�@�f�& �"�F�!�$�f����X/	�2@{�Hƈx�!��;�m#f�m�pٰ-��C��*;z��EbH�`!��$4%&B����a1��~`���HB�	)}�����C�XÄ����+�C�	A��,Z��\��)�.J��C�I�H0�D���\�RQ��� L�C�ɞV	z����D�/�0a���C�I<a��m3rU�|j܀A&& rC䉎#�sī0�]{5-x�HC�	�X*� �"�B2x4�Ȃ��u,C�.R�.U�T� v|�,� 8�!��Ŏ7����v�t���b�!��(<N���L�3a�Y���&9`!�Ί4�5%m�MT���E�D�sT!��%Q���G
�H��pK6�M�|k!�T�m�p�d���QaqC�푳~b!�$SW��ـ�ʚ"C�x+�Z73:!�$S
j2&M�K��K�fxyǉP& !�!J����H�8R���(U&	!�D�)b� ���s�����h�!�d�*[�:x1�FUo�z8��O�;w.!�ƾ1"�Q��H�>3�6���M�5&!���'(X(��=$G6@
͋�!򤏋�\� �`ʢwV���i!��,K~���ѥ� Cb������y�!�4}�Ly�A�^5(�\�	�'^�^!�B	I+
���m�;��瘡�!��4K@$Ɨ5,����E\�F�!�,g1�\��nD�Y[�mJ�%ӧ^�!��&�z�ٗkױIx�P�JãN�!�d# ʸ�r�j÷);����)!�!�$�:18Pp���.u) ���^�!��� NJx�hB�
R��d!�Z�!򤞤�B!CJ���!�/N�_|!�D_�x#�H2S�gY�N��6g!�Dڬ"v�|�B��gQ^ S�O+Sb!򤄥D�2��!JEnOX�� m�Z3a~�U��su�@����/K:V��U�$D�h�b�����Ɏ$�>�ӥ�"D�� �h�A���L �熀+`�ڹ��"O�A(2�\��޴딦��E�T�"Oj��կ�'W<
���f=R�nC�"O!�s!�p��A(hpl:Ap"Oh1�!N����:�0���"O���II�I����E�	/b�~���"OZ�d	Ν �t�%�Μ5��Xa"O�$� "�[����@)����xU"O��0V�Q-*E�yX5�B��lp4"O��[t��xv�35)=����"On��O��J��X��i�nل�z�"O���U�x��z�F�����x�"O6�2�_>Ͼ����8?�ƍ�A"O%ҤB�4|�D,+��ؕ@����"O$�zI�Ǣ��eZ2@r��"Obm��QX�D�"���1��ڃ"O�qGD�k7�59Ӏ�(gĬY�U"O�lBFAja�����l��	R$"O��ISl�4�~���B$t��m[S"O�} KY�&[�h��F��,�A�d"O��2�����1f�(�~���"O6`r!S�|�6��0E�eAl�3"O�\r���X�ޭ92c���P(c"Of=�b�$�tXr���sy�5�A"O �0��ԋ���á!Hud�X�p"O��-ՏM�|RT�Ə��ణ"O���"P	0��,��tH�"O���)�9r��$�dL 7'�Sa"O����"2Y|Z�"b��<T�J`P"O բEh�8xH+���%{�!��"O�a{7�+CX�Ԩ���gm�qy"O���4,
�sR�A�n� 'e�t '"OJ�!��Z�b��,2J�MKw"O�Ĩ��Z�N���E�pB���"O�]��aY��Q�ʊ�H)�Xx�"O��8�흊{�L`j`�E�xq��e"Oh��%0��-*��Ø;��K�"O�Qj�F	rt�:%J�aՖ\��"OzE�P�v�JD2��S��L)� "OX�z�!W<pf����,V2���"O� +���I�@�@<XbHH�"O>B�� �$&Z���B	e���i"Oz����҂&ۼ0jա�.�Ȝ"O���r�I�*�x�!�f�Ё�"O��Z��Y5���e�O,$A�4@�"O�Px3�G�a��r��
#�͠"O�9�#��pb��#�O-6�xy*4"ON�s��R�z� p��/U���!"O��s%I'!��8��u���O!�d������0*�>�Q���.�VB�0r�iK�ƕt�r���6K�B�	h��$rӠ��<	�DH�(k�C�I5>|�:�Ɩ+P�ՓgDݝ{�C�	���huA(^)A$Û�(��C䉗<�b��D����2Ԛ��-h�jC�U�A��� ڴQ���eLJC�)v;��b���r6A2��
S*�B�I���ݩa��(JK�9���F�j�B�ɣ t8�QD�{�hdrċ_*5�RB䉕a���Փ�J��� 6�dB�	z%�	Y��G�(	Re0�B� ˆB�	�'�\�H�)>H�P�^�mԜB�Q (�гe�:~6�q�ū܇>��B�I�8�:f̈́8PLY���jC�)� ���&���
�jL�,�2C�H��"O�$��P�p06xo��z�.�2�6D�2�ڑJ�8�9P+O0<�5���3D�D;� Aq�A�c�	4nĘu�v�/D��j�ܢd��Qg��>� ñ�9D��+ġD)	�܈�Ҋ�>[0�t8-D���5�$e�J�,�>h�8���+D����˭Y��33�[ }3F-�6
)D���r�σ8�p��Bg ~5�U�,D�<�3b�"d]RHR�eާ4%0��CD&D�$���v=�#��]<Q�"�n.D�̑�
#O��[a'y���B�ɴ|��(��ǉ���XɄ��;�B�	�P�:)ANK�Q�ٲ_0�C䉍D��YE�+7gBT�V)� r,8B�%~��Yk'����1���2��C�I*9z�Z4�|x�L+���~�C�	�|yt��t��n9��tdB<	�C�f(�Q�\�l~0�'�^�<URC�ɴ?�l3�N�be$9A�Ŝ�B���,�I��L!�^;2Q[v��my.C��F���N�({J9�q�_
0����=ʓ]
D�5�֒0�r4�A�0F_���ēQ����qh�9��Q�Q�u��Ą�I�t&���bC[̢mjp
�(}JpB�"L�j��QH��1�DtJ�HۊK4*C�I*"�ʰ�@��� ֵ��٫�C䉺^,V���Z�1��7��W��B�	*��[f��`�ip�.�4SC�		fxE��JL�K�0t����Z��B�It�l�B� w���"��4K�C䉄.08f�
����p H�%�C�	;b�������G�fztb�O��C��<']��1��$b�V$g�#o�B�	�E� �NL=P� �Q ��!�JB�I�D]�e��
4��l��i�<B�ɹ9�@�`3
��(z�}�ୁ���C��Gs@��l@�m� ��M�B�	�:�I�C������e�I�"�C��p���q��rN�4#��C�!u�N ����m���k��C��*���s��Yxe[�9v4B�I5j;�X+�kU� 	Pٻ�6��B�Ɏ>ڝ�"�E�v�F� P�!��B䉑S�MS��?�j���Ȥ@ˢB䉚<���3�A�l�N�)�LƧU�B�	={�4��nɪc2�#�جD�C�ɋ�̀r��+��S��4X��C�	=�Zu�`�ۛ�>�IճY�C䉏o�h�f.X,�D�&���|WB�	H�ʤ!�z��p�E%W`�C�	*"�d�
6cS+��0�� �y��C�	�bfq@0B�?h�qtB@=�C�	�3�@��IQ8.�
Qش�^iB�C�It~^�C�D/�A��\���C�I�Aغ��dLyἬ;�k�:@��C�I<!I��R�K�@"dh[�@��-~�B�I[S̔
T��z,@c�JJ�:2zB�I/�j���#ۚb����H�8�dB��:��%o�7׸�;3&H9PBB�	8�t�#�$Ͳ��(jfL$*~B�I�=m�%Y��Ԥ����C�nB��9{�2�	�. ��E�׍�0r�DB�	%/�LuS�"��ު�Q��C.J�`C�)� ��٦!^ ��䚁Oƈ�"OF������}n�X� H�Ӆ"O� �Ls� �����&(�%K�"O��	u�ѱ���"�/D.� �q�"O���$#�!I Qٶ�ՙtx$��"O��i�ρ6Q���9�At0i;�'<&)�H�
V��������P{	�'� Ej���x�ƽ{��;eޒ!	�'�j sJU3xdD����W�$<�
�'�m���y����w��,��0J�'
��2�ؑJ�x�Jf��N�� 
�'z��g��BP�D�ωE�xq	�'4E��ƾa����lT�[�� 	�'&PH�Q���CN�4Cv ����j�'����`��6Z؉�mv��� 
�' b���3)����H7`;��0�'�4 )2�^?���ȲQ���z�'�0@�U%��8��j��L> ,�
�'�d��L�F�3ք]�I�X���'��Q%�GB�a�6oɅB�,E��'!����,�h�R4���D�?���	�'�����ϥCv|���3Z�E�	�'�j �"Q(|g��R�eL�܍:	�'���2R���+x����7�N��	�'S�c�N(P �i�$��kϦ��	�'��(��ߋL��	�� �pB�$�'����E�?E�Yj��5n�6 ��'͊4JB�H!Q���Mɩ\U�0Y�'	��9@�?��0сhN_�nXb�'R�U�2�Ȗ��h��!T�yR�'�� ��B���qPL��mV��'Q��2��nu�x� $=e�R���'���P�,���AP���mBl]��'���8Ĉ���.X����^��	q�'M�����V��p0��!	�Q��R	�'	8�u"�	;�` �ʌ�&m��'|����0̶�аJ�!h@v1��'���!ӰS�=�P��Zp�D2�'Qܙ  P�l���R�
S�@}�'.��HV� [��R��T��aZ	�'W�a���P	Sv�UK�m�KbPE��'�> PW�)d�Z����@�^-��'�XC3 �3by)r�N6� �)�'���@�#O��}ӆ�W)?+���'LT� ���H�%{H��3��mq�'<��%O�&;�<}Su (.=�(j�'(A�Sn�Eh�`$��*$��d�'Ͷ�1F�@�v8	��g�rJ:��'Qڕ:��z9�,�����lx��'%Ձs@�+8���h�J�o:����'�|H��>��X��_�1�6љ�'1��8��U�d�P�PE%ӳ+(x$�'�ڡ9�E,-�J��*�+t��H�'H|�\"�Q#WN�;>j5�v�U�<�D���F���S�I[�h����HKM�<���� DX��O�6��0�_J�<a'��L0r�K�i_�uI�CdOGE�<�Vh�ZD�xr���2���Dh�<yE�5Qk=�wK��TsZ$�a�p�<�t�T9�X��"��Qr���Mu�<1�%3w���U�4A�I���y�<���I40G@@8�E�(3O<݉�"�t�<y���$@;N�����9.$ّ�F�o�<��+�9Gr�"�I­+���1�l�<� NDb�k5D����fr�T#�"O(�Чƹl��-�#��:*�`�8f"Ofͻǧ�&�6H�6���
K�(�"Oj@$�b�|�&@�/0D�a�f"Onh�5��[.�!��,EB���1"O`�2�kA�F��A�A��&W%dy�6"O�ؐ� 43 l�U^7B�I"OluY��F12�p`T,\3X�.�&"O@8��aZ�Br�ay���c�P�S"O�}۠$X��`rFh�#O�2E�"O�I��S�F���7�$4�ʭrW"Oj���kREN�1y���$xb3"OЈ�\�N�r9��A��P��Q�"O|����W�r��pp#��40Q"O��7� %*	Dd���H�+����"Ot�J҃Z�P��`��RQhz"OFԚ�Gסr�kY <�xU"O�ѻ���6*����K�'?�M8�"O^D��B�Af�}KA�S�^ �|�u"O��aN�k���ɑ�˦+�ꉹ�"O U2d�-�:!aa�9y �H�"Obġs(��"�H�
'���"O�r���Ĕ�7Ȇ�4�~a@'"OX��%.�mz�q�L���0�"O����[�oy �2 ��]�T�"O�}D��W�t�D/�
��$��"O�QE�%6wBiY�B����"O����mRO^�i�jF�s��y�"O�b�!,=!v�)�
��Š��"ORyV'��u���Y�m��	��"OF���&@�
���=1:�I0�"OXa�j�94���X�-99!ʕq"Oj���kӈM<�� T�xk���"OI�c�(2�>�J�L��/W ��"O��a ��y���ْkI8BLS"O�Y�a�Q0�d8��ʁ�H�4�!P"O�}��D���-c���aʄm�"O�I�4a�H�N\��K#*��iIQ"OB��u�ME`���fֽV��8"O>��d��_�J�ze��K�(���*OZ�nA��y{��E�3n�)��' 	�@� $t��kI6�n��'�LeH���4<�h�!R�Z�4<V-�'_��`����J���;�$O�0��=�	�'ޜz���+���L��8�ޑ��'"�Z�cW7Ic�Y��"Z�5v���
�'tE��%чcbq��ǈ@.j4k
�'1�1ӂJ�O�����:-���
�':>5#$hȿ5��c��L�:����'*����g[�7?�)��$�=]��4��'��� �S;<���a���Y�d�'ꚵ�1�1L�^ ���W�S�T�x	�'=:��U�#=�|R�m�/=�@%!
�'�^ݢ�#��"�E	�e[96Xz	�'�D�bE7 �@B�Ò|*��+	�'5�\Soo�*�Ӳ-��u��p��'׌�`�hG�ё�]%x �'dq��ٹ9Ҏ<��c].�\��	�'�.��T:}���2,��nX�P	�'�<�* ��Z���㉛^a��'B`<��L��L�H �P��� ��'Z�H a(ۺI�@�0	U3Ő�'�0�)!kR �L�Ԭڏf��'$'�V��-�G�7��̨��� �d�P�V�Cu
�ä�9r�M�"O3��ٶ��ɋ����U�*5�"O���p�ܪ3�N	� � "�6�g"Of]�S�X�b`�i��_?BD��� "O����\X�� ���%v�:a���'a��|��lf��Hm�x!����-Y�y��.e�t����;�T�%�O&�y�a���fH�/̅���	5�y��4�������, ��ٙ��*�y����jhO��꨻�i��y�߸m�B � FҖy���IQl�-�y· �z݃VTqx0�9�̓��y2�Ef-����#;�4�b�*F��0>aN>��a�3?��q¯T�q��<����e�<A�J�JrD�;g��h�T��|C�	p�84ocG~�����[� C�	FR�ICf&J�UFPaH1h)~��B�	
*�!�Cj��\� J(|�jB�!r< L�DF]�{j���C@��x C���BEy��<YF�%�%�����2�D!h�0��S۔ı�׀}��&���?v�L�f�XЋ��6#�@ۇ���<)C!�?�p �&��~�V��D�R�<�#a�(�����N<*н�!K�<���B �u�[�2>F)��`@D�<Y���P�Թ��T�p.��#���<9�$`�|1!w� 02��6��`��P��N�I] \� ��Ւz%ā�6��:��"<A(O�Ov�>�b w��2���x ""(���ȓ�F�j��Θz���`ܙ-����ȓA��
��I%*� fo��$6=��G$H�
���pevD�0�L��a�ȓ0��P�1��y�4����ܠ'�����Irbh"k� yP$����_8���	yy�I��E�A�dA��<��	�=��O\�:EE׫\\�x�Jl%�H�#(�P�<i���52���3%ڜ#�H!�\F�<֦Wda��aV�L"	B��{�<	�k��;�(Ȋbe����96.m̓�hO�����a���g�Ӝ|Ƽ���a5D�p1��-\�`5h�j�x��TY`'3D���-��_[P���e����DP1D��i"Y�NZ�\:���.�<r��/D���
dU�Hz*�4#��� �,D���eeR*	P�5"bh�~�c��/D���7�IY�:���5ߪ��B�8D����\k���Ҁ_����s��7D���D�W�U�:u��Ie����4D�p@����W9�k��rQ��⤅3D���!��;:X1v�����/r����I0M�qTfB�CK�����$�B�ɦ^��U�����B�T�[�-��F��B�I	A�PeQ�)6}���A�F�H�p��d?��/J�pA�%.�	-ޞ��DJ��@C�ɫHD���uHZ�>��@ϙw�nB䉑y�r��w!����9�V2c&���en���!�.dǦm[�n\-jh���?!�u_�YrtƝ�"�0�Ue�9@@�� �p�A���x�yq!-�W� P�ȓ/�.;��� +�6� �g�`��ȓ_g�@(`F�0&]8!阈=g,��ȓPVt͐��"74�A�L��_4����?)'�6YF07�?o$�p��Qt�<���!��i�ЇãP���mGF~�ާ� ��d��+y�
p��G�9rZ�<��"Or��Ǫn�B�0�Ƈ�P��I"O�5��+>~�ٷ")n*D à"O���N��O���˄�
�"O��NЩ5��$`�  :aR���'E��'dlQAf ��D3�M�+��x��'�J���
�Q�H@k�R�s��ar�'>* ��LlH
����ײWŊ���'X0yR��7�|	{����!H	�'��@��GC�	 |̐Q�eϤGHB�i�ē�`��41Ή��6$�Dd$D�8�A�]'�!�Qa͢:F8)vb6D�x�$�0��	�� UTxX��7D������\���j�#�z�8p�E�u�G{���G�6	�r@�C.C��� �'�`�!�dR�2>��a�*8	")��f��!��J<	���=�,��gT4z�!���6r����jא&�TI$h��YlB�I�C�H�'B�K�̱UgL� r�Ɠc�,,�`� oϮ�ц
X�xײфȓi|nX��'�7i�lٔnD,Ӣ)�ȓm���1�_9Kj09�L�?Ē4��M�`,��g#x�0T��U�d��ȓ��Є��;:|f���\&�����?QW�6�8YI2�W�"@��c��K�<A
��;���y��@�d<,D��� d��<����>Q`΂�U-�	h���j��`"}�<YD���YTXp���������oXz�<�b��G�(����i����<���U��`ݨQ)L�B�Z̀�	 A�<IW��9���a��K��ph�- g�<i�\�b����gǞ�vl2�B�)�d�<a���(6x��Ok	�H�M	w�tE{2b_.QNăS$^�+�ac�b��y���P�K�C܎�a�\	�y2��'�������4�L�2���y�.�fC�m�̈`V� i��	�yBJ�?KU��(dOá`՚�Fݪ�y��-P4�ys���/k���2��/�y�GN�?�� iP,�/u���gf�;�y��b�����,%5����.���O*�=�OI�(�Wc݀ ��a�1$]�0,��'* �3�,	atF8��V�T��`��'&i�Dn�O�(�(&?�����'qH�������JԊ4�4@�'pR�id�H�e���;B82�h$����D[w�"�api�N�T�ٷF���F��]�0q(�B�ݦ�t�zF��y�/C9>*(��L�0TT���5���y��2j��A�W]e�1P�%�4�yB�U�r��]��'�N��1$GG2�y2��(�R%���E�7|4��3%���y�,����z�$FOpx0���0>yN>�$�|ؖXK ���7���s�OVp�<����&1����&+d�"=��KKl�<r�WVD�óK��~A�I�f�<���5zÒ\��� /�|���^�<��I_�&����ޗ[�(�cΝX�<	�h'=ۈ=��&ϖ	�0����W�<���'zx�\`�A�3{h8U�S�<�����iVjx��`\�� �AU�S�<q�T0Y�]h!�8*���
���M�<@�ck>�B0e��6�Eb5E�'�ў�/�������	�(!S��;C���S�? ��X�J��c������:���A"OJ�*���1F��=��mY�@��zb"O�u`�oɲl�N����� ���;�"O|@��#0=|@CF���X2H�
�"O|��&n��� d�M z�^je!�G�7*�����A��8�ƈ`��wy�|��	;P�6���F�k�%��$9N!�$����'&�Z�d�ӣ�4�!�䈈p�x��7镭jo�����!4!�D�,l�-�AG��[ZBP��|0�I]x�\xj�G���8 ƋGH4�HV@0D��P�xaw��<�͊�Â��C�I�8a��9r�  ����� 7�HB�	;O���"LR���Q�t�\B��� ��H�mG�c-DҠ7D�܀��ԒqHc��X���Am)?!���$P��S�e�N*��;���ьB䉵'��tS#s��B2���j &3D�t �K˓Z��#�m�d��@��.D�4!KŜ?V�Tc��	3s��r�,"D�$��o�x�����B/S��Qu�>D�����+7 �r =�dݡ�2D�xr�eY��y�g�I��Z铥�"?ъ�4�f�ı<�E��$ ve�L����qM�j�<qG/�M�D�����5m��#�dTB�<��FX����"e�-�vDi��z��$�̠�@�d	��R������/)D�P0�� 1����W�~6�3�-&D� �f�|��9�'�S|���A#&D�ۅ���
^����Ğ������`����ʓ=��)�	r��Z�h˔"M舆�t@qT��	!^�jPE�ir���/t��QCG�8!�:���)\�����P�'gF��Ђ�1�~ �v,�(XS4A��'�h�r`��.Ų�1�xC�!�'>������nt*���FB"!��H�'������J�0��.�01�'�T��d�&�R!#	�<:���'����틴���WH��1����'iF��ȑ9
ā�/Ґ K�i*ӓ��'D��I��T����J���A�'��[�i�1S�B b�{���'�~$ҥ'�0B�dU{�O1kz���'��0B�gY��	���&r�	�'������4"XD5��F5l�>�:	�'\ܽR��	
-\��S��8~�xK�'Lm��#�$�|����A�#^���'I8�)`cTC����k�9!p ���'�h!�ˎY������\��'�F|��/J[P�(ч��;�Lu��'`��ej��\��-դFm��*�'4�,A�[!N�ne�$T�q
��S�'dn<*�F�I|y��Y03� �q�'��(�0CȫK���!�m\6c���'1��0F*O�2�[R.�25	�<��'���� R������.�[���'�(��G�6, -�4g1e���q�'��uj�8/��`s��7Hb�(@
�'d����^%Cު-Jr�1s>`%�	�'&֑�Qn�	K����cžl�(���'(8�C�JCL�� ��3d�)�'ݞ��B�����*��*2ā2�y��ؗZ{�)�@IӸ%s����y��֊F{H�� ��v�N9c棅�y
� R�c��4殉�Ӎ3�ʨ�4"Oؔz�\�x�Ԙ��l�W���"OR]�f����id�&o�:�U"Oz�&ʇ��Lr��� �{R"O*-#�R-}nA�f*X��"��Q"Ou���Q�z�&�0TO-nxI{s"O����[1-X�cU�}�"O0[�� �t�Px� �be�U"O�d��#�5ꂉ2�O/c|�I斟X�	J��D��L^�.��aqsa�qg�X:��)D�����-6��WO�!Q�:����&D��E\�(�&�	�JN��G��Bh<9U�A	 ��)�	�e7`����Wv�<9�� 5b,m9�߈y���gs�<�a� x���e�"t3 fo�<��E����� jъgl�k�@��<9����>!th9��E�e�Ǆ�jsa�S�<$+|JNE�D@���q�CV<I��/���d ՙG�dQ�E�5%����A&B�1���\̪#2���,Y��C� �'�b�B5b�)�l��H�ȓG�*����~$a�C�O���%�<�
ߓR�F(K!݇Sx�*$Ʉ"��)���?qd&��`�PY��#�+)D�+D��p�<��޾"���Q���Tl��+Fc�G�<�3@�7FK�N\�9�.��#�O���x��+��e+c�]���F(��y�@'2�uh�a�$>[�!���%�y���d����@"7��C�������!�On�j ��8+`�׺'v�0b�"OxU
�i�m4Tp��D�8��8�$"O\�AD
L�����)>��<�g"Of�P���\S� �!lsƍZ"O@5���8͞����J�=�&�"O�PY���<6���d�[5����y¬Q���C��J%;ul Θ'��{2���O�����Y"d ��d�A�yb"��%e���Q9@Ȕ��.�y��� 8�)�ˋG�ru���
�y⮛�c0�]ҕŚR!���LҮ�y��N
����ȋH_(��DӍ�y��L!��ke
��-��`j�y"�4)��؁%�ô,TE�RJU��y�PQ2AJ�D����H6)2z�k�'�� FB�.Y�q�U$_?p�X�'*� �ԝR�t���+�7�Ρ;�'���9F�V���z�ǘax��':~UZ�`�7"�Xj6g ���P�'/F�#C��3�ʝ!k_�-�x��
�'��aC�ƯID�!ҡ뒢$t��
�'d8lj" =薹@�DY�F���	�'��H�S�˹'�5�/Ʋ( D:	�'��Y�Ď(��m0+%[�d	��'�8 �h8ڽ�ML�W���
�';�5HT�������-ҬUJ��Z�'Xlp��V�de[��SrQi�'�P1xcO�eD`RD�D���)�'��@��OY�T� �P�KVh��'7~(�F��6u,nm���G�F�v�A
�'���Y�Fح9Z�P����"-���r
�'pJb�GSf�����(��0�'�1QaFʐg���B����TB*$��'̹���+{ ���#�9�Z�9
�'Ю�{b�N_$�a��W;6!l����"<O� ����V�~��P�s(K�/O���"O��)ّf F!"���/:7b�ɰ"OE��k�$Ep��1�ɀ�:)t]�6"O2�:7P:^�>`i�ꅔF¨�w"O�D��B�9����A'��eY�"OB�r���T��[��3Ey�L��"OV�a�B&�3�}W���"O�)���,4TE! .0X+P"Of\ �_�Ez@Zu���A�X��"O����� �w�F�Õ��f�R�"O��8!/<!�N&Dx2��f��*|OP��ЀZ�ccL!�fY�@̤h��"OĘӵ��;_�Ik�ϕ�SSf1!�"O,R��ߧf�<��a.˚E���1"O:�s��H�(���+4�R6O+2E�"O , &Ӂ7]-��FCA5$(�"O���&k�-ig��`DX�E0��k�"O`5���ێZ�B�����_��L�v"O6!�e�p��"Ũ�V|U"O2ɀbo^.Q�*��"X60�A�"O�A2�`�(᪔#�C�1(!\�K�"OHU	���*
��Ӓ� i��w"O�툠��b��|� 2L��"O�u�ҁ��~�% �7c��#"O
�"#�Z�����jB��4"O�!S�~0pM��!� -_>�Q�"O��
�y������"�t`�"O(���ĺ�����&L\L9a��D{��	�m��'��?<��I��S�bD!�;v�j�Ϗ	M�*�3� �!��װOl,��%������e��f!�$-u���Ef])��%#��=]!�D�4W���q�Y�-Y<�I�'J�~�!򤈍Z��@��#?�� �gp!�ųvl�(�"�2)-J��1�5@���֟X�?E�A�3?�,$;�����N�y�L��x���� �U�
�J�'h�y��	#��I���)nzf�
'E��y"�L�`$K��*g �L������y�%ӽ1��ES�Q�h�8�����y�-1H��W�3��8Q�E��y���h��x�3(yZ�C�Ž�y��)�'Z<���h�����DBĢ$����&Ӣ4����D]^x�1NO�|��ȓ��	@k�G�T�#@�"y�$���qK~�y�NH�#F��#h�a�<�ȓF<���VAƁ!Tʝ�)M�W#��f\Գ+�9����Q�FH��?茘��_S�Hc�ϒ	�A��$���ʄ B',���2kˌ]��ȓ#����ҎC�up((P�hN� �ȓlB8lI�e��dHش-�| v���+��`��`C�5���bJ
+K
M�ȓ��H���q��a��樀��p�6��3'I-k���� 7	�JI��'W�m3�m��WX�+����@��'�ў"|b2B�	�h3І9J7R�K�,p�<��瘏D��C��/��cp�j�<��)�,�l(�s)N&5Hl��"�c�<����f#�91�A&L7���*�K�<I&�؏P��\y�
D"A�>�:&�G�<)%
N5�u��b��j�*E��a�D�<a1"Bn �@(ƐD8 �#0/Fy̓�hO1� 1B�*� ��@ap�^,?� A	S"O� 0u�֢�|x��
���^�p�*�"Od ` �8j<� 	�Y���"O���eV22�2�P���~��H� "O�� *�zřVcı�
��F"O�8R��>B� A���?�Ry��"O����)��P�0��?>��q����D{��	��EO�|��S4 ɧ�.1!���@d���ő�]��bň )!�ĺD*�MSD�^�X�r�L�O#!򄌃{�X"B�
�"�����b!�D� mw�lx+�=qÌ�Bfʁ�L!�ߙ���s.�>E��D��H���!��6.�Z�(�%��-�&MҶL�1O�=�|��&ۅ>M��Z�Yb�h Yz�<���Gk��"�[�%Ⱝ\�!��ߩk�%�AO%�Q�fZ3!�TY��u�Q-��H��_$a!��q<<�B��4�,HP�	�!�
�M<,"��	5x��[��ȍFR!�D��(��)�`�U����t`�/63��F{ʟh�(s��$�)��oX�=L�-�"O�9F-�+I����R�".>���"O�з監��AB�M3	n$�s"O,�A� S�F<j	�Ү��Wc��;O����S�O��Yp�LF�mҖO)z4�@�'�pPc��I���B�/xl�!�'n֜��fQ(P�^9j�?z�~y��')@��W�ǹVe�򊕼l�l� �'������=Z}*pE�f��'�	ѫ@�jw$��g��W��<��'O.��)۲T�p�x�`B�^�J���'�^�pW��l���0�
P���'�,u2Bp-J]bvፐ>��'��t8lӦj�h*���hd���<�'_�X�8�BR�f�Z$R5�>����ȓ`^ٻ��W�xRuYEM8v<0E��F5<�'K�X8�\a�G�ID�ȓ)�r)�d�
4Q���EC�?��5��=L��w���9~iS&aϭi����(���
bd��<Ʈ��L$P�\��T>0�iwÑ-�,3w  l\tȇ��l�'8ΕX�L�=f�UAf!�#[�h�',tS0��*<4PZ`��wP	�'�q`�<u��	�JQ�}�)��'�\%r�d�$u����8
w��3�']lh�Wm˳l��'�7�*��'��@�6ĈLO�)��ף^�s�'� y�"e�
��p��I_�li,�[���'J�Ĵ�2�L�6�y���6�!�;)�bYڀj�
J�`m!K�&st!�dS�,C���c �%J��!q���C�!��թ&�DĻ�
��*�*�fd( I!�dN�i�������%U�85!�$Y,J(-�sa�:�Vu�e�
!��6q�Xf��N�I� ؄Qa|�|�*=cz(p��O<(:� ��S��y�h�1��b2�%k�����0>�K>�DD\�Xء!�Y���9�Et�<qq�� c�\�po�r�����f�<A�A'(�	C�*Ug�} m�x�<���*UF�1RAZ�VpZ�8� �[�<�f�T1:8� �͟�aZg+IV�D&����!Vʙ�g
1r�,�u&D���*��
�n� ��7@���#֟T&��E{ʟ� �tHs㟽r��i���=	���"��P�O�)C6Ō>p��jC&˾Qk�*�'�&`��Èlk�@38:(Ҙ{�'��Ж�_�>�QqM�8�(���'e@M�V� 7_�=��1�D�B�'�p�!!D�41����l��+[�+�'��ܡ3�X��ea�j;�B}s�'>ў�F{���X���Ug��_���r�%
`�ў"~ΓP1ZQpmY�-�ʨb7) �RT��ȓ$�j�RCәkk(qB$�A7�֡��R�1�t�4zϦ����Q�V���eZ��������CF�S��@��,\`Y��uo�AH0>�ȓP��葅�@�s��H�P�,�GxB�IeyR	�C�N9"����B9Y�o\=�yB�'e�O?�2U#��l��(�£J�(1�8D�x�C�3~�)���@��
����2D���b�|`��V�ߏL-���%1D��s#�M��6)�B��d-D��t	/�~��@	�L�P)y4e)D���?M�t�H�g�
��`P�*D�\�Uߒo���0�S(/��B��'?��ᓽn���$O�c}�]Pp�J}u�C� `/��*�I�;S��	�(Ǔ�xC�	(9�����z���I�B��B��.[ʤTK�Tp���D�zX~B�	3YS�P'L�9��kG�~vB�I�P�Zm	�A�C}���b���<��C�I/\�8� [7J5�Q� �5q#<9��$�OB��g�
X����Q�Z�n��G>O���d� :݊x���
*Ș`��D �!򄟦V><I�L���Tp�F��t�!�ċ�*���t�N�`~�8%�	h�!�ԠT6�%r����b��ha!>�!򤖵82�juk�[d����c��f�az2�Ċ�s�����(�@�4��9Fx��'�d�"Q�Y���1��Cɞ^a���
�'`��3ǃ�!^�+�<��b�)D��sd��;~.�{ᯑ,��cs*5D����P�x�[�d��d�23�4D�T���[�n�C�M���h��1D��x�b�&Xv��`���;�z�� �#?y��$)�䞛r���Ԫ��!R�(yw��4*�!�dE`��i���Ⱦ`2tI��ˆ���=E��'�\���(����`��;O��H�'�(��Pk2�J�&�J��H	�'R�li����S��yia�ќ@`nB
�'i��ӱ��^y�����D��-c	�'WF�RQl�t��&L�~��� �'b>���׽c����Ҁt*�
�y"�)��Sp<�ƃG; ���ڕFn�NC�I].n|aE���\�(�Ѣz�:C�1[�OD�2ڳ��0D. C�	П��&R>-��ɸ��\X�`9iC//D��Iv��D,(�/������.(��|���O�PzBиf�AR��P�g,X 	�'`��%A��\h0�A�5�u�㓿?I.O�1C!K�i`k����k�1�"O>}�@(�m�pA1�]'Rߎu"�"O|X��Ʉ3G�lX�n�˒��"Op ���Ө`��  g-�;1�6l#$4O���v9�zC/ 
r�|��fO�Q!�dP{#2����	�	:6#�3!���>��k�@W����lτu��H�'��� ��ᶂ�� |�J�_,u���q"O��� �b��IP5�vaC�"OԄ0���S���go�k:A��"O�\r喭�aCeO]<c6NM�ů�OL���,@<�P���H+Z�`�0�#�>V��&�S�Oj����b���7eZ=�vu��'$�8i��R��0ڶC�-H�y��$)��7���(�6E��%!Nj~�BF���)6\C�I7����TeM.Mdl����g�8C䉒#D�EaƁ�7zB�٫D.�0!��B�;(y��w�H!�`� ��U�B��Kw���.�!!:Yi2��a/���Qx�`$�(���5�ɸi.j֐Ct
=D�$�S(�B��S���>���!"8?����4E��ɛ o1�� �g _'�@C䉛��N�N$f�ؤ�� (�}�6A2D��J�@�3P���((Jd\aC�x�<1P���|�)�hׯq�2Y�Ԉv�<1!�[�S�����^�pˢ����	��?��zwV�@ �QF`bV��!�H�'%�}�Z�+�=�f�зZڈ!����y�֯"|Q� fΔL蕂����y��K�DR$��5_�A2�c���yr�s�Z��C
�ڭX�G�y2&��"�,�B�`�)~9l�����x��'f4l2V��	� �A#T��ț�']l�b�M�V�ҘH�n\�Fr�ؐ�'��O��r��?qn�;X���`�)&���[��Vz�'	�y��-%�䅠��ե]��5R� Ҳ�y�N>6e:�R��SW,�񪂨�y�/�B������Е&� �i" ��y)�2a~S���4�L��"+��y�a΍B�d��M�3*)�EZw���y���@�Z���!B�����,�%�0?�,O �����x�H�8��P.A�D�5"Oh=#dD�y1��P��I�f��̑�"O<�v��1�Bq+��Z���@��"O��q��5fD��P؜&�T��"O*� ��*�)m��hH�z�!�Du��9�bЉ.Ж������g�!���k� ,���RW�>�#���T!��L�~�ΠJëL9$�b\�2��/4!�E�U!!�U'��� �F+`y!��#/ʹXp*Ͼ�(�C
^�gf!�ڶM�fg(
=a��p�'��SL!��=9h2ջ�恦R�i�h�'U!�dԷ3�:�s$�A
7e򵢅�ȑ!U!�։%?V�4,O+c�DZc�48!򤙺<k 1[dH7��h@N� !��6.���*&́���9V��-t=!�d��"b-��C�>9�(����J0b5��L�h��Ƌ�K8��jWK�
�y�%1�B(Q����Pd�Z��/�yr*g�2�j���@�@��(�y���|���B��C�F�$§I�5�y��mk.�2D�F�B��'&�y�#Z)<����
�\pZ4Gˆ�yb
��Y��c�Y)|�dH[��2�y�lѡh�\�q�� -"���3�V��y���t�8H� �T6!*�L��a��d$�S�O~�#O��nWv٢�hA't4�H�'�J�ن��~����D9h�S�O:�D8�)��ϟX�T�7�������cS5D����"ߣJ`�	�H�
�����=D�� ���� v��˂GʖS���"O����ӷK�Z$��x�ޡ�"Of]�g���@�cO�LU���"O�@�1�� sp�Cfa��|9$�"O"�YrHȄ/"(	��NX�m���)�S�'���z��<6��\��kԎz>v���|�tt�ƌ�]��pj�8�Z��ȓ/+�E�& 6<�Ѳn�
761�ȓi��(�'ցwG�9��$Q
>����ȓl�a���b��BWLE�)��`��|�~��pG��%�D�:�'�;Ј��ȓ`�i�"
)�A�� �ܠDx��'L�O��'JRn��t`Q�C����� =�m��*�� DkК(?$�@�e1l62̇ȓ3T�D�9�<�3"�J�Y����8�,,)�ߋP�@��DO<j��(�ȓP�2h���Ud���ċ\�X9�ȓJ�)�ΧT���D,Բ����ȓQ�]��Pg5`�� [%�ȓm�FTd�	wpv���R�(�ȓ-����^�/�(�C�O"�ćȓK�,l��h��(y��Fƕ&_>C前 Q�� b�5���+�
֡T\B�	�r��� �p��֨H�_g�B�ɢ$��PUn���cK�Y�B�o�����"�$��m��
���B�	K����ǧ���CɎSx$B�Ik��p�D!�<��	
�)�"`SB�	JC*t*7&��6<�=�2�ޜqz
B��f`��$iňx~�Ͱ�'�)=  C��T�g��H�V������t%�B�\0���0MW�7*(�2����%�B�Is���
�@@�^�L���AŴb�B�	�[���I	�8��x§%�9��C�I�˺��]F����E�o��B�	+�H�X�W�q�V��hZ�B�	*A�8�8�a�pp|���l�+�fB�	�3O�ᑧ%G�*~�a���x�,B䉽|�0�BB��9�t|��A[�8�bC�I8yr�h�N�X/t�a҇4u|vB�I�<�%�6&،k2�Ҷ�W�f��B��"c �+A��H��M���a��B�	�eUr��Q�z��88�DC�Ɇ �� ¦�Q�T����O�v'TC�	�4�������5+�����ά|�BC�I6e�
��%�K8�x�p��,�\B�ɑ~�P�+�%> �ыE.�)H��C�	'l-4T��F�u��1��G_5r�B䉖7��5�',��:���@!	&{hzB䉈I��5��:�X؁g�&�.C䉞=*�`�a`D�`�V�#�oJ� ��C�	�l������D�{��G��C䉖@a� I�%q1��s4�D6�C䉵Wx�d:��e4�'-A���B䉇O������%�d�:��Y�A�BC䉜b�z��ɒ��� f��p�B�	,5�����*�l5�!ʰ���B��TL�h���|}�siǴ@5�C�I�5a	�]#5D)�#�D�$�C��/��W$IQX$y'Hߚ:�C䉣��t�T�ߨq���+D��<g�DC䉬x���� سmx� ���=�nC�	�.C�i��%{M�8
��S>*�C�	����bVXV��3P�+�B�)� $i�w��1>�!B��'Wlt@X�"O�h�AٮHg�M:P��+e*,��"O��h�$� �(���%_��"Ozx��"�.m�|06�F�W���"O��BB��`�,`zD/g�"�p�"O�L�F�� �z���K�i�~lYp"OpmZ3�˟]u��*`�TI $"O��0�a��>!�TQ�Ϝ3a���2"O,YH���
�r��͟��R}ht"O�ѧ+ċf��%�\Hl��F,7�!��o��M`��$��rQ�.;!򄔊%�r�R���c~!��D�<~�!�d�3%��h�K��l�� T�6[!�d�b�nx���<P��V��	P!�.��a��q�.�ᄧ7�!�R�+�p�,Q�����CO�4S ��'����k����E���t1��
�'y��G�
�]{C+��l4vA��'�u�sj��%��hS�b2���'L� ��@ɝh�y�j��@�8�'c�����O~�k�iɼ����'�^���V�
�r��]z�&m�'+�ճ���q^������:|-*p�
�'�x���S12}�LA�D�w�\Ii�'�Z1���b�0��UtZr�
�'7�7<#�qP�ѵd���c�'�Q�,��8��ܶ�����'���h�Ĵ��B6?rN�I�'`xTi聗Pʚ�ńk��<Q�'�q t(�R��p�UM�9�xj�'��4P��%S*Щe��.��)��'چ�Z�X&�|U�$�$2!R	�'1T ��E5�ȴM�*� =9	�'�P5��hS,`�:�)g��%Ͱ���'`�e�U2���P�P�1����'`1�D�!LTy��l�|�Y��'���U㝙PF�J�Ň����'ۚ`i�5�(r����Z���'L-�f�	�z2�]��'Q�Y{T�B�'>P�qw+�$|�H���-C���k
�'��2ˈ��LkD�T�f�np��'�����%dD��Q�'KVҼr�'�$�i�c��k"�;qNކ@���'5��3Q*lq������1�e8
�'��;��X�$	�_�@�Af��x�<��ǃ�l@��H�E>?���P��~�<Q��_�Z�!�j@> ��9V�9T��HTCF�1�Ҽ�A'4(��<�)9D������Q�1�V�^D��s&�6D�*L2,Y9��T�nƪ<��&D�(�X�����}��X�(B�I	>;`�1A�?����瑖YRB�	�'�p�U��.�1c2d̐e.�C�	�O���B#B£?׈��c�9M��C�I�f�]��	��B09ag%�M�C�	�=��e�R
H�/��)�''E~�C�ɆTo��K� �%�� �y�tC�	  u�gZ�J���#�F�xC�	#���Y�nj��pQ
b�B�I�l0���%JB��|��ڏ&�B�Ɂx���	�:R9��j�+wC�ɴA��u�%l�'X��O�
C�	��J�3�K�"O
�ks.�%~C�	�`�x�i(E��D��d�B�)� |��2F�?}V�;Fe��A��s"O�q8PNԃ}Xp�@�C�0Ĳ�!%"O �JO"	����"�w�����"O��;�H��t]*шg!�4f�F�J�"O��`��M3m�Hʖ%F
�}�"O��B0k9TX����$�N8g"O��h_].�A"I�M�����"O؜�r�ة)߸�����i�"O�Dx����1��<ڲ��8-y>K�"ORy����7-�-�#�I(vf����"O�ԃ�.x�ȱ�g�Cc��6"O�i�bL&@::R�ЂyX��"�"O�L�0���Ol��c��N�vD��
�"O��#���W��{wGòu:��@"O� U�ƪ)�9�b�ݳ#7Vh�!"Op@�p�/^�(#��#BP�*�"O��'�̞ᖱ�G���T��a2u"O���#��>�H��@�+ڼŋ"O�y��E�r��*D ł5+�Q�"O��Ǣ�x������
<�L��"Ox�(�.܄:�r�#��3�eK&"O2 ����" hl J(	�-�*�U"O~ w��s�~(c2&E�p�RxT"O&���=|��$���{>1X "O��c���sl�	���4Y@"O�űA#6/����G$�z�s�"O�8��%N}��0 ��ɽ{$
v"Op$��.	�����C�%)Hx�"O !���I$D��cμ����"O�P�V1-�H�2��1�<��"OʴX��I
bs|t�f֥f5x��""ORl�d� �.����K����"O@GJ 17��S�$_l{XHa�"Or<��dƺ��	�#����"Oԥ��%g@�u��}M��:G"OR�{C�;/S���� iG���3"O�졓b�n��2�[�0WtX�"O�t��� {$�t�g��8AF���"OE���$��᳔!$�����"O^Ԡ���3�MZԯ>�>��A�&D�8	��%-[�Y����70���$D�� G�
,�� �-.�(y��$D���DBlT=�G!��v���"@!D�0�E�Ij�1 �� A@�Z�o?D���C��L%6bd�2�dȪb(?D�� U�%zF�`�/ݨo�S�/D��X��Η[�6�` O2tm��/D���7i@�R�|ѐ�/�q ����,D�'��F��߃*φ�h�,D��@�K�1����Be )㲭3��?D�p���Z��ʙ��(ݚS���:�a>D��3���&R8|����?(6�n=D�d3
�����ǉԠq�(���9D��@g�60���-�����f�.�ybΓV�X5��g�:8)Ұ��oV��y��(}��a�,f.��s��>�yŭ�`�5���m�f��fC��y��M"��q"F>VEV�h���y��D�t��!�c�\����eϹ�y��[�{�� ���<��ғ��y����X�$����9�6�؋�ybȼ'����ʊ�I��E2�H�(�y2ω�nQ������H��x����>�y��Ga�@�7�� =/�@�bB��y
� $�eD',c�I+��;<N\
�"O|T�R*�!F1X�a���+]R��	7"O"%����+}��d!�.�D%I�"Or���₦2j��E@�c�2�{�"Ou"U�ry���7`KP�����"O���QjËT�Aѕ,�01|��Yp"O�y���]��%ؐa�$YTf@(�"O���/
���+g��>J�!��"O���`��X@A�
�F1H;�"O�}A�M
�9n����IE�� �"OP��E�o1B���:&|�Ո$"O.��n�DX��!�F�=dx{"O�������L��d(�=ʂ"OJ����6�V]0"
�ku.��"O�!�$�4#��d��I�f ��2"O���'�X�L,���q�֛R�豸`"O��#��D�g,мH^tA���"OV�[�D�tmN�F����6"Oz,��#��,-�(zq���F�[6"Of�
�f�.ui�ě�aȽ��MZ�"O~�񁊮�aX�c $�z���"O�4Y�Y��T9�O;9[�Y�0"OAR���9؜��Q�΄B� U"O�t:�G�
Ð�����%�~���"O^���,��	�����L:[����"O��G��]f��U}+���`"Oʤb���dw.xHF`S%�@ 1"Ol�ң�sDi��OJ�)&2���"O�@2���:NU��Ufqr�t"O�hiF��m�p4��.ޑvdeXS"O���N#��02��|V���E"O��AW�D�(�,��I%�>a!@"O
ͨZR�i!� 1GO`$�䯁��yJ84S\7��z�b�hbC�I�^p�+|$�5��e�1W_�B��/¹9��P�5]f�bG ��A�C�I�ﾹ�� �2N%@�[SMJ$��C䉾]V�Iy H�r(M������C�	��A�З(M�{T�E&3t�C�	ê0a��N�U��$��� �C��I��(@_�D�#��C<�C�		w����ð$'`����ݵ#�lC��&U��Q�PN�%h��;��ZnXC䉖��n���mxǉ�{� 
�'T��Ss�� ՞p�M�)���'����c�7+�r��5���-�A �'�Xtұ�`�J��*�,�}��'TЀyGn�z?\U2d@G�u��'�p1юU,R�x�B�k��d�y�	�'r���fKƽ$����j�b $1�'�H*�ٟub�����G�^���'/NTX���EPp)��O�X�A9�'�Ni�äF�&�Fɉ1$�>&��
�'F�pт8r0�"�+�%~��y��'�������i�Bͫ��L����	�'��ip5D��w��ld���b�l*	�'HH�4@w,qS��N�}"	�'�La	'��&Y�(㋐!}+����'��(E�0��Q��
>%K��Q�'�,�X�G&|dP��hШ`��[	�'IY`$�9.b:��Bk#��	�'�6�[0�[0��Й�?L+�A�'�����pd�)�̎�=�R���'"ݚ5��{P4�L��e|,����� �d�0-��\�"Ȉ �CB¦H!"O���a"^J�>4�뇂O�t�x�"O(-Q�_;b�fL�r�<Z5J1r"O`�R�F�4���x90t�"O �{Vj̬�T��f�9+��	�"O<�;��Z�w��}(���I���A"O��S��O���q��6W�Fl�u"ONa���2^>�E  j����YC"O`�u"
]�~$��O~�F�:C�!�dϺZ��Q��'��(�N��%l@�{k!򄔿F����(�cO�!�+�3�!�^����� 
1��!A��94�!��yU��� ��d����ϖ �!�$�f�2YP20C��Z���1�!��-c*�x��0��Q�e���/o!��4�"��eHV��P�a�Oi!�\!`hi�q搾V�n��2��B"O�m�t�@�B���$Ϩ(z�)b�"O��q�����:�f�\w����"Oԕ8�OD}j<��A$ӱ`[>d{�"O&�3�&U��p�X�#Q�$���W"O}k�#֣p�|-��d��!��X3�"O`���'N<}H�<�c�:���"O��ժ-Uhh(��j����"O���ÍA�9x����/�8��s"O�s�0�`�S��6/^��"O� ���`6��Q97@Y2�"O�	�҇ɵ	�$�5�R�\���"O�d�&�گF��%@�9}�$��"O�TSf�����u��2tp��"O\�rBG�Y�i�CEј!��"O�L"��<�lȢQ�u� �B0"O���1JN�2���`&) �?��ЋT"O@hI �M�xq Ur O#���X"O$9"�U4BX~`j�k�6�$T��"O8�z�&�^9�yXU��Uj<q�b"OD��m_�/�qV�V4XX<���"O�X��쒋e�h�{� �2���"O�u��!�)\yD���ߨxl ��"O�qCd��
i���c'&Xr=�"O�5X��MzXXaq]Lʐ33"OT���[�zV(Ӥ��#B���"Or��1���wV��炌h,J4+7"O�<#����,�"��xl��"O&<�/Ü|��h*��M�	��L �"O����U�;r<ô�^�W���8�"O������"3��1#w�`P�"O>��E'G���Pu�<6���)�"O���a&G!m��� �`�=����"O>%�!���7�}���YT~y�"O�( C��~�Ψ�4�ٝ9g(���"OP=W�U�S�����焑79:ᛂ"O�tjޞ��V����$��t"On��b���T ��3y{�t2"O��(�"2��p�2�P=if�i�"O̐��)H�$,�P2�����@��"O�����	�1`��S(Slؤ"OB��Ӱ$���VƚDH����"O���0�©_�(C2��+=�$�g"Oj��ՋĖc,*�����'��Y9A"O���td�@�!�9_�:@�"O*}���ϘM��d1��ɘ0�H���"OP	�d��07^4��yA�"O��1��Ğ(���R�g�)kPlɑ"O� J�ءb�$Z?��;�ϧ$V� �"O4+CL�vPԫ���{92���"O�l���X%kW"j!e�&[�.|0�"O��i5��G¦A
�c��"O>\+E�͞���7��:g�����"O��ɓ�X���4���yŎ�6"O�M�N]9��3��n̲�5"O�Q�sM�/rp��"�>,�����"Of��R�՜L��������HK�"O0���Ѳ�R/��e�hCG"OD`ke��!,���q�  ��	�"O&�JbnY�9֮y�0@:?�2���"O���W��	
!� �н��"O&���@@�U��xc$��1*^,��"O�u�����z�����H�-��E"Oڍy��<qj�a���"�$�A4"O�iz�G'i%�e��B!�4�:�"OJh`.R+Wg���qV��b�F"OL��2���m"��u-�4���"O�z�I������
�>z~���&"O�E�r✪#�e0rHLv��"O^��Ү[3#	�AĠ�0 ��]�F"O0yC�Iɳ4u�����	 �Fu�!"O���2j�/\�X@��*]���"O❸�hB�,P�D����4>�!�"OZe��^�t�{U�	&N4<�C�"O���t,�/6z1g�8E�`m�E"O$�AL�8\�[p����"O�!B�4,�|0Q�JvR,�3g"O� R��� �3 (�8.�	�"O�Z�Jζn��Yৗ0` �5SF"Ob �"�+$j�3��Z��""O�=��a�W�=J���=��Hd"O&�۵oԉ9N$)��쑘v����W"O��	��T�y�����.3����6"O��Y�`��Ë%r�Ы "O��󆐺�>8��>�Y�*O�AFK���p��G*EtD�*�'[�u��/�(d��A��
46�d��'��<��Υӌ@��a�B���'P���E,KtT�,���R�+� u+�'W���-&H༡��N (>�%�
�'ZXhք�n¥���1�$�	
�'�~U�$`VND9��0{M�9��'��t)�Z� ��!�e�OI��[	�'IX�@�ES7=�.A�dIȘ���	�'��X�EBT�ҁ4lE(]G�d��'��ʡ�/-a�k�@N*N^�A��'/�q�4C.U~@�nەKi��';�<��oO ��A��K���(�'h�]��u".��pf� t�D�X�'��Y�Ch�a��G	)q���(�'v���DJ�>c�P'O�#�a��'���@3o��]Nx!Iw��P4���'T�\w
�!|e�!�"�'igv���']��+�'3^ ��0��4.a���',ݳ�5[��=*P��:*��'Ȥ
/�#̀I��Z�_P�'MN��7j�
�2�i����f1
�'�����ǒyz�Y�+�Pr��'�4�'!�cɖ��E)]6|+���']6 	%5� �b�lΖQs�'h)�e��W�L��* t�r���'��!xL��b��u㝯NxUB���� <��D�	t�a���V�|^�B�"O���AH�#6��`��cVL1QR�<G{��)V��]�ֆ�,J͒���#!�?Q&�@L͚;��Q�Wyɉ'S�|�M�H[:�2s�-
���� 5�y��3kt�{��D����+@(��y���Q��U���x��r2`ط�yB��Q%��C�k�i���s����<cō�g��@�']�dڌt" AYh�<��cG�D1�$ȡb�|�1��e�<)##['u�L9��Z!ټ�Bx≬BL�{"�ї��Z���1�tU��K��?��'plZ���5�T bGD�1�8-�
�'�zIBS�9n&){�h�&,8D�Ȍ��:ORH�A��c!��o�Nx�"�'��lƑ{�͘�>f$��#y����'�ў"}Bg�A	G�����~=���A�<��J\�lM�!(��Qb1��}�<����3%�,&!ƽr��qr��|��`��0G+]���Ď&^�t���<D�0I3LS7�XpQ�N�0�����>Y��~�X����i�p1��ݖ
����S\�a�T'H��D a� ߍ a�4��T��<#ENJz5xۅI�:��]�ȓ`A�a�'#!tL�9{���s���ȓUw^�q���2�Zl����cu`���-�	�F_	S�]� );C���ȓ75LIxCn��}5Z��R��3T��?q���~���d��ʳ ��?�>`	`(�U�<!E�M9��lRm����0E�Q�<y��ǂ;&՛��ϓ�RJD"Zd�<�o�y>t0�K��v�Z
�Z?�M��g[�Y�]���P�h��*�q8�8&��pk��&#��k� ^�E'��Q�5Oh"=�'_�� �0�&�<bG\d�<i�(O�[���P�^4rpF	�t�]d�<���y�6a[b�D/k��QxGi�`�<A��e�,)�R�Z�(����Y�<E�g����0��9�hᓦ�}�<� Gɚ͐��d�(|�����S�<a�#�]p`!�F-��(CvBQ�<�e�ec�Q�B��n��)�6��J�'�ў�'i�~�0E��<B�܅3�	ǋay��ȓe�$"�!YK����q
J�ȓH��M&&��@r E#w@��ڀчȓ+;��A��B�	�Z#��$���ȓ<���¶%Ҫb�b��?@E���L��@+�*s�\���
_���͆�+s�m����H�8yjcJ]˪�E{��O������]���i$�&�t �'�V��W�ٿL��0ڣ�� �x�b
�'����d�4�ks���I��uB��dt�(�}��^�tʄ��c�W���Ua\���$�p��I8m~  j�-:`���R���,ieNC�*k	��p��o�¬�p�:c#>����a����2�D�@�*D�">	��i��O��c¥� 
Z��]"�o�����`a�#VlN��4�]�?����.*D�HC��.>��U��[ ����k������'�ўJ���P���[<��-� 5D���`��6��k�
�<S���Æ�0?ɍ�$=�G��hˢB�+N���8��<��9��`���E��}��I-&L �m@-����ɄrvIpNɬ5��� ��E&�}R��� �8�F�؅G�R����Z&d�>�z�"OD@UF��f���˙�`ʲ��� �	w�'����'�f�api����
I7�(R����l�����2f�`�ԍ�d�Er��#Z���%�R5h��xa�� ,�B�>9�Ă�ͤ}�j5C��9{ĎB�^�DQ�A�%�BQ0�Lα��C�ɇH"�c��=>��9h2؜),^B�Ig9�YZl��T���T-W3 2B��LwV=���Q�Tq#���0p�C�Il�{2B�kH^�s�,��t��C�I!eVNM:��T
l�F�pa�
7+�C�	��
����03��r����C�ɪ04H���N�M����FGH� b�b���.���ɺ�,XV�<X)�H]�3���#T D��J� eKR�H2�X�Q��JҢ<D���͍�"�ě�c�ns�쩶�:��<'�S��4��c���0��t�<���sϰ�ʶ��n�|d�宅n�<���	 D|A��o�/`�����n�<��] Q��7�^�k� ��	e�<�� �:����P��lv�<�4e�G�<��DH/��K��ȴK�B�FA�<��-H4}0� �.��C�e�z�<�D�+[TD=�PgZ��!�aj�yܓw���<%?�s&cۈSb�D� H�:����N5D�<�"�^f�N�����O�I⣋6�	q���'\H��@'K�n`1�h�^E�ɆȓȈT! ��)��aD)u�4�Ez��'cJ�Q�ԓr�� ÷J)N芷�'�F��Ë�6�=�D�߃?�a��'��۴ Y2�*S��"��H���D�4�hO�)_�\����C�'}�8����%�!���:#N*��"[���p O�]�ay�I*v`R�`�(9ֽ��dݷRÖC� H8.���Ɔ���DGA�J��B�I�5�<�!W��~�i��K�B�I�����䆝}f�P�%�*<HB�ɦ
G����N�0u���!��,h���)?�O<��1O��)RL��%�������"s	��r2�Iz�'��$�"�&!�Ą9v�윹gFF���d)�I�D�ԋ�*L��hV'�#Z�-��	��~��)��<���ia���E�@���K�c<�Ԅȓ�|��))��ak{tN�D|���x�~���y�����V'wph��WG4T��r��ң~���gC%{�N�ZQ;�O��Ox�1���Y��I���$a�Ѓ��'=�~�,(	�Lى���z�o�j\�E�?����~:�
݌��=ǉ�wF�p�t��v�'/ў�u:,��d�6Fr�@G��̴[���s����@�n���v��­��7D�4����~��n��D���F6D��B��Q�����*Nf���j7B5D�`Zp�L�k.�8�r���yn�y�s�7O��=Q��݌2��U2���"Z��z�EO�<A�@P�*�����=l������N�<�v���#b�EƑ�=F^)�@�K�<҈_2��x℘_ݔ4��/�]����?A`��#^7V��W+�&��`���MW�<qB��=D֮|p�L�\���z�$9(�<%?�K��ͥa�s�l�6y�D�;D�(�A��.�2"�A�1OMz�.=D�������P���M��M���x��5D��8���%)\�qƦCx3¼p��4D�� ��7�]�'q -���' ����"O8%��ˌp"�P����~!�A"Ony�DE����W��/�(�!��U�<��$ȍ<�D'�V ��,!�gHf�<I�g���ja�J��i����bPe�<��&߂4_ �S��ɿs.ą�dk�J�<���.�0�Wb� "s�H�+B�<	�a�_Y�J��M�]�bPF�u�<!snQ�lF�X��E�^�"ū��Y�<)�A=y�`:W�F� ɎAS%!�Z�<����l!�]�M�&�d�j�&�O�<�!� ��:����|(J�"�H�<a���|qd��C��Y(�E�F�<@��t��3��w�Hmq"c_X�<�&��RvZ���H�)Q�P@���K�<��퇙)�����+A?�(Ƀ�IE�<���ބD�&*�V�x<kb��B�<YA�*uZ
Hl�1W'�������y��T����ӳb�P���o�+�y���kh����eJV-����ܵ�y�y�p���̍�N�(����C�yb��W���*S+�<�t�"K$�y��[�Qn\�+��#�9�P8�y��A<_;j�Ce���h�@���y�k\�Q��9t��	|Nd;QG��y2�ܨ1I����)odi�@ڛ�y�X����eԔ}�py����yr�	��(a�!f�vC6�ч��yb��#�\,	��C������y�J&Z�nY��VP���)��ع�yBH�:k!X���&6M-�*����y��ҕf�~<�+����pR����yb�Ψ �$������<	{�f��y2���	!��!%�A4��#�!�y�`O�w���3j��{����s"��p>�VJ
� �#KA�>�`��cL5:)�UQ�	��iVB��-
´T��^�V͑L�R��B��6L�܋!K><�=��X��B�ɭmF�Z�#K,W&�WD�4ٞ)�
�'�T�K@��+l@�s��\-G.�;�'���s�Nex3E��. >�R�' BɊr L1|�.��� ��W����'Fnt"��Ե%.���]�^�8�'�2�aȉ)]�=�׊ԪV����'�R]�Uk�f H8�aY4��(�'*�d	��M�b�DT���#[s`�C�'J&PP�K*����`�[�hݰ	�'�H] E�G���'E�1RAz��'=�	�`�P�(z-G)O���
�'Z4��gAN4��(;���<�>���'��ɗ�հT�Y�$hR�D�!�'Hb���NϾ!e���V�
#���
�'���
�2��3��Y�x���x
�'jL�!0��$��i�XI4�r	�'s�g���#�he��oϐkV�J�'	�|�p�]�iK�,��)�2f����'n�H�
L�=���`�`1]�h�	�'�0�Z��*���0�@�gF�E�	�'Q��e�ܢ 
eI�NM'[H {
�'�4i(��*`�9��c�$a�'��2�#U�k�D��F5HoZ,
�'�H ��ωP� Ī���� ����'��XR��y\���N[�� �H�'̨��"��6O��d��m8��� \���D��Ԡ�"I�)��(�6"O>�qRO�k'h�Ba�I��Pr"O�pQW�\ yvlkE�F�e�d�is"O@��;��`(���~����"O$�R"��u�j��S/#|�Q��"O��g� 4k�ŚC��vg��J�"O y�AO�>�ԵEǔG�8��U"O`��0���-���dҨa|@X�"O��CRMx��;�C�!\�"O�)c��$v�䨺���	~�pC�"O�3��N><���耊y�9@"Oz A���9@!G�]U���D"Odq ��W3p�,P�a4��r"O���5m�2m� U��K�58���"O�<`�/1⼑iB�Y�����f"O�$��o��B��̓Q�L�g����%"O�D�G�ǂ]��x���Y�U����"O>��AK������;��q#"O��S�	, ^|� �
��`�H�F"O��qnD���A#�F0	�XL�b"Od�3���u��Hc(�H@R��"O �Y"E̱x��л@&̶*=���"Of�i0�B� ���&��F"O$���k��Vm� �T62��4;D"O�}H��ϸ'� :RN�:��`r"O�Ă�>K����p懐i��Y"OT���̊	d��l��h�0\�@�H�"O8t1Ӡ� ��й疴e>���v"O� 
ҙ&������݁f	�i�"O������R�h�&��0nܹ�"On��5EҶK��`C2�!Y@���"O�=�q�=�hYT���*0�"OΠj�CM�"$�C��Zz�ɱ�"O��QV$W�>��⁓)P� �"Op���cF�\��O�=rG L8��'�L�OL%�{!�0X`��-4�{����8��Q��X��e+t��(1m�M~��'���O��E��o� �^T���m��ġ�e�+�y� !U^���fȀ YUb�b�%��y�E??Ր���'�P@3jB5	M���払�z�Ɖc�';��3UaCy��M:V	Ӳt�AP�'Q5��
��~2���Bc*l����l���Eq��� )X%~z���Y;���e"ONu��d���l5��c���@���e�Hy�����D��~��H�O��P�%& �QH��I�A�["�x3�'���xь��1�P�IQ! �I��8�r�]� �9�lś @�+�(���p��T5�2�q�du����ˈT�RVhUX����P4+�"�NX���E�bT)%�# +N������V�@Q��3Q�0Zw:<m	,F�0T�y�>���+.�ZL@��+���ZU�'ϤE�S �*/��܄)�2�요8���Ū�`@���iLec1��R����&]�x�аF�Ƅ8�	ÓJ�Bϗ��3q��80��������r�'`�f�82���!$@�(��h�A�޺��c#ML $�D�D526
��k8!A��F�C�B�����-��ę1?E�m����_������ -F��sY�[X��\	��9�B�i~����;z����$�&�`'oY���%��!��-����dY��\Ʉ��Ad�0q�S	��X4n��/%��P#�W��.Q� �F�Ărb�3�f�(!o��� �.��+"�ʓaN+D���Ż �$2�L ��g2�%s�dz��"I."U�G� 5Jl�����'dD�$�SJ�.%�qD�V�{��)b�ܦ>�L�2�"�E�`�W�ޓ$|�y���D��wCЅP	O���uц@��2(�}C��\S��`8��o�Yp�۵pNȩ ��υ��]����0/�A�D҄[ ]�Վ��
�
���b��q <e�5@0�O��2�$]"
;��b���([�\+&��-wE�	��c��5r�� �]Vtם:Br�I�"S��!���_�\q0��0T���s�� ����$� g�Z]J`+ȍФ0��4Lh�@�S�u}6(K�8{�]��f�*yw�1#�ƙ���\4Nm�H��rp.�J�<�aȌ��HE���r���@BT̓s����F����X �T$osr�׋��!hq��荍/�-P���@�D�)��QE����)��W�
I���S�x$�OL��   ���6�RT��'F�e�ݩVi�
�{�Ŧ�8���:�,5H�`��{e���όs�8�#� ��������iÁE�p����E����U����	ٽ>%2���^�h �X{�o^:]��ݛ����J���&"��T����X?= 6�gy��}��2t#��3+qBv����0=��$E�� 	�����#��]u�QӢP>Pl���ЀÁ8�RM��g�0%�;��۟:��$��Y�Tq:�G0y^�ICw���1O�Ys���.��-O�ma���8�P`����.li�d
Ӧ��t�YR�ǟ�m�v(�f,�hBV�	%�L�k�*�����[�gr�D@r[����k&j���QቬR�^��]�(a�;sΙ�a� ��Ea��đ[�2цȓf"�=B嚨^��P9d�̌U �HZ�bZ�'Y���]��:�'`,5�mQ�(�L��͟�ɾ29��o˻}���&fǠ#���O�5���,OD�{���:w$ن)�����i�����ڠT�(��%LOV�P��4-����ҳ&���pT�'9$���`DEE̦���������S��-�1��?D�q�.�/1FX1���!zz��7�<��B�#�=�Jw�xi��P<#,�02'��<����ȓ<ǜ��#Ո)��\Pw�$���Qi0�@'�Ze$R�ar >��-�ȓ ���s��U�{�b !U��;<N�`�ȓ_��l�jL�~Ԁ�2fFQ�剘1���!K�m�d@g��ysg] H��a>!�D��;V.�37'^�W-��S�NܯXe�@�R��ݹ]����)�B!,�̕�D7:�)EbPA!��C�EQ"E�#kP��rX�Bؖw+0<p4�<��Պb\б�|�<	�.��"�
`r�g*p\��I�N�M<��. ��9���N���PLI�P�l�>���\�̅4�S�W��ӂ�"nH�,��	 K�֌z4��!�y�' ̲ńY�XO���3oLK��{�'<r���+�&�z�R��MZ����O��%�:��Y��'�'B��D�%_%�ΠSa��_ �P�ȓ�Ց$�<ڈE;4�sK�]ZA	�򤐙(������Dj�D0b�A�m�5�1aC'a�!��Di���Խn����ܫ&��e�И4;Z�ۦ�/�OH���
wr��J������W�'=P��cL����h�U�(���j`��a���`��;�-D� �#-��YS4��3f��5� p�h+}�'̽=n`)�d�V�OA�@ۑ��17��!g�ܖmdt�"m�R>�l0|�AS��Z"S���Q����&�'��QP����5���H�e�q�I;+�1�'�W�øx� FBK��	�ȓX��JW��=j)����@� Z�~��'��E{�-�ԦO�>��UF�5 ���^�6�Ujf�(D��3O�lb\,�d � u�qgUq�$�=�i��#�k�3�I�Z�r��`K�*1�!�-Ő5f���tQ��Z�	J�}��Խ`��x�1lלG+z�� �6��?�d��:s�IBd�
,��q�eSR�'�܅���!^��X$?��q���O�tI��R�hp��&D�����#�4Hb F<9���ʮ>���
=��al&}����z]�(��h�f!˅J!�A�<��(ȄoS�3�pɱ
�t$�'e8̡2#���@��O�5K�,��4pQ���D�� &�'��@[��>*� 7�j=�A�%��� �
M��BK���q����]a2�y��p�*�zga0��b�~���fM3טO�>Y��H�bR�qw�,@�b���'��ۑ��=sJa#k�=�����O�,"�V�����l�9�YA`r����+a���[&�'���(�o��V��/%��P���i@�� v�%B�茄ȓ#�N��0�E)�����N����q�O�uˁ!ݭO(v���'5��@�'u��0�'���_ -�ȓR�T����B�-(v�ɶh��5@A̥��X�$ݬ�¦��$�
e������\��c��S!�d�f����I��:r(	�(��a �n�j%�С�!�Ob|�p%�!�t�^�}�4��e�'Ӟ�XA&��6�����Y��d#Bb� &�ʎ@���#�$4D���4ɇ1[�m3�.G�5���+�D~�m������R��&K��?� :u�c��:-��Q�IفL��a�"O������._x����(ϝt6�������˓=r��H�LT�g�;���[��X]�RY2d���^9d��:������#$@� ֌V�F+�u�A#^ox��^ ��>��@D�!o�j���&�p{sk�icΐo
�(q���[yR�4A%�=
dI�/���{ƭΟ�y�-Md��J��L��h�&�� ���<d�2M�4��@#a���_%��I�VP��6���y�I�zs���٪�h�5D�:~9�p%�l�T:���ēh�n���Ȩ��%�G%P Ip�ȓC��u�U�,*!�m�Ar��ȓ՞��uǆ��U#�$Վ��X����̲�U�C`d���#CD����V{N��QHC�V�bhcqf�lEFh�ȓ��q�-0���5D��x��0��-�P����ԑtጝP���8��ȓO�Q�5�(LC"U��ePE4&���ioV��TdU�EtX�0T�ز	aJ�ȓM�ԛ�	�,W�}�@jI.QǢH�ȓ}�B�	�%��6����6!��A�ȓg��Ka��M�2)ن˶?(��ȓoW	�F�D�
�\����[.�(��ȓF; l��疁t�~�1�J�*9m���ȓ)�~���6;������B�͇���+��]�6Ҁ�A�%Q�`�n��ȓт�]�=�BP�r"�le��/��}����
�:�jROC�x�t`��E�DZB�l�X���;�&���fؤtp�j1+!F��M]4yڠ<��%Qj�Z�̀>U۠dɢ!�7n�]��������=Ɍ9�UP�r�B���z#�i↙8d$dls�,ܡaBC�	?N)���!�)%E��ҁI|� B�	#l�ïG4s�9����k6B�3J��:�N©xgy��JÄ$�&B�I�O��Q;ƪ��P�i`���~J�B�	S����"�+������*��B�I�9@4�"KWN�n��+��NC䉘S���$D�F�`䅿�RC�ɥi#`���M�ZP��(@T��B�xg�U҄�\>`� ����˙B^dC�ɖ3���t(�n�SCɈ/+T~C�		���tL2�^ ;t(��XH�B��5_��R���x.�P6�e��B�	�E�-p�*@��`k/\�P��B��`��H��	�dz����M\8#3�B��V��Jv��
E�j�r�FΔ\D�B�b�j��$��P�t�`s#���C�I.W���a��3�N�@G��gАC�I�L",�c#,UTHj��U9j8C�	�y��mag�A5�$y��7U��B䉚;��:&�v�HY¶�)C�fB�	�� (�'��0s8���N?y�B�I,Q��ِ��"0.d�h��̙`�lB䉼x���c�J�M��c��	L B䉌_���%O�	:r8Qҥ��B䉽N��!��޷ S<�B�	�zL�	a0oPӦ��(x��C��%mf����} N@��Jʬ\�C�I�?�|�CD��X��L��{�C�Iy�<�8C��|���։¢B�	'4��J��;�2@�7@U�B�	�D��H��� Y�� 6�Ҋ<�B䉦P�L<9�/`�Qq��0:ưC�)� �u!��N0^�ra�ԯ-�<�X�"O���� &�޽�$�Q�� �E"O��P�.��X��$�UV���"O���⑘7����A� �ZG"O�u�p U\�p`�^�3���"O�Xڶ��Jd8���_%�X*�"O�j�FY� ����jA�c!����"O�h��d�'6xX����+d�XF"O<�X� ¨mo��q�E��x쨒"O����˯1>���2'�)�`��"OʤhĞ�,_��R3�H%sV�s"O���CJ�
�n����U�i�"O���ě9:D�\{��5#^鹣"O2T��F�N�c�� {�b�H"O�MCD���W�� 6��c�X �"OԒ�����C�U�d s�"O(�J��;"Xx�t!��'üI۴"O����Ny�<�������X��"O0�c�)+^�0ig��7va9��"OP3��&&����FZ�\mHP)�"O�t�4�īb ;�DY.-BnX�"OLAgJ/�҈zf�]eЬd�$"O��P��iL<��%���5X�"O�X��+�^���۠�F@Q$"O��tNG�U���K�� �5�(P�!"O&�����x��@�D�H@(�"O2D�Gf�!�����)u:��"O����D�>\����/Z� L�4"Of��Sc�N[�2EżC���"O�a�3�Y(�h����*|�1�"OVq4e<8�1��
�N}n�@6"O���_�7�x���̈́~,@�t"O�)�Ȇ^�d��N]c�$"O��;��"\�
�m� ���B"O�XX�(f��
E+ڭF.���"O(�#4��&Tq	��}�"OB���*Nj�qC"矴P�K�"O�|�2$�0�V�9w��%	����'¾ԙ (I<Pv8�*C�]�F`H�'7jhCB�#!z�b��`�,�h�'z��ʝ g�Ѝcu���̃�'lP�@CK�(j?��$c�8\�z<��'��at���n�d��$�6IR&���'^�9@���,��8*N�D8�Y�',<@��LYAۆ����ػ4i�p�'�REZ$�B�Q	`-�v`�7N���	�'ަ���KژS�( ��eE	0����' ̝����Y�8����C�0��<K�Ef���ǹ����"
�iŤT���*T��i� D��Ɓ��v��Ԙw�#Z	́cf�4��9q����CE�O-�-��"�'uֲ���ɴng����i��is��OԨ��!׽7Vy��V��E����y|�SsA'
�j�P*�$ky>�i�xz2"ػ~���.8�r�G�_�'|@�&,��&"Q>b�k|�n8Y�c����I��F]>*.z�S���@4��z�O�%]h��
Ó4�dPQ�H�� A*���T���B�놔v���ه(0}��������%!56�(��.6�jL-u�v�#5Kăy�09��/N�j�dYQe)Wz���.)�,$�����ur���hW�N��B��a��'�b����8~�$����yz��H?y ��I���B����bK��I0�O� c�DΛN�2P���,x����Ǌ)�v��w(�v���'��~9�n��w���z���	�(O�4��MN�Rk�8�G�Xs��Q�2ቼ^P�Z ��|i�%O��h� �;V�X:u� Z�<��q/�[�����K�U�����&�hRS�G=;�T�vH;S2uY���%3�v��+ON��Oh����Ǒ)5� UR'��") T��6���O�Ι�`U�n,�B�خj�����ޔ!@K�>��8����Q�����Y����qN��|7$A�qe���u��. �l��(^O�� xA	c��N��ٛ�KP�.�dЛ0�'��Y�UH�P5�Q(�K
C}R�˅�E�|4���$�Y�N�TS���]\(�7���M����հ����ł}6����O���-Lق��$��%]������S�"��b�����Җ'����ĭ�(�~�iz4Q	b(쟀x� -��0���o�}�e���
��}+ӡ�O����
J���Ul˂��G{�ԂҦ̆\^B%��Ȁ:�z�I�7b0䚢jH�d@��c��<lnEisƃ/*��hK6.�ެ[����}���!�
�%�5�@�j(#�Ŗ�n%��K��,P�(��21^xA�"�<Q�bP8��X�EE;�əs*tX����?V��qs� �.�����_*w�	( �W��~�Ѯ
��4e0x<�(�(��M���?6���:V�'|O�83� g���r�4݂�`��D�7Ֆ�0.�2��d��C�Hk�b�������<|�!f��Y��a�s�<Y�$h�~a�u�@~"�%�#�G/FJ|H�6ɷ<Q��:��A:�	8������1��P�*ҭPBA�<�!��	�΀&_;+ta��`Wj��đM�Mc�O�z��>1e�яr�a���-�0#^��g��"�=�!D�֥]�sT�&}�"h9��R-���be�|����o��.a\YB
ߓS�x��4E�::�:8�7�J0<�L��ɣ|���S���<��$�2�BCb*�mC:�����k�<y'e#Ġ��!e��O`"�)G�e�'䬝���f�OtY���\�`9���,����'���A�$>_T�hu,G�&M�{�'�*� u���P��)!I�jܢ�'��*sR�9S��|����\��y���Om�����2o�Gc�#��<�1@�d��K�|c!��)g�訢��h���;D���5fY�tTrM;T�?l�� A�*}b��|��e�U>��pG:�Hֆ~O�%c3$4D���GL�&����o�8�01�D�t�@�'IV��$@�ΘϘ'�� �/ޖ{Ծ\�p�[�*��'��`c��8�HKs�!��Dx����7|(���� �6��}2��&�ҸD,��A���0<)�&M2&nxI�Sl����Եw&��Q����q���h�!�d�!z��A6����hf�T�	i��7=#xx,�cؤF���@X�ā��?J�<������y��"l�	x���#G�t���ƛH��<��Q�\���c:c>c��"d�9�D��(A�P��bH.� �Bd�t��i��NڃA*�
�-#2����8�5��	6~��2"Jw 
�QO�3M������W$�;! x8��|t��`��ΊRi�F���G%�P�ȓ�@i��ܓ=̖���S
I�t-�O�%@�&�L�R��	(R/Ui S�$Lh�
���k�5��@I�h
�:8D�q#�΂4x�'9@�a��:��]�f���O��X��D0(b�,�d�T�3B D� �����q�4� E拣*� ����>م鄩1XM1�$(}��iB�$|� �_�M���t� �!�D�5�8��� ���"a��> �P�'���	�y4��O ���H��Np,D6��U��#�aBD�:���U	ӝ���,��P<X�paCX�:Յ�I�^�T�f
�W8�Y�=`�"?1�E�7U/䠀�)-��Z���r7�<O�P�X� d!W"OҨ�N�i!r:��iB�52pW�@#��ъyq|P;�>E����>F�ԅ��D�u�d9����y®V>/�4�Y`�g�ԉV�D0r��������c����'�\a�u�O�	x���E�ҨY������svΡ��+ b?@��Ċ<TYX܊�a��7j�
�#4�O|D�ïh�%���R����!�U�'�����@V�[1�.��X{��(�P䒯8�H	G"O�(���f�R���S�X�������K��qO>E�6흻8�9;Ug0�{(?,O�)bV�Nb(�'䪍�d���
8^X�����r���@�'���FC'5Hx�� 	?���O��
��S�{�8��OJbxA3a�:�|aE�	�c�\3�'Y�xĄL���q��A*_��,A��̦@M�ɺ�pi���=�3�ɘR6 ��&*��i#%�ה,��C�I�P00� ���t��|'��.߸.���ڒ�J�O=��7"?�O��sRH!C�ɐ 'ؼB�L�3�'��H2̇>��	�VP�|��,СS�#Rg �m��6D������7y������eS�x �+7?q5MA�+žh�����蟎t;���lȰ�DQ�65��D"O
�Ra��E������	Hv`��*��v��".E�Aeh�g̓G���V��$/^�`W��P`�����C����'��K���猏<Ɇ�2�8Lv��h1�ʹ��>y��P!d]�D��=�B)$m�l�$���s�E�G
�`y��P]�6QK��בiP��
K�y��X���8a3��4d^z	���^+��I�h̶�:�a�W�a�d]�J]H *��A�������yR �@ @If�	(C�N��⇘f�$���������ē�AKQ*C��p�a� (I2�!�ȓ`@ [c��}�@	�P�p��x�ȓ}��Me��
3�N�&�����ȓv�p��Ӫ4~�"a��I��j���ȓ?@��b J�u��)�D�\-����JUXqK��1$�r}�����\�ȓp��MPEB�^<p� #l$]�
��~xh����x���hߚ�l=��_��g-�>O��3bOՐ<D���=��U,�$TsC��zņ�����*�"Cg�3�BS*1p�ȓp�Y��J�x���䁕�~���ȓx2�i
a!�#���*%.���Q"O�[��˹
&>��Bo�@�����"OB��#�8Z'���V� �"Of�X1L�#v�;V�8����"O��'/߲ov�����J\p��*�"O�(�S�R�0��8VfP(D���(s"O88p�KE;b=�p��$��(�ؙt"O=Q쀲@E3?ް93�!��?w��8JT��V�-{%L�h�!�G�N_R(�d'���:�'E�m%!�]$&�̱S�'��vd:����^�<y-�U����ۨ�j=bc�<�㘇d`L�F��`�H��V�T�<���MD���C���'�U�<��Е|�`	sV
8n�#Gd�^�<�T^?�:�@��=0�ɲ��Zq�<�*+0���a�Ҿiq�hm�<�a˅��ޱ���ǂ8�� �Jj8�ܸgcɫ,�z�
���tM�)	E�ݪazT��F5�!�S*�`���C`m| z�i�y����)+C���A�%/�Ꝩ���yb.�� �>�+f"X��%���y���¡Arb�K0N���M�y�bS�")C�f�A:�P؃�R��y"e��V)��2l�H [�>�yIб#�j�h�c��aP� WΙ̨OoZ��x��~*���3JD*T����,���F)��0-�-�$Bd?��m�1H�L��i�k+bԒӁT�&�0��5�ڒ`�p���F,;@�KR��_w�=)��O`�ZL��r�Q:X�$��
ԻVdH�UA�	,���e�H=�H�K�OQ>7͂![3z�*��ޞv��l˒��,�u#�p���I�i̷����[���*���2�*����  c �<���-Ok�O���8�	��}QzPJ�mΠB�,���Z����'��9xP�����Y&	��� �
�P"\HB$&p�u�H>)T�B%$t���r=Jq���$P$L�p��S��ĕU؞�YHA�{C����J�����eo!D����E0�ͻ� B��[Ш=D�t�6+# 6��0
�}9��(��7D��CC��?��@+��	�~-�p8��3D�`�.� >d�(bF��5�T˂�/D�� <Y�j�qJ�i��
FC8�X�"O�|hf O�u��P��4I�M�"Oµ� ��[r��A�+�9&B)Ӓ"O4�:�f��2I�wj�{�~P@"O�9�LΊ)�@����J��1J�"O���c,p�
��N�H|x���"O:� �*g�8���YA�t�+�"O�+v�C864�Z�G��9� xx�"O�@�jپU�Ե��@�F��Ku"O����+E�qZ�Xã�*@c���@"O�uy� � *�p�UD�7���c"O^�lO�H-�;��H��9�P"O:RU��v��9SE�V1m�v�0�"Oh�J�Dׇ�0M�gU�"�2�	R"OZ�ׁB�p��E0�e(�2�8�"OX����]��|*�DO����!�"O�%��lM�)��1�Y�NP��`�"O�����2VVX󄏇pI�H��'B  �qf��>B��kIǖX���'��$r�c�>kK�� $�۱}^hx�'�`A�3I�< R��fc�!+ ��'2�� ,P�[,��W�a"�4	�'l��"j#[�n]�a\�e�֭��'�L�i���%���jZg�}a�'Y��Hc�Q�@����Iƪ^�TLH�'@z͒c�.u����� 2 [f	j�':�ɓ�N����CHf����
�'�f�8gR�'U�e`Z-` .���'�LY���$���j�)�@�����'|n�X-�2 T�{��G*=,���'�R��� �
A.�&��6$$�y�'�D5+�iO�;�D����2.�����'� �;pm��MƄS��6 ��UP�'���:��yᦠ��A�����K��yR�ֆ}Z��&B�=���f�ybd�6Y��iw/!<[�A�&c\,�y�	��r����܄5��q���Q#�y�H� �܁5n��0��\颥�?�y��V�hNKs�ӁX�ԙc����y2#��m�M�֫�)9����tH�9�y�,҂iD�r���4��R�g[��ybb�{�6��С�z{�P�� 
��yD�E�Ƅ96NI�w�^0�[<�Ņ�bLN��u�}�R��Ҩ��n,��ȓ
���[�I_9U����6��ćȓ����w�/H���90��1L��ȓ!�l�\�sQ����gϤ)2!���Z*4lѵ��%w��`*UH�	)�!�C7"UQ(�.�~Dd��͆�R`!�[���3�*�y��h*��E�!��P�o�)�"lV 6��թ�",!�d`��)�QCK>%���!@��6* !��۰B�:�+�oK�+[�
pd��!�=]��\�@�/"r�ҺPW!�8s'�A��0{v]H3�G�OH!�D��Nvt)��+��=a�!��K�?!��!Y���B�6`D���ŏ�3!򤞟2�(�E�B�q	�hR�_�e�!�dV�jlP"�����9R�'�!�Zl�|Y`��Q�>OTBԯ��!���5|��=�%i�$j��\���T=Q1!�ĉ2o�>�5�ʜ �8���ܗ�!�$��
Y~�22��?�0�B@�(l>!�=�}j�
�&V������^0!�� �����Ry�n̹$3��:�"O�Ep�)��D��ȍ`�>��5"O @�k�9]���A���Z��"Oz	!i�>����Ŷ\�j)Av"O%��c_�0�>	-C�Q;�(
�"O�����<A����пS����"OŲ7�,���ءA�sNH\�"O �����YK�㊲l�P��"O���Q�z�T`₁��2�|x�T"O��)dE����ۖJ�K���2r"O��r7��h�H<+�R�3q*���"O}a .=:᪷(ɜ:�Y��"O$X��M��.�BTI7�ٻS��)"O��+�����p�����z"OA�vY*Bf�<� O�����"Ot��iʐ6�89pp��ܪ���"Od��fEF�g��Dz��V�)��Cs"Oҹ�4��>hS��{7GQ�\
XĐ0"O������
S��m��x��"O��եl�aĂ1E��P��"O2P�b&e�ĵ����.\�<��"OVp�&Ab����.		xa��r�"O�¢��O��dq�N�S骜+�"O��RiZ� R5yҁ��"A�d��"O����g¯1ޅ�q�Q�>�H��"O�� ,]&s*^ �7-J="�4�`�^H<QK "��Āv�ҭ�i��'�\�<��B�<7��M+��E�;�h�ڄ�W�<���;�z�s'�+P��UR�  P�<�V���b͖�#�o��K��zp�D�<�'��R���&���IU��a�B䉌�
��ѮV$?��mPqJ�gj$C䉀u�t�/���I�&6�B䉪M�V-H�d�(f�)(*��k�B�I�T@t�B�S��	qC�D3v�B�	�r�\�zFF^�M�@Qq��1),DB�I>7n��yM #m��p��R�CB�I-�z�XpA��x� #J�	gp B�əvu�<�v�|�h�bWe�М3�"O��9�Ό�+�" t�l��4H�"O�diɐ�r9Pܸ�G�W��!k�"OΡ�#�QI�hTY��;?�"���"O
	���"<+�H�1JA�b�J!��"O�2U��:�\*��؝�0$�w"OZtㄋ� @���!�oI�m��\1�"O�!U@6L �`I�,ʻMm�}"�"O�86��g�iq�*��XHP��"O(<cq!]3���H���\�媖"O�5Aͅ��.���&֜{nt-�"OJ��!�D ����tVJ�Г"O:}�����"����>#=�}��"Oz��FҚE�nyqfF$;29�"O�e���X ���%P���e
""O�1av��9.��p3&V�w�*P�d"Op�`Z2���` �0	�-�d�H�yR��V^���JԪ.��H(�])�yb�¬`wlL�k��0��h�Ԇ
��yRa)E���{Ċ�/x���'��y�	�*!]�!�!�������y��+¼�QU�ЂG��,����>�y�LӍ�I+�A��C]`��ԁ�y�*2T&���$����a�:�yBc�2���@�dC�Q�Jdi���y"�е4Z@CH<��S`b�
�y
� �-��?^BZ���M��U"O�h��Ե3�a��
5��"O��F�R T{��9B�ڄz�B��"O2<�щ��6����(QzE2"Ob�ڐO�
{ߔ@���D5:��s"O�\�w�N5����/0&��"O�%V)����C�F�?/y�k5"O��Æ�}'�Ƽm:t���"OT�Y��̏:_�Mه�Q,���"O0����u�ބ+��EY�"O�%�5D�?販9p�I	Y�nA�Q"O~� P��u&�ҩK*��"O��z��F}:�L�aB�9��	�"O����ka�`jՁ��B�t"O�L���Sr�� �Z�Xx9"O�9�2)ӽ�`��U��� ��a��"OH�jlt3�ÀH߶2�<�Y�"O8ź�E� �
����˕�2EI�"O���_���<䨀Z���$�yO�;��g�;.n�� F(�<�y����Htd)ʓ ؍�ع�4�S��y�"�g9�����	%}n>��d���y�Ϛ
2��e�4�W6"͐��s��)�yҍ�1x$������(���Ě�y,�R7���_T���� �y��R{$���n	V�-���	 �y2G[��c�Bы��h:�,ɉ�y��*�T�H��A�?�z�3cɋ7�y�NS6 )���@I�c*�s�с�y��$9ܽ�� U�Xp婟2�yBd29�y�F@Z H���Y�d���y��1k�]P�)�G��us/Y��y���o���y�d����p@2�yҀȱq�� ����8i����y�F�5Z�z �*G�U�����9�yr�и3����<w�A����y�'���j�K�G���1B	:�y�jS!s�z{�̚�=z��M���y������h�L�8�X-[R���y�D��>��Q��+u�Q`���+�yҡ�w����C�NL��qgQ��y� ̱_�ج���\N�Iv�G��y���x�RXH���dҘ�y��J4{v�\�5%ăw�y������y2	��nߔixP��j�@a��
�yR�P+X�Z��ʗ;k�����y�� �� ��u�z���>�y��Ī6��d�B�\<�J���T��y2�#]rUXEHY�7:
�ye@Ƕ�yr,J4o���#�̟*X��xi�B�1�y�o�=%���6�"�1� /�0B�IB+LxK7/�(#}U�A�c B�I`v Xf.P�e����։�;�.B��2M	|- �G^6�r��jA/F�,B� *�Q�B�޽�R8�у�RHC�ɦ��D�Dį&����fb���C䉳6_���V��|�f��K�\C�ɬb`pr0e�%^��q� &$�8C�I�f��8 ���q� �!����C�	�PL�QS�ןd��a1�C�@Z*C�I4R�v쪗m�	.��Ů,~�B�I�Czbh�'��5Gi
���-?#�C�	?\��#RG&, �Q!�mx�C䉁0JZ��	Ã#�䨹E�
!A�C�)� l(��-�!�@����|@D��"O�#��9J��- ;�L�r"Oq��/ߎ%�rX9�m��gGd�;�"OR5�A�v<��C��+���e"O$Q�c�8�.����U�T���"On����46��يeFЁ(`ܠ�"Ori*`��&pzśF�Y����E"O �#�X Z)�5˲��-�ذZ��'j���}� ��gGl���P�C̼"�Z���ئ���П�Io�i>��	+3t(`�\�&� ��n�.(m�Dr� ^9U�a�N��}���JܼX)��zA�ٯ_7Z�a��Q6,�
Q���γ$D|Y�V�	q�ў<z�mm�L8�ʥ�%��Cn^�˔Iӹ&���ئ��jy"�'��k��2f��D[1ü�S�珃i�B�ɳ:��q�DFD8�I����N�<�$�i��$d���lZ���S�h�R�H�4�?��O�*Ҏ�!e��LN���$Xd�	ߟd�	 ��'�`����@��CK�*���$!�1Nh�d�e�	�)4`�Q4I�ܧV:��4g�C��{���� ��D~��ť�?I���ħY����&ݞ[&�eۤ�*I'����'a��|B�S�" nE*�#��n�^,�A��Z`��d���El��]��6�	�5��Mh�"�	U�6	��X�!@����$7���nZ�&q`cY��|�	�716�����rT�Q��/}��'�"Kʜ8�Di��Ϻ}�nJ �����w"y�6O��[JX�FcJ�T�P�J�1�ӕu�s�ݺ8J� z�A�h��'�ҭ���?��i��Ӭt�0���(��Bșקۦbk��Z/O$�d�<���'�l](��T������M�k�6T!���c��lZ۟���!�Mè�hU����I|�YB���(^{|��拖�ؕ'��f�{�(���O��D �Jp�A��R>���k�K�2W�d�O���%	3lO�Lx�+V>R��@�C�'Æ�qÃ��d�Y��*�U�3�ɋ)��#󆆸�`x���'e�ּx�O����'�J?��O���kӐ �R�ѓo�"Љ$��y��Ի��	}X�d�V�Ѣ��tbض����gd��H#�4�?�I>ͧ�?I(O��q�T/"T�b��U6Tb\|�Õ-�D�n៼��ӟ�&���˟��W���E��T4tt\,K1����as�'�O�e	W�M2_:�xwH
o�<�î�]�j��aE�A�\(�
�A�1n�#�0�Q��I�kS���J�Xkj,`	�ډ'��O�O������F�(�ݸ�$́��B��<P1.鉐+�!����5��5���'�47�y�'qR��Kr����>����)m �����u����)�'���'�SU�|�����h:�mdC�7�`�2�F�'�1q��9�B! 4�~*ȓ2�x�%c���� j�F�y�'�p�9��?AG�~j��˙[D���+�.k�^Y{��V�v���'��O�)7�I3J�4�#-\@�<����3����Y�YH�E�T!A�`��w�0%�0���Z�'����͟<��'̪� @ ��